// This is the unpowered netlist.
module mult_32 (clk,
    done,
    init,
    rst,
    A,
    B,
    pp);
 input clk;
 output done;
 input init;
 input rst;
 input [15:0] A;
 input [15:0] B;
 output [31:0] pp;

 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire \acc0.A[0] ;
 wire \acc0.A[10] ;
 wire \acc0.A[11] ;
 wire \acc0.A[12] ;
 wire \acc0.A[13] ;
 wire \acc0.A[14] ;
 wire \acc0.A[15] ;
 wire \acc0.A[16] ;
 wire \acc0.A[17] ;
 wire \acc0.A[18] ;
 wire \acc0.A[19] ;
 wire \acc0.A[1] ;
 wire \acc0.A[20] ;
 wire \acc0.A[21] ;
 wire \acc0.A[22] ;
 wire \acc0.A[23] ;
 wire \acc0.A[24] ;
 wire \acc0.A[25] ;
 wire \acc0.A[26] ;
 wire \acc0.A[27] ;
 wire \acc0.A[28] ;
 wire \acc0.A[29] ;
 wire \acc0.A[2] ;
 wire \acc0.A[30] ;
 wire \acc0.A[31] ;
 wire \acc0.A[3] ;
 wire \acc0.A[4] ;
 wire \acc0.A[5] ;
 wire \acc0.A[6] ;
 wire \acc0.A[7] ;
 wire \acc0.A[8] ;
 wire \acc0.A[9] ;
 wire clknet_0__0457_;
 wire clknet_0__0458_;
 wire clknet_0__0459_;
 wire clknet_0__0460_;
 wire clknet_0__0461_;
 wire clknet_0__0462_;
 wire clknet_0__0463_;
 wire clknet_0__0464_;
 wire clknet_0__0465_;
 wire clknet_0_clk;
 wire clknet_1_0__leaf__0457_;
 wire clknet_1_0__leaf__0458_;
 wire clknet_1_0__leaf__0459_;
 wire clknet_1_0__leaf__0460_;
 wire clknet_1_0__leaf__0461_;
 wire clknet_1_0__leaf__0462_;
 wire clknet_1_0__leaf__0463_;
 wire clknet_1_0__leaf__0464_;
 wire clknet_1_0__leaf__0465_;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf__0457_;
 wire clknet_1_1__leaf__0458_;
 wire clknet_1_1__leaf__0459_;
 wire clknet_1_1__leaf__0460_;
 wire clknet_1_1__leaf__0461_;
 wire clknet_1_1__leaf__0462_;
 wire clknet_1_1__leaf__0463_;
 wire clknet_1_1__leaf__0464_;
 wire clknet_1_1__leaf__0465_;
 wire clknet_1_1__leaf_clk;
 wire \comp0.B[0] ;
 wire \comp0.B[10] ;
 wire \comp0.B[11] ;
 wire \comp0.B[12] ;
 wire \comp0.B[13] ;
 wire \comp0.B[14] ;
 wire \comp0.B[15] ;
 wire \comp0.B[1] ;
 wire \comp0.B[2] ;
 wire \comp0.B[3] ;
 wire \comp0.B[4] ;
 wire \comp0.B[5] ;
 wire \comp0.B[6] ;
 wire \comp0.B[7] ;
 wire \comp0.B[8] ;
 wire \comp0.B[9] ;
 wire \control0.add ;
 wire \control0.count[0] ;
 wire \control0.count[1] ;
 wire \control0.count[2] ;
 wire \control0.count[3] ;
 wire \control0.reset ;
 wire \control0.sh ;
 wire \control0.state[0] ;
 wire \control0.state[1] ;
 wire \control0.state[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_121 ();
 sky130_fd_sc_hd__inv_2 _0491_ (.A(\control0.reset ),
    .Y(_0171_));
 sky130_fd_sc_hd__buf_2 _0492_ (.A(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__nand2_2 _0493_ (.A(_0171_),
    .B(\control0.sh ),
    .Y(_0173_));
 sky130_fd_sc_hd__buf_2 _0494_ (.A(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__or2_1 _0495_ (.A(\control0.reset ),
    .B(\control0.sh ),
    .X(_0175_));
 sky130_fd_sc_hd__clkbuf_2 _0496_ (.A(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__or2_1 _0497_ (.A(\acc0.A[15] ),
    .B(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__o221a_1 _0498_ (.A1(_0172_),
    .A2(net7),
    .B1(_0174_),
    .B2(net247),
    .C1(_0177_),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _0499_ (.A(_0171_),
    .B(\control0.sh ),
    .X(_0178_));
 sky130_fd_sc_hd__clkbuf_4 _0500_ (.A(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__buf_2 _0501_ (.A(\control0.reset ),
    .X(_0180_));
 sky130_fd_sc_hd__clkbuf_4 _0502_ (.A(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__nor2_1 _0503_ (.A(_0180_),
    .B(\control0.sh ),
    .Y(_0182_));
 sky130_fd_sc_hd__clkbuf_4 _0504_ (.A(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__a22o_1 _0505_ (.A1(_0181_),
    .A2(net6),
    .B1(_0183_),
    .B2(\acc0.A[14] ),
    .X(_0184_));
 sky130_fd_sc_hd__a21o_1 _0506_ (.A1(net229),
    .A2(_0179_),
    .B1(_0184_),
    .X(_0158_));
 sky130_fd_sc_hd__a22o_1 _0507_ (.A1(_0181_),
    .A2(net5),
    .B1(_0183_),
    .B2(\acc0.A[13] ),
    .X(_0185_));
 sky130_fd_sc_hd__a21o_1 _0508_ (.A1(net228),
    .A2(_0179_),
    .B1(_0185_),
    .X(_0157_));
 sky130_fd_sc_hd__buf_2 _0509_ (.A(_0182_),
    .X(_0186_));
 sky130_fd_sc_hd__a22o_1 _0510_ (.A1(_0181_),
    .A2(net4),
    .B1(_0186_),
    .B2(\acc0.A[12] ),
    .X(_0187_));
 sky130_fd_sc_hd__a21o_1 _0511_ (.A1(net192),
    .A2(_0179_),
    .B1(_0187_),
    .X(_0156_));
 sky130_fd_sc_hd__a22o_1 _0512_ (.A1(_0181_),
    .A2(net3),
    .B1(_0186_),
    .B2(\acc0.A[11] ),
    .X(_0188_));
 sky130_fd_sc_hd__a21o_1 _0513_ (.A1(net188),
    .A2(_0179_),
    .B1(_0188_),
    .X(_0155_));
 sky130_fd_sc_hd__a22o_1 _0514_ (.A1(_0181_),
    .A2(net2),
    .B1(_0186_),
    .B2(\acc0.A[10] ),
    .X(_0189_));
 sky130_fd_sc_hd__a21o_1 _0515_ (.A1(net181),
    .A2(_0179_),
    .B1(_0189_),
    .X(_0154_));
 sky130_fd_sc_hd__a22o_1 _0516_ (.A1(_0181_),
    .A2(net16),
    .B1(_0186_),
    .B2(\acc0.A[9] ),
    .X(_0190_));
 sky130_fd_sc_hd__a21o_1 _0517_ (.A1(net178),
    .A2(_0179_),
    .B1(_0190_),
    .X(_0153_));
 sky130_fd_sc_hd__a22o_1 _0518_ (.A1(_0180_),
    .A2(net15),
    .B1(_0186_),
    .B2(\acc0.A[8] ),
    .X(_0191_));
 sky130_fd_sc_hd__a21o_1 _0519_ (.A1(net168),
    .A2(_0179_),
    .B1(_0191_),
    .X(_0152_));
 sky130_fd_sc_hd__a22o_1 _0520_ (.A1(_0180_),
    .A2(net14),
    .B1(_0186_),
    .B2(net168),
    .X(_0192_));
 sky130_fd_sc_hd__a21o_1 _0521_ (.A1(net230),
    .A2(_0179_),
    .B1(_0192_),
    .X(_0151_));
 sky130_fd_sc_hd__a22o_1 _0522_ (.A1(_0180_),
    .A2(net13),
    .B1(_0186_),
    .B2(\acc0.A[6] ),
    .X(_0193_));
 sky130_fd_sc_hd__a21o_1 _0523_ (.A1(net148),
    .A2(_0179_),
    .B1(_0193_),
    .X(_0150_));
 sky130_fd_sc_hd__a22o_1 _0524_ (.A1(_0180_),
    .A2(net12),
    .B1(_0186_),
    .B2(net148),
    .X(_0194_));
 sky130_fd_sc_hd__a21o_1 _0525_ (.A1(net154),
    .A2(_0179_),
    .B1(_0194_),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_4 _0526_ (.A(_0178_),
    .X(_0195_));
 sky130_fd_sc_hd__a22o_1 _0527_ (.A1(_0180_),
    .A2(net11),
    .B1(_0186_),
    .B2(net154),
    .X(_0196_));
 sky130_fd_sc_hd__a21o_1 _0528_ (.A1(net170),
    .A2(_0195_),
    .B1(_0196_),
    .X(_0148_));
 sky130_fd_sc_hd__a22o_1 _0529_ (.A1(_0180_),
    .A2(net10),
    .B1(_0186_),
    .B2(net170),
    .X(_0197_));
 sky130_fd_sc_hd__a21o_1 _0530_ (.A1(net175),
    .A2(_0195_),
    .B1(_0197_),
    .X(_0147_));
 sky130_fd_sc_hd__a22o_1 _0531_ (.A1(_0180_),
    .A2(net9),
    .B1(_0182_),
    .B2(net175),
    .X(_0198_));
 sky130_fd_sc_hd__a21o_1 _0532_ (.A1(net218),
    .A2(_0195_),
    .B1(_0198_),
    .X(_0146_));
 sky130_fd_sc_hd__a22o_1 _0533_ (.A1(_0180_),
    .A2(net8),
    .B1(_0182_),
    .B2(\acc0.A[1] ),
    .X(_0199_));
 sky130_fd_sc_hd__a21o_1 _0534_ (.A1(net149),
    .A2(_0195_),
    .B1(_0199_),
    .X(_0145_));
 sky130_fd_sc_hd__or2_1 _0535_ (.A(\comp0.B[14] ),
    .B(_0176_),
    .X(_0200_));
 sky130_fd_sc_hd__o221a_1 _0536_ (.A1(_0172_),
    .A2(net22),
    .B1(_0174_),
    .B2(net157),
    .C1(_0200_),
    .X(_0144_));
 sky130_fd_sc_hd__or2_1 _0537_ (.A(\comp0.B[13] ),
    .B(_0176_),
    .X(_0201_));
 sky130_fd_sc_hd__o221a_1 _0538_ (.A1(_0172_),
    .A2(net21),
    .B1(_0174_),
    .B2(net183),
    .C1(_0201_),
    .X(_0143_));
 sky130_fd_sc_hd__or2_1 _0539_ (.A(\comp0.B[12] ),
    .B(_0176_),
    .X(_0202_));
 sky130_fd_sc_hd__o221a_1 _0540_ (.A1(_0172_),
    .A2(net20),
    .B1(_0174_),
    .B2(net193),
    .C1(_0202_),
    .X(_0142_));
 sky130_fd_sc_hd__or2_1 _0541_ (.A(\comp0.B[11] ),
    .B(_0176_),
    .X(_0203_));
 sky130_fd_sc_hd__o221a_1 _0542_ (.A1(_0172_),
    .A2(net19),
    .B1(_0174_),
    .B2(net195),
    .C1(_0203_),
    .X(_0141_));
 sky130_fd_sc_hd__or2_1 _0543_ (.A(net152),
    .B(_0176_),
    .X(_0204_));
 sky130_fd_sc_hd__o221a_1 _0544_ (.A1(_0172_),
    .A2(net18),
    .B1(_0174_),
    .B2(net198),
    .C1(_0204_),
    .X(_0140_));
 sky130_fd_sc_hd__or2_1 _0545_ (.A(\comp0.B[9] ),
    .B(_0176_),
    .X(_0205_));
 sky130_fd_sc_hd__o221a_1 _0546_ (.A1(_0172_),
    .A2(net32),
    .B1(_0174_),
    .B2(net152),
    .C1(_0205_),
    .X(_0139_));
 sky130_fd_sc_hd__or2_1 _0547_ (.A(\comp0.B[8] ),
    .B(_0176_),
    .X(_0206_));
 sky130_fd_sc_hd__o221a_1 _0548_ (.A1(_0172_),
    .A2(net31),
    .B1(_0174_),
    .B2(net173),
    .C1(_0206_),
    .X(_0138_));
 sky130_fd_sc_hd__or2_1 _0549_ (.A(net171),
    .B(_0176_),
    .X(_0207_));
 sky130_fd_sc_hd__o221a_1 _0550_ (.A1(_0172_),
    .A2(net30),
    .B1(_0174_),
    .B2(net180),
    .C1(_0207_),
    .X(_0137_));
 sky130_fd_sc_hd__buf_2 _0551_ (.A(_0171_),
    .X(_0208_));
 sky130_fd_sc_hd__or2_1 _0552_ (.A(\comp0.B[6] ),
    .B(_0176_),
    .X(_0209_));
 sky130_fd_sc_hd__o221a_1 _0553_ (.A1(_0208_),
    .A2(net29),
    .B1(_0174_),
    .B2(net171),
    .C1(_0209_),
    .X(_0136_));
 sky130_fd_sc_hd__or2_1 _0554_ (.A(net160),
    .B(_0175_),
    .X(_0210_));
 sky130_fd_sc_hd__o221a_1 _0555_ (.A1(_0208_),
    .A2(net28),
    .B1(_0173_),
    .B2(net204),
    .C1(_0210_),
    .X(_0135_));
 sky130_fd_sc_hd__or2_1 _0556_ (.A(\comp0.B[4] ),
    .B(_0175_),
    .X(_0211_));
 sky130_fd_sc_hd__o221a_1 _0557_ (.A1(_0208_),
    .A2(net27),
    .B1(_0173_),
    .B2(net160),
    .C1(_0211_),
    .X(_0134_));
 sky130_fd_sc_hd__or2_1 _0558_ (.A(net185),
    .B(_0175_),
    .X(_0212_));
 sky130_fd_sc_hd__o221a_1 _0559_ (.A1(_0208_),
    .A2(net26),
    .B1(_0173_),
    .B2(net205),
    .C1(_0212_),
    .X(_0133_));
 sky130_fd_sc_hd__or2_1 _0560_ (.A(\comp0.B[2] ),
    .B(_0175_),
    .X(_0213_));
 sky130_fd_sc_hd__o221a_1 _0561_ (.A1(_0208_),
    .A2(net25),
    .B1(_0173_),
    .B2(net185),
    .C1(_0213_),
    .X(_0132_));
 sky130_fd_sc_hd__or2_1 _0562_ (.A(net201),
    .B(_0175_),
    .X(_0214_));
 sky130_fd_sc_hd__o221a_1 _0563_ (.A1(_0208_),
    .A2(net24),
    .B1(_0173_),
    .B2(net203),
    .C1(_0214_),
    .X(_0131_));
 sky130_fd_sc_hd__or2_1 _0564_ (.A(\comp0.B[0] ),
    .B(_0175_),
    .X(_0215_));
 sky130_fd_sc_hd__o221a_1 _0565_ (.A1(_0208_),
    .A2(net17),
    .B1(_0173_),
    .B2(net201),
    .C1(_0215_),
    .X(_0130_));
 sky130_fd_sc_hd__clkbuf_4 _0566_ (.A(_0182_),
    .X(_0216_));
 sky130_fd_sc_hd__a22o_1 _0567_ (.A1(net162),
    .A2(_0216_),
    .B1(_0195_),
    .B2(\acc0.A[30] ),
    .X(_0129_));
 sky130_fd_sc_hd__a22o_1 _0568_ (.A1(net208),
    .A2(_0216_),
    .B1(_0195_),
    .B2(\acc0.A[29] ),
    .X(_0128_));
 sky130_fd_sc_hd__a22o_1 _0569_ (.A1(\acc0.A[29] ),
    .A2(_0216_),
    .B1(_0195_),
    .B2(net190),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_1 _0570_ (.A1(net190),
    .A2(_0216_),
    .B1(_0195_),
    .B2(net197),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_1 _0571_ (.A1(\acc0.A[27] ),
    .A2(_0216_),
    .B1(_0195_),
    .B2(net155),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _0572_ (.A1(net155),
    .A2(_0216_),
    .B1(_0195_),
    .B2(net210),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_4 _0573_ (.A(_0178_),
    .X(_0217_));
 sky130_fd_sc_hd__a22o_1 _0574_ (.A1(\acc0.A[25] ),
    .A2(_0216_),
    .B1(_0217_),
    .B2(net199),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_1 _0575_ (.A1(net199),
    .A2(_0216_),
    .B1(_0217_),
    .B2(net215),
    .X(_0122_));
 sky130_fd_sc_hd__a22o_1 _0576_ (.A1(\acc0.A[23] ),
    .A2(_0183_),
    .B1(_0217_),
    .B2(net176),
    .X(_0121_));
 sky130_fd_sc_hd__a22o_1 _0577_ (.A1(\acc0.A[22] ),
    .A2(_0183_),
    .B1(_0217_),
    .B2(net150),
    .X(_0120_));
 sky130_fd_sc_hd__a22o_1 _0578_ (.A1(net150),
    .A2(_0183_),
    .B1(_0217_),
    .B2(net187),
    .X(_0119_));
 sky130_fd_sc_hd__a22o_1 _0579_ (.A1(net187),
    .A2(_0183_),
    .B1(_0217_),
    .B2(net211),
    .X(_0118_));
 sky130_fd_sc_hd__a22o_1 _0580_ (.A1(\acc0.A[19] ),
    .A2(_0183_),
    .B1(_0217_),
    .B2(net206),
    .X(_0117_));
 sky130_fd_sc_hd__a22o_1 _0581_ (.A1(net206),
    .A2(_0183_),
    .B1(_0217_),
    .B2(net219),
    .X(_0116_));
 sky130_fd_sc_hd__a22o_1 _0582_ (.A1(net219),
    .A2(_0183_),
    .B1(_0217_),
    .B2(net221),
    .X(_0115_));
 sky130_fd_sc_hd__a22o_1 _0583_ (.A1(\acc0.A[16] ),
    .A2(_0183_),
    .B1(_0217_),
    .B2(net165),
    .X(_0114_));
 sky130_fd_sc_hd__a22o_1 _0584_ (.A1(_0181_),
    .A2(net23),
    .B1(_0216_),
    .B2(net157),
    .X(_0113_));
 sky130_fd_sc_hd__a22o_1 _0585_ (.A1(_0181_),
    .A2(net1),
    .B1(_0216_),
    .B2(net149),
    .X(_0112_));
 sky130_fd_sc_hd__buf_2 _0586_ (.A(\control0.add ),
    .X(_0218_));
 sky130_fd_sc_hd__clkbuf_4 _0587_ (.A(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__nand2_1 _0588_ (.A(\acc0.A[30] ),
    .B(net59),
    .Y(_0220_));
 sky130_fd_sc_hd__nand2_1 _0589_ (.A(\acc0.A[28] ),
    .B(net56),
    .Y(_0221_));
 sky130_fd_sc_hd__nand2_1 _0590_ (.A(\acc0.A[22] ),
    .B(net50),
    .Y(_0222_));
 sky130_fd_sc_hd__nor2_1 _0591_ (.A(\acc0.A[23] ),
    .B(net51),
    .Y(_0223_));
 sky130_fd_sc_hd__or2_1 _0592_ (.A(\acc0.A[22] ),
    .B(net50),
    .X(_0224_));
 sky130_fd_sc_hd__nand2_1 _0593_ (.A(_0222_),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__nand2_1 _0594_ (.A(\acc0.A[20] ),
    .B(net48),
    .Y(_0226_));
 sky130_fd_sc_hd__nor2_1 _0595_ (.A(\acc0.A[21] ),
    .B(net49),
    .Y(_0227_));
 sky130_fd_sc_hd__and2_1 _0596_ (.A(\acc0.A[21] ),
    .B(net49),
    .X(_0228_));
 sky130_fd_sc_hd__inv_2 _0597_ (.A(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__o21a_1 _0598_ (.A1(_0226_),
    .A2(_0227_),
    .B1(_0229_),
    .X(_0230_));
 sky130_fd_sc_hd__nand2_1 _0599_ (.A(\acc0.A[23] ),
    .B(net51),
    .Y(_0231_));
 sky130_fd_sc_hd__o31a_1 _0600_ (.A1(_0225_),
    .A2(_0223_),
    .A3(_0230_),
    .B1(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__or2_1 _0601_ (.A(\acc0.A[23] ),
    .B(net51),
    .X(_0233_));
 sky130_fd_sc_hd__nand2_1 _0602_ (.A(_0233_),
    .B(_0231_),
    .Y(_0234_));
 sky130_fd_sc_hd__or2_1 _0603_ (.A(\acc0.A[20] ),
    .B(net48),
    .X(_0235_));
 sky130_fd_sc_hd__nand2_1 _0604_ (.A(_0226_),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__nor2_1 _0605_ (.A(_0228_),
    .B(_0227_),
    .Y(_0237_));
 sky130_fd_sc_hd__or4b_1 _0606_ (.A(_0225_),
    .B(_0234_),
    .C(_0236_),
    .D_N(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__a22o_1 _0607_ (.A1(\acc0.A[17] ),
    .A2(net44),
    .B1(net43),
    .B2(\acc0.A[16] ),
    .X(_0239_));
 sky130_fd_sc_hd__o21ai_1 _0608_ (.A1(\acc0.A[17] ),
    .A2(net44),
    .B1(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__nor2_1 _0609_ (.A(\acc0.A[19] ),
    .B(net46),
    .Y(_0241_));
 sky130_fd_sc_hd__and2_1 _0610_ (.A(\acc0.A[19] ),
    .B(net46),
    .X(_0242_));
 sky130_fd_sc_hd__or2_1 _0611_ (.A(_0241_),
    .B(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__and2_1 _0612_ (.A(\acc0.A[18] ),
    .B(net45),
    .X(_0244_));
 sky130_fd_sc_hd__nor2_1 _0613_ (.A(\acc0.A[18] ),
    .B(net45),
    .Y(_0245_));
 sky130_fd_sc_hd__or3_1 _0614_ (.A(_0243_),
    .B(_0244_),
    .C(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__nor2_1 _0615_ (.A(_0242_),
    .B(_0244_),
    .Y(_0247_));
 sky130_fd_sc_hd__o22a_1 _0616_ (.A1(_0240_),
    .A2(_0246_),
    .B1(_0247_),
    .B2(_0241_),
    .X(_0248_));
 sky130_fd_sc_hd__or2_1 _0617_ (.A(_0238_),
    .B(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__o211a_1 _0618_ (.A1(_0222_),
    .A2(_0223_),
    .B1(_0232_),
    .C1(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__or2_1 _0619_ (.A(\acc0.A[7] ),
    .B(net65),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_1 _0620_ (.A(\acc0.A[7] ),
    .B(net65),
    .Y(_0252_));
 sky130_fd_sc_hd__xor2_1 _0621_ (.A(\acc0.A[6] ),
    .B(net64),
    .X(_0253_));
 sky130_fd_sc_hd__nand3_1 _0622_ (.A(_0251_),
    .B(_0252_),
    .C(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__nor2_1 _0623_ (.A(\acc0.A[5] ),
    .B(net63),
    .Y(_0255_));
 sky130_fd_sc_hd__and2_1 _0624_ (.A(\acc0.A[4] ),
    .B(net62),
    .X(_0256_));
 sky130_fd_sc_hd__and2_1 _0625_ (.A(\acc0.A[5] ),
    .B(net63),
    .X(_0257_));
 sky130_fd_sc_hd__or2_1 _0626_ (.A(_0256_),
    .B(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__or3b_1 _0627_ (.A(_0254_),
    .B(_0255_),
    .C_N(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__nor2_1 _0628_ (.A(\acc0.A[3] ),
    .B(net61),
    .Y(_0260_));
 sky130_fd_sc_hd__and2_1 _0629_ (.A(\acc0.A[2] ),
    .B(net58),
    .X(_0261_));
 sky130_fd_sc_hd__nor2_1 _0630_ (.A(\acc0.A[2] ),
    .B(net58),
    .Y(_0262_));
 sky130_fd_sc_hd__nor2_1 _0631_ (.A(_0261_),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__nand2_1 _0632_ (.A(net149),
    .B(net36),
    .Y(_0264_));
 sky130_fd_sc_hd__nor2_1 _0633_ (.A(\acc0.A[1] ),
    .B(net47),
    .Y(_0265_));
 sky130_fd_sc_hd__nand2_1 _0634_ (.A(\acc0.A[1] ),
    .B(net47),
    .Y(_0266_));
 sky130_fd_sc_hd__o21ai_1 _0635_ (.A1(_0264_),
    .A2(_0265_),
    .B1(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__and2_1 _0636_ (.A(\acc0.A[3] ),
    .B(net61),
    .X(_0268_));
 sky130_fd_sc_hd__a211oi_1 _0637_ (.A1(_0263_),
    .A2(_0267_),
    .B1(_0268_),
    .C1(_0261_),
    .Y(_0269_));
 sky130_fd_sc_hd__nor2_1 _0638_ (.A(\acc0.A[4] ),
    .B(net62),
    .Y(_0270_));
 sky130_fd_sc_hd__nor2_1 _0639_ (.A(_0256_),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__or4b_1 _0640_ (.A(_0254_),
    .B(_0257_),
    .C(_0255_),
    .D_N(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__nand2_1 _0641_ (.A(\acc0.A[6] ),
    .B(net64),
    .Y(_0273_));
 sky130_fd_sc_hd__a21bo_1 _0642_ (.A1(_0252_),
    .A2(_0273_),
    .B1_N(_0251_),
    .X(_0274_));
 sky130_fd_sc_hd__o31a_1 _0643_ (.A1(_0260_),
    .A2(_0269_),
    .A3(_0272_),
    .B1(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__xnor2_1 _0644_ (.A(\acc0.A[15] ),
    .B(net42),
    .Y(_0276_));
 sky130_fd_sc_hd__xnor2_1 _0645_ (.A(\acc0.A[14] ),
    .B(net41),
    .Y(_0277_));
 sky130_fd_sc_hd__xnor2_1 _0646_ (.A(\acc0.A[13] ),
    .B(net40),
    .Y(_0278_));
 sky130_fd_sc_hd__xnor2_1 _0647_ (.A(\acc0.A[12] ),
    .B(net39),
    .Y(_0279_));
 sky130_fd_sc_hd__or4_1 _0648_ (.A(_0276_),
    .B(_0277_),
    .C(_0278_),
    .D(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__nand2_1 _0649_ (.A(\acc0.A[10] ),
    .B(net37),
    .Y(_0281_));
 sky130_fd_sc_hd__or2_1 _0650_ (.A(\acc0.A[10] ),
    .B(net37),
    .X(_0282_));
 sky130_fd_sc_hd__nand2_1 _0651_ (.A(_0281_),
    .B(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__nor2_1 _0652_ (.A(\acc0.A[11] ),
    .B(net38),
    .Y(_0284_));
 sky130_fd_sc_hd__nand2_1 _0653_ (.A(\acc0.A[11] ),
    .B(net38),
    .Y(_0285_));
 sky130_fd_sc_hd__and2b_1 _0654_ (.A_N(_0284_),
    .B(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__or3b_1 _0655_ (.A(_0280_),
    .B(_0283_),
    .C_N(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__and2_1 _0656_ (.A(\acc0.A[9] ),
    .B(net67),
    .X(_0288_));
 sky130_fd_sc_hd__nor2_1 _0657_ (.A(\acc0.A[9] ),
    .B(net67),
    .Y(_0289_));
 sky130_fd_sc_hd__nand2_1 _0658_ (.A(\acc0.A[8] ),
    .B(net66),
    .Y(_0290_));
 sky130_fd_sc_hd__or2_1 _0659_ (.A(\acc0.A[8] ),
    .B(net66),
    .X(_0291_));
 sky130_fd_sc_hd__nand2_1 _0660_ (.A(_0290_),
    .B(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__or4_1 _0661_ (.A(_0287_),
    .B(_0288_),
    .C(_0289_),
    .D(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__a21o_1 _0662_ (.A1(_0259_),
    .A2(_0275_),
    .B1(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__and2b_1 _0663_ (.A_N(_0288_),
    .B(_0290_),
    .X(_0295_));
 sky130_fd_sc_hd__o21a_1 _0664_ (.A1(_0281_),
    .A2(_0284_),
    .B1(_0285_),
    .X(_0296_));
 sky130_fd_sc_hd__nor2_1 _0665_ (.A(\acc0.A[13] ),
    .B(net40),
    .Y(_0297_));
 sky130_fd_sc_hd__nand2_1 _0666_ (.A(\acc0.A[12] ),
    .B(net39),
    .Y(_0298_));
 sky130_fd_sc_hd__nand2_1 _0667_ (.A(\acc0.A[13] ),
    .B(net40),
    .Y(_0299_));
 sky130_fd_sc_hd__o21a_1 _0668_ (.A1(_0297_),
    .A2(_0298_),
    .B1(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__or3_1 _0669_ (.A(_0276_),
    .B(_0277_),
    .C(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__o211a_1 _0670_ (.A1(\acc0.A[15] ),
    .A2(net42),
    .B1(net41),
    .C1(\acc0.A[14] ),
    .X(_0302_));
 sky130_fd_sc_hd__a21oi_1 _0671_ (.A1(\acc0.A[15] ),
    .A2(net42),
    .B1(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__o211a_1 _0672_ (.A1(_0280_),
    .A2(_0296_),
    .B1(_0301_),
    .C1(_0303_),
    .X(_0304_));
 sky130_fd_sc_hd__o31a_1 _0673_ (.A1(_0287_),
    .A2(_0289_),
    .A3(_0295_),
    .B1(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__nand2_1 _0674_ (.A(\acc0.A[16] ),
    .B(net43),
    .Y(_0306_));
 sky130_fd_sc_hd__or2_1 _0675_ (.A(\acc0.A[16] ),
    .B(net43),
    .X(_0307_));
 sky130_fd_sc_hd__nand2_1 _0676_ (.A(_0306_),
    .B(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__xnor2_1 _0677_ (.A(\acc0.A[17] ),
    .B(net44),
    .Y(_0309_));
 sky130_fd_sc_hd__or2_1 _0678_ (.A(_0308_),
    .B(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__or2_1 _0679_ (.A(_0246_),
    .B(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__a211o_1 _0680_ (.A1(_0294_),
    .A2(_0305_),
    .B1(_0311_),
    .C1(_0238_),
    .X(_0312_));
 sky130_fd_sc_hd__nand2_1 _0681_ (.A(\acc0.A[25] ),
    .B(net53),
    .Y(_0313_));
 sky130_fd_sc_hd__or2_1 _0682_ (.A(\acc0.A[25] ),
    .B(net53),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _0683_ (.A(_0313_),
    .B(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__and2_1 _0684_ (.A(\acc0.A[27] ),
    .B(net55),
    .X(_0316_));
 sky130_fd_sc_hd__or2_1 _0685_ (.A(\acc0.A[27] ),
    .B(net55),
    .X(_0317_));
 sky130_fd_sc_hd__or2b_1 _0686_ (.A(_0316_),
    .B_N(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__and2_1 _0687_ (.A(\acc0.A[26] ),
    .B(net54),
    .X(_0319_));
 sky130_fd_sc_hd__nor2_1 _0688_ (.A(\acc0.A[26] ),
    .B(net54),
    .Y(_0320_));
 sky130_fd_sc_hd__or2_1 _0689_ (.A(_0319_),
    .B(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__or2_1 _0690_ (.A(_0318_),
    .B(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _0691_ (.A(_0315_),
    .B(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__nand2_1 _0692_ (.A(\acc0.A[24] ),
    .B(net52),
    .Y(_0324_));
 sky130_fd_sc_hd__or2_1 _0693_ (.A(\acc0.A[24] ),
    .B(net52),
    .X(_0325_));
 sky130_fd_sc_hd__nand2_1 _0694_ (.A(_0324_),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__a211o_1 _0695_ (.A1(_0250_),
    .A2(_0312_),
    .B1(_0323_),
    .C1(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__nor2_1 _0696_ (.A(\acc0.A[25] ),
    .B(net53),
    .Y(_0328_));
 sky130_fd_sc_hd__a211o_1 _0697_ (.A1(_0324_),
    .A2(_0313_),
    .B1(_0328_),
    .C1(_0322_),
    .X(_0329_));
 sky130_fd_sc_hd__a21oi_1 _0698_ (.A1(_0317_),
    .A2(_0319_),
    .B1(_0316_),
    .Y(_0330_));
 sky130_fd_sc_hd__or2_1 _0699_ (.A(\acc0.A[28] ),
    .B(net56),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_1 _0700_ (.A(_0221_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__a31o_1 _0701_ (.A1(_0327_),
    .A2(_0329_),
    .A3(_0330_),
    .B1(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__nand2_1 _0702_ (.A(\acc0.A[29] ),
    .B(net57),
    .Y(_0334_));
 sky130_fd_sc_hd__nor2_1 _0703_ (.A(\acc0.A[29] ),
    .B(net57),
    .Y(_0335_));
 sky130_fd_sc_hd__or2_1 _0704_ (.A(\acc0.A[30] ),
    .B(net59),
    .X(_0336_));
 sky130_fd_sc_hd__and2_1 _0705_ (.A(_0220_),
    .B(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__inv_2 _0706_ (.A(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__a311o_1 _0707_ (.A1(_0221_),
    .A2(_0333_),
    .A3(_0334_),
    .B1(_0335_),
    .C1(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__or2_1 _0708_ (.A(\acc0.A[31] ),
    .B(net60),
    .X(_0340_));
 sky130_fd_sc_hd__nand2_1 _0709_ (.A(\acc0.A[31] ),
    .B(net60),
    .Y(_0341_));
 sky130_fd_sc_hd__a22oi_1 _0710_ (.A1(_0220_),
    .A2(_0339_),
    .B1(_0340_),
    .B2(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_2 _0711_ (.A(\control0.add ),
    .Y(_0343_));
 sky130_fd_sc_hd__a41o_1 _0712_ (.A1(_0220_),
    .A2(_0339_),
    .A3(_0340_),
    .A4(_0341_),
    .B1(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_4 _0713_ (.A(_0208_),
    .X(_0345_));
 sky130_fd_sc_hd__o221a_1 _0714_ (.A1(net225),
    .A2(_0219_),
    .B1(_0342_),
    .B2(_0344_),
    .C1(_0345_),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_4 _0715_ (.A(_0343_),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_4 _0716_ (.A(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__a31o_1 _0717_ (.A1(_0221_),
    .A2(_0333_),
    .A3(_0334_),
    .B1(_0335_),
    .X(_0348_));
 sky130_fd_sc_hd__xnor2_1 _0718_ (.A(_0337_),
    .B(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__buf_2 _0719_ (.A(\control0.add ),
    .X(_0350_));
 sky130_fd_sc_hd__or2_1 _0720_ (.A(_0350_),
    .B(net239),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_4 _0721_ (.A(_0208_),
    .X(_0352_));
 sky130_fd_sc_hd__o211a_1 _0722_ (.A1(_0347_),
    .A2(_0349_),
    .B1(_0351_),
    .C1(_0352_),
    .X(_0110_));
 sky130_fd_sc_hd__and2b_1 _0723_ (.A_N(_0335_),
    .B(_0334_),
    .X(_0353_));
 sky130_fd_sc_hd__a21oi_1 _0724_ (.A1(_0221_),
    .A2(_0333_),
    .B1(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__a31o_1 _0725_ (.A1(_0221_),
    .A2(_0333_),
    .A3(_0353_),
    .B1(_0343_),
    .X(_0355_));
 sky130_fd_sc_hd__o221a_1 _0726_ (.A1(_0219_),
    .A2(net227),
    .B1(_0354_),
    .B2(_0355_),
    .C1(_0345_),
    .X(_0109_));
 sky130_fd_sc_hd__nand4_1 _0727_ (.A(_0332_),
    .B(_0327_),
    .C(_0329_),
    .D(_0330_),
    .Y(_0356_));
 sky130_fd_sc_hd__and2_1 _0728_ (.A(_0333_),
    .B(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__or2_1 _0729_ (.A(_0350_),
    .B(net242),
    .X(_0358_));
 sky130_fd_sc_hd__o211a_1 _0730_ (.A1(_0347_),
    .A2(_0357_),
    .B1(_0358_),
    .C1(_0352_),
    .X(_0108_));
 sky130_fd_sc_hd__a21o_1 _0731_ (.A1(_0250_),
    .A2(_0312_),
    .B1(_0326_),
    .X(_0359_));
 sky130_fd_sc_hd__a31o_1 _0732_ (.A1(_0324_),
    .A2(_0359_),
    .A3(_0313_),
    .B1(_0328_),
    .X(_0360_));
 sky130_fd_sc_hd__o21ba_1 _0733_ (.A1(_0321_),
    .A2(_0360_),
    .B1_N(_0319_),
    .X(_0361_));
 sky130_fd_sc_hd__xnor2_1 _0734_ (.A(_0318_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__nor2_1 _0735_ (.A(_0350_),
    .B(net224),
    .Y(_0363_));
 sky130_fd_sc_hd__a211oi_1 _0736_ (.A1(_0219_),
    .A2(_0362_),
    .B1(_0363_),
    .C1(_0181_),
    .Y(_0107_));
 sky130_fd_sc_hd__xor2_1 _0737_ (.A(_0321_),
    .B(_0360_),
    .X(_0364_));
 sky130_fd_sc_hd__or2_1 _0738_ (.A(_0350_),
    .B(net244),
    .X(_0365_));
 sky130_fd_sc_hd__o211a_1 _0739_ (.A1(_0347_),
    .A2(_0364_),
    .B1(_0365_),
    .C1(_0352_),
    .X(_0106_));
 sky130_fd_sc_hd__nand2_1 _0740_ (.A(_0324_),
    .B(_0359_),
    .Y(_0366_));
 sky130_fd_sc_hd__nor2_1 _0741_ (.A(_0315_),
    .B(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__a21o_1 _0742_ (.A1(_0315_),
    .A2(_0366_),
    .B1(_0343_),
    .X(_0368_));
 sky130_fd_sc_hd__o221a_1 _0743_ (.A1(_0219_),
    .A2(net237),
    .B1(_0367_),
    .B2(_0368_),
    .C1(_0345_),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_4 _0744_ (.A(_0350_),
    .X(_0369_));
 sky130_fd_sc_hd__nand3_1 _0745_ (.A(_0326_),
    .B(_0250_),
    .C(_0312_),
    .Y(_0370_));
 sky130_fd_sc_hd__a21o_1 _0746_ (.A1(_0359_),
    .A2(_0370_),
    .B1(_0346_),
    .X(_0371_));
 sky130_fd_sc_hd__o211a_1 _0747_ (.A1(_0369_),
    .A2(net216),
    .B1(_0371_),
    .C1(_0352_),
    .X(_0104_));
 sky130_fd_sc_hd__a21o_1 _0748_ (.A1(_0294_),
    .A2(_0305_),
    .B1(_0311_),
    .X(_0372_));
 sky130_fd_sc_hd__a21o_1 _0749_ (.A1(_0248_),
    .A2(_0372_),
    .B1(_0236_),
    .X(_0373_));
 sky130_fd_sc_hd__and3_1 _0750_ (.A(_0226_),
    .B(_0229_),
    .C(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__or3_1 _0751_ (.A(_0225_),
    .B(_0227_),
    .C(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__a21boi_1 _0752_ (.A1(_0222_),
    .A2(_0375_),
    .B1_N(_0234_),
    .Y(_0376_));
 sky130_fd_sc_hd__a41o_1 _0753_ (.A1(_0222_),
    .A2(_0233_),
    .A3(_0231_),
    .A4(_0375_),
    .B1(_0343_),
    .X(_0377_));
 sky130_fd_sc_hd__o221a_1 _0754_ (.A1(_0219_),
    .A2(net241),
    .B1(_0376_),
    .B2(_0377_),
    .C1(_0345_),
    .X(_0103_));
 sky130_fd_sc_hd__nor2_1 _0755_ (.A(_0227_),
    .B(_0374_),
    .Y(_0378_));
 sky130_fd_sc_hd__xnor2_1 _0756_ (.A(_0225_),
    .B(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__or2_1 _0757_ (.A(_0350_),
    .B(net243),
    .X(_0380_));
 sky130_fd_sc_hd__o211a_1 _0758_ (.A1(_0347_),
    .A2(_0379_),
    .B1(_0380_),
    .C1(_0352_),
    .X(_0102_));
 sky130_fd_sc_hd__nand2_1 _0759_ (.A(_0226_),
    .B(_0373_),
    .Y(_0381_));
 sky130_fd_sc_hd__xnor2_1 _0760_ (.A(_0237_),
    .B(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__nand2_1 _0761_ (.A(_0219_),
    .B(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__o211a_1 _0762_ (.A1(_0369_),
    .A2(net213),
    .B1(_0383_),
    .C1(_0352_),
    .X(_0101_));
 sky130_fd_sc_hd__nand3_1 _0763_ (.A(_0236_),
    .B(_0248_),
    .C(_0372_),
    .Y(_0384_));
 sky130_fd_sc_hd__a21o_1 _0764_ (.A1(_0373_),
    .A2(_0384_),
    .B1(_0346_),
    .X(_0385_));
 sky130_fd_sc_hd__o211a_1 _0765_ (.A1(_0369_),
    .A2(net220),
    .B1(_0385_),
    .C1(_0352_),
    .X(_0100_));
 sky130_fd_sc_hd__nor2_1 _0766_ (.A(_0244_),
    .B(_0245_),
    .Y(_0386_));
 sky130_fd_sc_hd__and2_1 _0767_ (.A(_0294_),
    .B(_0305_),
    .X(_0387_));
 sky130_fd_sc_hd__o21ai_1 _0768_ (.A1(_0387_),
    .A2(_0310_),
    .B1(_0240_),
    .Y(_0388_));
 sky130_fd_sc_hd__a21o_1 _0769_ (.A1(_0386_),
    .A2(_0388_),
    .B1(_0244_),
    .X(_0389_));
 sky130_fd_sc_hd__o21a_1 _0770_ (.A1(_0243_),
    .A2(_0389_),
    .B1(\control0.add ),
    .X(_0390_));
 sky130_fd_sc_hd__a21bo_1 _0771_ (.A1(_0243_),
    .A2(_0389_),
    .B1_N(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__o211a_1 _0772_ (.A1(_0369_),
    .A2(net223),
    .B1(_0391_),
    .C1(_0352_),
    .X(_0099_));
 sky130_fd_sc_hd__xor2_1 _0773_ (.A(_0386_),
    .B(_0388_),
    .X(_0392_));
 sky130_fd_sc_hd__or2_1 _0774_ (.A(_0218_),
    .B(net45),
    .X(_0393_));
 sky130_fd_sc_hd__o211a_1 _0775_ (.A1(_0347_),
    .A2(_0392_),
    .B1(_0393_),
    .C1(_0352_),
    .X(_0098_));
 sky130_fd_sc_hd__o21ai_1 _0776_ (.A1(_0387_),
    .A2(_0308_),
    .B1(_0306_),
    .Y(_0394_));
 sky130_fd_sc_hd__xnor2_1 _0777_ (.A(_0309_),
    .B(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__or2_1 _0778_ (.A(_0218_),
    .B(net44),
    .X(_0396_));
 sky130_fd_sc_hd__o211a_1 _0779_ (.A1(_0347_),
    .A2(_0395_),
    .B1(_0396_),
    .C1(_0352_),
    .X(_0097_));
 sky130_fd_sc_hd__xor2_1 _0780_ (.A(_0387_),
    .B(_0308_),
    .X(_0397_));
 sky130_fd_sc_hd__or2_1 _0781_ (.A(_0218_),
    .B(net43),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_4 _0782_ (.A(_0208_),
    .X(_0399_));
 sky130_fd_sc_hd__o211a_1 _0783_ (.A1(_0347_),
    .A2(_0397_),
    .B1(_0398_),
    .C1(_0399_),
    .X(_0096_));
 sky130_fd_sc_hd__nand2_1 _0784_ (.A(\acc0.A[14] ),
    .B(net41),
    .Y(_0400_));
 sky130_fd_sc_hd__a21o_1 _0785_ (.A1(_0259_),
    .A2(_0275_),
    .B1(_0292_),
    .X(_0401_));
 sky130_fd_sc_hd__a211o_1 _0786_ (.A1(_0295_),
    .A2(_0401_),
    .B1(_0283_),
    .C1(_0289_),
    .X(_0402_));
 sky130_fd_sc_hd__a31o_1 _0787_ (.A1(_0281_),
    .A2(_0285_),
    .A3(_0402_),
    .B1(_0284_),
    .X(_0403_));
 sky130_fd_sc_hd__or2_1 _0788_ (.A(_0279_),
    .B(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__a311o_1 _0789_ (.A1(_0299_),
    .A2(_0298_),
    .A3(_0404_),
    .B1(_0297_),
    .C1(_0277_),
    .X(_0405_));
 sky130_fd_sc_hd__xor2_1 _0790_ (.A(\acc0.A[15] ),
    .B(net42),
    .X(_0406_));
 sky130_fd_sc_hd__a21oi_1 _0791_ (.A1(_0400_),
    .A2(_0405_),
    .B1(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__a31o_1 _0792_ (.A1(_0406_),
    .A2(_0400_),
    .A3(_0405_),
    .B1(_0343_),
    .X(_0408_));
 sky130_fd_sc_hd__o221a_1 _0793_ (.A1(_0219_),
    .A2(net42),
    .B1(_0407_),
    .B2(_0408_),
    .C1(_0345_),
    .X(_0095_));
 sky130_fd_sc_hd__o211ai_1 _0794_ (.A1(_0297_),
    .A2(_0404_),
    .B1(_0300_),
    .C1(_0277_),
    .Y(_0409_));
 sky130_fd_sc_hd__a21o_1 _0795_ (.A1(_0405_),
    .A2(_0409_),
    .B1(_0346_),
    .X(_0410_));
 sky130_fd_sc_hd__o211a_1 _0796_ (.A1(_0369_),
    .A2(net238),
    .B1(_0410_),
    .C1(_0399_),
    .X(_0094_));
 sky130_fd_sc_hd__and2b_1 _0797_ (.A_N(_0297_),
    .B(_0299_),
    .X(_0411_));
 sky130_fd_sc_hd__a21oi_1 _0798_ (.A1(_0298_),
    .A2(_0404_),
    .B1(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__a31o_1 _0799_ (.A1(_0411_),
    .A2(_0298_),
    .A3(_0404_),
    .B1(_0343_),
    .X(_0413_));
 sky130_fd_sc_hd__o221a_1 _0800_ (.A1(_0219_),
    .A2(net245),
    .B1(_0412_),
    .B2(_0413_),
    .C1(_0345_),
    .X(_0093_));
 sky130_fd_sc_hd__nand2_1 _0801_ (.A(_0279_),
    .B(_0403_),
    .Y(_0414_));
 sky130_fd_sc_hd__and2_1 _0802_ (.A(_0404_),
    .B(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__or2_1 _0803_ (.A(_0218_),
    .B(net39),
    .X(_0416_));
 sky130_fd_sc_hd__o211a_1 _0804_ (.A1(_0347_),
    .A2(_0415_),
    .B1(_0416_),
    .C1(_0399_),
    .X(_0092_));
 sky130_fd_sc_hd__and3_1 _0805_ (.A(_0281_),
    .B(_0286_),
    .C(_0402_),
    .X(_0417_));
 sky130_fd_sc_hd__a21oi_1 _0806_ (.A1(_0281_),
    .A2(_0402_),
    .B1(_0286_),
    .Y(_0418_));
 sky130_fd_sc_hd__or2_1 _0807_ (.A(_0218_),
    .B(net246),
    .X(_0419_));
 sky130_fd_sc_hd__o311a_1 _0808_ (.A1(_0346_),
    .A2(_0417_),
    .A3(_0418_),
    .B1(_0419_),
    .C1(_0345_),
    .X(_0091_));
 sky130_fd_sc_hd__a21o_1 _0809_ (.A1(_0295_),
    .A2(_0401_),
    .B1(_0289_),
    .X(_0420_));
 sky130_fd_sc_hd__nand2_1 _0810_ (.A(_0283_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__a21o_1 _0811_ (.A1(_0402_),
    .A2(_0421_),
    .B1(_0346_),
    .X(_0422_));
 sky130_fd_sc_hd__o211a_1 _0812_ (.A1(_0369_),
    .A2(net217),
    .B1(_0422_),
    .C1(_0399_),
    .X(_0090_));
 sky130_fd_sc_hd__nor2_1 _0813_ (.A(_0288_),
    .B(_0289_),
    .Y(_0423_));
 sky130_fd_sc_hd__and3_1 _0814_ (.A(_0423_),
    .B(_0290_),
    .C(_0401_),
    .X(_0424_));
 sky130_fd_sc_hd__a21oi_1 _0815_ (.A1(_0290_),
    .A2(_0401_),
    .B1(_0423_),
    .Y(_0425_));
 sky130_fd_sc_hd__or2_1 _0816_ (.A(_0218_),
    .B(net67),
    .X(_0426_));
 sky130_fd_sc_hd__o311a_1 _0817_ (.A1(_0346_),
    .A2(_0424_),
    .A3(_0425_),
    .B1(_0426_),
    .C1(_0345_),
    .X(_0089_));
 sky130_fd_sc_hd__nand3_1 _0818_ (.A(_0259_),
    .B(_0275_),
    .C(_0292_),
    .Y(_0427_));
 sky130_fd_sc_hd__a21o_1 _0819_ (.A1(_0401_),
    .A2(_0427_),
    .B1(_0346_),
    .X(_0428_));
 sky130_fd_sc_hd__o211a_1 _0820_ (.A1(_0369_),
    .A2(net214),
    .B1(_0428_),
    .C1(_0399_),
    .X(_0088_));
 sky130_fd_sc_hd__nand2_1 _0821_ (.A(_0251_),
    .B(_0252_),
    .Y(_0429_));
 sky130_fd_sc_hd__nor2_1 _0822_ (.A(\acc0.A[6] ),
    .B(net64),
    .Y(_0430_));
 sky130_fd_sc_hd__nor2_1 _0823_ (.A(_0260_),
    .B(_0269_),
    .Y(_0431_));
 sky130_fd_sc_hd__and2_1 _0824_ (.A(_0431_),
    .B(_0271_),
    .X(_0432_));
 sky130_fd_sc_hd__or2_1 _0825_ (.A(_0258_),
    .B(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__or2b_1 _0826_ (.A(_0255_),
    .B_N(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__o21ai_1 _0827_ (.A1(_0430_),
    .A2(_0434_),
    .B1(_0273_),
    .Y(_0435_));
 sky130_fd_sc_hd__a21oi_1 _0828_ (.A1(_0429_),
    .A2(_0435_),
    .B1(_0343_),
    .Y(_0436_));
 sky130_fd_sc_hd__o21ai_1 _0829_ (.A1(_0429_),
    .A2(_0435_),
    .B1(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__o211a_1 _0830_ (.A1(_0369_),
    .A2(net212),
    .B1(_0437_),
    .C1(_0399_),
    .X(_0087_));
 sky130_fd_sc_hd__xor2_1 _0831_ (.A(_0253_),
    .B(_0434_),
    .X(_0438_));
 sky130_fd_sc_hd__nand2_1 _0832_ (.A(_0350_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__o211a_1 _0833_ (.A1(_0369_),
    .A2(net235),
    .B1(_0439_),
    .C1(_0399_),
    .X(_0086_));
 sky130_fd_sc_hd__nor2_1 _0834_ (.A(_0255_),
    .B(_0433_),
    .Y(_0440_));
 sky130_fd_sc_hd__o22a_1 _0835_ (.A1(_0257_),
    .A2(_0255_),
    .B1(_0432_),
    .B2(_0256_),
    .X(_0441_));
 sky130_fd_sc_hd__or2_1 _0836_ (.A(_0218_),
    .B(net248),
    .X(_0442_));
 sky130_fd_sc_hd__o311a_1 _0837_ (.A1(_0346_),
    .A2(_0440_),
    .A3(_0441_),
    .B1(_0442_),
    .C1(_0172_),
    .X(_0085_));
 sky130_fd_sc_hd__nor2_1 _0838_ (.A(_0431_),
    .B(_0271_),
    .Y(_0443_));
 sky130_fd_sc_hd__nor2_1 _0839_ (.A(_0432_),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__or2_1 _0840_ (.A(_0218_),
    .B(net62),
    .X(_0445_));
 sky130_fd_sc_hd__o211a_1 _0841_ (.A1(_0347_),
    .A2(_0444_),
    .B1(_0445_),
    .C1(_0399_),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _0842_ (.A(_0263_),
    .B(_0267_),
    .X(_0446_));
 sky130_fd_sc_hd__or2_1 _0843_ (.A(_0260_),
    .B(_0268_),
    .X(_0447_));
 sky130_fd_sc_hd__o21a_1 _0844_ (.A1(_0261_),
    .A2(_0446_),
    .B1(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__o31ai_1 _0845_ (.A1(_0261_),
    .A2(_0446_),
    .A3(_0447_),
    .B1(_0350_),
    .Y(_0449_));
 sky130_fd_sc_hd__o221a_1 _0846_ (.A1(_0219_),
    .A2(net233),
    .B1(_0448_),
    .B2(_0449_),
    .C1(_0345_),
    .X(_0083_));
 sky130_fd_sc_hd__nor2_1 _0847_ (.A(_0263_),
    .B(_0267_),
    .Y(_0450_));
 sky130_fd_sc_hd__o21ai_1 _0848_ (.A1(_0446_),
    .A2(_0450_),
    .B1(_0350_),
    .Y(_0451_));
 sky130_fd_sc_hd__o211a_1 _0849_ (.A1(_0219_),
    .A2(net222),
    .B1(_0451_),
    .C1(_0399_),
    .X(_0082_));
 sky130_fd_sc_hd__or2_1 _0850_ (.A(\acc0.A[1] ),
    .B(net47),
    .X(_0452_));
 sky130_fd_sc_hd__nand2_1 _0851_ (.A(_0266_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__xor2_1 _0852_ (.A(_0264_),
    .B(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__or2_1 _0853_ (.A(_0218_),
    .B(net47),
    .X(_0455_));
 sky130_fd_sc_hd__o211a_1 _0854_ (.A1(_0347_),
    .A2(_0454_),
    .B1(_0455_),
    .C1(_0399_),
    .X(_0081_));
 sky130_fd_sc_hd__a21o_1 _0855_ (.A1(net149),
    .A2(_0350_),
    .B1(net234),
    .X(_0456_));
 sky130_fd_sc_hd__o211a_1 _0856_ (.A1(_0346_),
    .A2(_0264_),
    .B1(_0456_),
    .C1(_0345_),
    .X(_0080_));
 sky130_fd_sc_hd__buf_1 _0857_ (.A(clknet_1_1__leaf_clk),
    .X(_0457_));
 sky130_fd_sc_hd__buf_1 _0858_ (.A(clknet_1_1__leaf__0457_),
    .X(_0458_));
 sky130_fd_sc_hd__inv_2 _0859__1 (.A(clknet_1_0__leaf__0458_),
    .Y(net68));
 sky130_fd_sc_hd__inv_2 _0860__2 (.A(clknet_1_0__leaf__0458_),
    .Y(net69));
 sky130_fd_sc_hd__inv_2 _0861__3 (.A(clknet_1_0__leaf__0458_),
    .Y(net70));
 sky130_fd_sc_hd__inv_2 _0862__4 (.A(clknet_1_0__leaf__0458_),
    .Y(net71));
 sky130_fd_sc_hd__inv_2 _0863__5 (.A(clknet_1_1__leaf__0458_),
    .Y(net72));
 sky130_fd_sc_hd__inv_2 _0864__6 (.A(clknet_1_1__leaf__0458_),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _0865__7 (.A(clknet_1_1__leaf__0458_),
    .Y(net74));
 sky130_fd_sc_hd__inv_2 _0866__8 (.A(clknet_1_1__leaf__0458_),
    .Y(net75));
 sky130_fd_sc_hd__inv_2 _0867__9 (.A(clknet_1_1__leaf__0458_),
    .Y(net76));
 sky130_fd_sc_hd__inv_2 _0868__10 (.A(clknet_1_0__leaf__0458_),
    .Y(net77));
 sky130_fd_sc_hd__buf_1 _0869_ (.A(clknet_1_0__leaf__0457_),
    .X(_0459_));
 sky130_fd_sc_hd__inv_2 _0870__11 (.A(clknet_1_1__leaf__0459_),
    .Y(net78));
 sky130_fd_sc_hd__inv_2 _0871__12 (.A(clknet_1_1__leaf__0459_),
    .Y(net79));
 sky130_fd_sc_hd__inv_2 _0872__13 (.A(clknet_1_1__leaf__0459_),
    .Y(net80));
 sky130_fd_sc_hd__inv_2 _0873__14 (.A(clknet_1_1__leaf__0459_),
    .Y(net81));
 sky130_fd_sc_hd__inv_2 _0874__15 (.A(clknet_1_0__leaf__0459_),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _0875__16 (.A(clknet_1_1__leaf__0459_),
    .Y(net83));
 sky130_fd_sc_hd__inv_2 _0876__17 (.A(clknet_1_0__leaf__0459_),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _0877__18 (.A(clknet_1_1__leaf__0459_),
    .Y(net85));
 sky130_fd_sc_hd__inv_2 _0878__19 (.A(clknet_1_0__leaf__0459_),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 _0879__20 (.A(clknet_1_0__leaf__0459_),
    .Y(net87));
 sky130_fd_sc_hd__buf_1 _0880_ (.A(clknet_1_0__leaf__0457_),
    .X(_0460_));
 sky130_fd_sc_hd__inv_2 _0881__21 (.A(clknet_1_0__leaf__0460_),
    .Y(net88));
 sky130_fd_sc_hd__inv_2 _0882__22 (.A(clknet_1_0__leaf__0460_),
    .Y(net89));
 sky130_fd_sc_hd__inv_2 _0883__23 (.A(clknet_1_0__leaf__0460_),
    .Y(net90));
 sky130_fd_sc_hd__inv_2 _0884__24 (.A(clknet_1_0__leaf__0460_),
    .Y(net91));
 sky130_fd_sc_hd__inv_2 _0885__25 (.A(clknet_1_0__leaf__0460_),
    .Y(net92));
 sky130_fd_sc_hd__inv_2 _0886__26 (.A(clknet_1_1__leaf__0460_),
    .Y(net93));
 sky130_fd_sc_hd__inv_2 _0887__27 (.A(clknet_1_1__leaf__0460_),
    .Y(net94));
 sky130_fd_sc_hd__inv_2 _0888__28 (.A(clknet_1_1__leaf__0460_),
    .Y(net95));
 sky130_fd_sc_hd__inv_2 _0889__29 (.A(clknet_1_1__leaf__0460_),
    .Y(net96));
 sky130_fd_sc_hd__inv_2 _0890__30 (.A(clknet_1_1__leaf__0460_),
    .Y(net97));
 sky130_fd_sc_hd__buf_1 _0891_ (.A(clknet_1_0__leaf__0457_),
    .X(_0461_));
 sky130_fd_sc_hd__inv_2 _0892__31 (.A(clknet_1_1__leaf__0461_),
    .Y(net98));
 sky130_fd_sc_hd__inv_2 _0893__32 (.A(clknet_1_1__leaf__0461_),
    .Y(net99));
 sky130_fd_sc_hd__inv_2 _0894__33 (.A(clknet_1_0__leaf__0461_),
    .Y(net100));
 sky130_fd_sc_hd__inv_2 _0895__34 (.A(clknet_1_0__leaf__0461_),
    .Y(net101));
 sky130_fd_sc_hd__inv_2 _0896__35 (.A(clknet_1_1__leaf__0461_),
    .Y(net102));
 sky130_fd_sc_hd__inv_2 _0897__36 (.A(clknet_1_1__leaf__0461_),
    .Y(net103));
 sky130_fd_sc_hd__inv_2 _0898__37 (.A(clknet_1_0__leaf__0461_),
    .Y(net104));
 sky130_fd_sc_hd__inv_2 _0899__38 (.A(clknet_1_0__leaf__0461_),
    .Y(net105));
 sky130_fd_sc_hd__inv_2 _0900__39 (.A(clknet_1_0__leaf__0461_),
    .Y(net106));
 sky130_fd_sc_hd__inv_2 _0901__40 (.A(clknet_1_0__leaf__0461_),
    .Y(net107));
 sky130_fd_sc_hd__buf_1 _0902_ (.A(clknet_1_0__leaf__0457_),
    .X(_0462_));
 sky130_fd_sc_hd__inv_2 _0903__41 (.A(clknet_1_0__leaf__0462_),
    .Y(net108));
 sky130_fd_sc_hd__inv_2 _0904__42 (.A(clknet_1_0__leaf__0462_),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _0905__43 (.A(clknet_1_0__leaf__0462_),
    .Y(net110));
 sky130_fd_sc_hd__inv_2 _0906__44 (.A(clknet_1_0__leaf__0462_),
    .Y(net111));
 sky130_fd_sc_hd__inv_2 _0907__45 (.A(clknet_1_0__leaf__0462_),
    .Y(net112));
 sky130_fd_sc_hd__inv_2 _0908__46 (.A(clknet_1_1__leaf__0462_),
    .Y(net113));
 sky130_fd_sc_hd__inv_2 _0909__47 (.A(clknet_1_1__leaf__0462_),
    .Y(net114));
 sky130_fd_sc_hd__inv_2 _0910__48 (.A(clknet_1_1__leaf__0462_),
    .Y(net115));
 sky130_fd_sc_hd__inv_2 _0911__49 (.A(clknet_1_1__leaf__0462_),
    .Y(net116));
 sky130_fd_sc_hd__inv_2 _0912__50 (.A(clknet_1_1__leaf__0462_),
    .Y(net117));
 sky130_fd_sc_hd__buf_1 _0913_ (.A(clknet_1_1__leaf__0457_),
    .X(_0463_));
 sky130_fd_sc_hd__inv_2 _0914__51 (.A(clknet_1_1__leaf__0463_),
    .Y(net118));
 sky130_fd_sc_hd__inv_2 _0915__52 (.A(clknet_1_1__leaf__0463_),
    .Y(net119));
 sky130_fd_sc_hd__inv_2 _0916__53 (.A(clknet_1_1__leaf__0463_),
    .Y(net120));
 sky130_fd_sc_hd__inv_2 _0917__54 (.A(clknet_1_1__leaf__0463_),
    .Y(net121));
 sky130_fd_sc_hd__inv_2 _0918__55 (.A(clknet_1_1__leaf__0463_),
    .Y(net122));
 sky130_fd_sc_hd__inv_2 _0919__56 (.A(clknet_1_0__leaf__0463_),
    .Y(net123));
 sky130_fd_sc_hd__inv_2 _0920__57 (.A(clknet_1_0__leaf__0463_),
    .Y(net124));
 sky130_fd_sc_hd__inv_2 _0921__58 (.A(clknet_1_0__leaf__0463_),
    .Y(net125));
 sky130_fd_sc_hd__inv_2 _0922__59 (.A(clknet_1_0__leaf__0463_),
    .Y(net126));
 sky130_fd_sc_hd__inv_2 _0923__60 (.A(clknet_1_0__leaf__0463_),
    .Y(net127));
 sky130_fd_sc_hd__buf_1 _0924_ (.A(clknet_1_1__leaf__0457_),
    .X(_0464_));
 sky130_fd_sc_hd__inv_2 _0925__61 (.A(clknet_1_1__leaf__0464_),
    .Y(net128));
 sky130_fd_sc_hd__inv_2 _0926__62 (.A(clknet_1_1__leaf__0464_),
    .Y(net129));
 sky130_fd_sc_hd__inv_2 _0927__63 (.A(clknet_1_1__leaf__0464_),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _0928__64 (.A(clknet_1_1__leaf__0464_),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _0929__65 (.A(clknet_1_1__leaf__0464_),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _0930__66 (.A(clknet_1_0__leaf__0464_),
    .Y(net133));
 sky130_fd_sc_hd__inv_2 _0931__67 (.A(clknet_1_0__leaf__0464_),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _0932__68 (.A(clknet_1_0__leaf__0464_),
    .Y(net135));
 sky130_fd_sc_hd__inv_2 _0933__69 (.A(clknet_1_0__leaf__0464_),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _0934__70 (.A(clknet_1_1__leaf__0464_),
    .Y(net137));
 sky130_fd_sc_hd__buf_1 _0935_ (.A(clknet_1_1__leaf__0457_),
    .X(_0465_));
 sky130_fd_sc_hd__inv_2 _0936__71 (.A(clknet_1_0__leaf__0465_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _0937__72 (.A(clknet_1_0__leaf__0465_),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _0938__73 (.A(clknet_1_0__leaf__0465_),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _0939__74 (.A(clknet_1_1__leaf__0465_),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _0940__75 (.A(clknet_1_1__leaf__0465_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _0941__76 (.A(clknet_1_1__leaf__0465_),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _0942__77 (.A(clknet_1_1__leaf__0465_),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _0943__78 (.A(clknet_1_1__leaf__0465_),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _0944__79 (.A(clknet_1_1__leaf__0465_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _0945__80 (.A(clknet_1_0__leaf__0465_),
    .Y(net147));
 sky130_fd_sc_hd__or3_2 _0946_ (.A(net34),
    .B(\control0.state[1] ),
    .C(\control0.state[0] ),
    .X(_0466_));
 sky130_fd_sc_hd__nor2_1 _0947_ (.A(\control0.state[2] ),
    .B(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__nor2_1 _0948_ (.A(net34),
    .B(\control0.state[2] ),
    .Y(_0468_));
 sky130_fd_sc_hd__and2_1 _0949_ (.A(\control0.state[0] ),
    .B(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_1 _0950_ (.A(_0469_),
    .X(_0161_));
 sky130_fd_sc_hd__and3b_1 _0951_ (.A_N(\control0.state[1] ),
    .B(_0161_),
    .C(\comp0.B[0] ),
    .X(_0470_));
 sky130_fd_sc_hd__inv_2 _0952_ (.A(\control0.state[0] ),
    .Y(_0471_));
 sky130_fd_sc_hd__or4_4 _0953_ (.A(\comp0.B[10] ),
    .B(\comp0.B[9] ),
    .C(\comp0.B[8] ),
    .D(\comp0.B[7] ),
    .X(_0472_));
 sky130_fd_sc_hd__or4_4 _0954_ (.A(\comp0.B[14] ),
    .B(\comp0.B[13] ),
    .C(\comp0.B[12] ),
    .D(\comp0.B[11] ),
    .X(_0473_));
 sky130_fd_sc_hd__or4_4 _0955_ (.A(\comp0.B[6] ),
    .B(\comp0.B[5] ),
    .C(\comp0.B[4] ),
    .D(\comp0.B[3] ),
    .X(_0474_));
 sky130_fd_sc_hd__or4_4 _0956_ (.A(\comp0.B[2] ),
    .B(\comp0.B[1] ),
    .C(\comp0.B[0] ),
    .D(\comp0.B[15] ),
    .X(_0475_));
 sky130_fd_sc_hd__or4_4 _0957_ (.A(_0475_),
    .B(_0472_),
    .C(_0474_),
    .D(_0473_),
    .X(_0476_));
 sky130_fd_sc_hd__and4_1 _0958_ (.A(\control0.state[1] ),
    .B(_0471_),
    .C(_0476_),
    .D(_0468_),
    .X(_0477_));
 sky130_fd_sc_hd__a211o_1 _0959_ (.A1(net33),
    .A2(_0467_),
    .B1(_0470_),
    .C1(_0477_),
    .X(_0160_));
 sky130_fd_sc_hd__and3_1 _0960_ (.A(\control0.count[1] ),
    .B(\control0.count[0] ),
    .C(\control0.count[2] ),
    .X(_0478_));
 sky130_fd_sc_hd__a21oi_1 _0961_ (.A1(\control0.count[1] ),
    .A2(\control0.count[0] ),
    .B1(\control0.count[2] ),
    .Y(_0479_));
 sky130_fd_sc_hd__nor2_1 _0962_ (.A(_0478_),
    .B(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__xor2_1 _0963_ (.A(\control0.count[1] ),
    .B(\control0.count[0] ),
    .X(_0481_));
 sky130_fd_sc_hd__nor2_1 _0964_ (.A(_0480_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__xnor2_1 _0965_ (.A(\control0.count[3] ),
    .B(_0478_),
    .Y(_0483_));
 sky130_fd_sc_hd__o21ai_1 _0966_ (.A1(_0482_),
    .A2(_0483_),
    .B1(net236),
    .Y(_0484_));
 sky130_fd_sc_hd__or4b_4 _0967_ (.A(\control0.state[0] ),
    .B(\control0.state[2] ),
    .C(_0476_),
    .D_N(\control0.state[1] ),
    .X(_0485_));
 sky130_fd_sc_hd__nor3_1 _0968_ (.A(net34),
    .B(\control0.state[1] ),
    .C(\control0.state[0] ),
    .Y(_0486_));
 sky130_fd_sc_hd__nor2_1 _0969_ (.A(_0468_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__a21oi_2 _0970_ (.A1(_0485_),
    .A2(_0484_),
    .B1(_0487_),
    .Y(_0162_));
 sky130_fd_sc_hd__a21o_1 _0971_ (.A1(_0181_),
    .A2(_0487_),
    .B1(_0467_),
    .X(_0163_));
 sky130_fd_sc_hd__a32o_1 _0972_ (.A1(\control0.state[1] ),
    .A2(_0471_),
    .A3(_0468_),
    .B1(_0487_),
    .B2(net231),
    .X(_0164_));
 sky130_fd_sc_hd__a22o_1 _0973_ (.A1(net240),
    .A2(_0161_),
    .B1(_0487_),
    .B2(_0369_),
    .X(_0165_));
 sky130_fd_sc_hd__o21ba_1 _0974_ (.A1(net159),
    .A2(_0486_),
    .B1_N(_0468_),
    .X(_0166_));
 sky130_fd_sc_hd__and2_1 _0975_ (.A(\control0.state[2] ),
    .B(_0486_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _0976_ (.A0(_0488_),
    .A1(_0466_),
    .S(\control0.count[0] ),
    .X(_0489_));
 sky130_fd_sc_hd__clkbuf_1 _0977_ (.A(_0489_),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_1 _0978_ (.A1(net226),
    .A2(_0466_),
    .B1(_0481_),
    .B2(_0488_),
    .X(_0168_));
 sky130_fd_sc_hd__a22o_1 _0979_ (.A1(net164),
    .A2(_0466_),
    .B1(_0480_),
    .B2(_0488_),
    .X(_0169_));
 sky130_fd_sc_hd__inv_2 _0980_ (.A(_0483_),
    .Y(_0490_));
 sky130_fd_sc_hd__a22o_1 _0981_ (.A1(net167),
    .A2(_0466_),
    .B1(_0490_),
    .B2(_0488_),
    .X(_0170_));
 sky130_fd_sc_hd__dfxtp_1 _0982_ (.CLK(net68),
    .D(_0080_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _0983_ (.CLK(net69),
    .D(_0081_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _0984_ (.CLK(net70),
    .D(_0082_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _0985_ (.CLK(net71),
    .D(_0083_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _0986_ (.CLK(net72),
    .D(_0084_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 _0987_ (.CLK(net73),
    .D(_0085_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_1 _0988_ (.CLK(net74),
    .D(_0086_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _0989_ (.CLK(net75),
    .D(_0087_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_1 _0990_ (.CLK(net76),
    .D(_0088_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _0991_ (.CLK(net77),
    .D(_0089_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _0992_ (.CLK(net78),
    .D(_0090_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _0993_ (.CLK(net79),
    .D(_0091_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _0994_ (.CLK(net80),
    .D(_0092_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(net81),
    .D(_0093_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _0996_ (.CLK(net82),
    .D(_0094_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _0997_ (.CLK(net83),
    .D(_0095_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _0998_ (.CLK(net84),
    .D(_0096_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _0999_ (.CLK(net85),
    .D(_0097_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _1000_ (.CLK(net86),
    .D(_0098_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(net87),
    .D(_0099_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _1002_ (.CLK(net88),
    .D(_0100_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(net89),
    .D(_0101_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(net90),
    .D(_0102_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(net91),
    .D(_0103_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(net92),
    .D(_0104_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _1007_ (.CLK(net93),
    .D(_0105_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _1008_ (.CLK(net94),
    .D(_0106_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _1009_ (.CLK(net95),
    .D(_0107_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _1010_ (.CLK(net96),
    .D(_0108_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _1011_ (.CLK(net97),
    .D(_0109_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _1012_ (.CLK(net98),
    .D(_0110_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _1013_ (.CLK(net99),
    .D(_0111_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _1014_ (.CLK(net100),
    .D(_0112_),
    .Q(\acc0.A[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1015_ (.CLK(net101),
    .D(_0113_),
    .Q(\comp0.B[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(net102),
    .D(net166),
    .Q(\acc0.A[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1017_ (.CLK(net103),
    .D(_0115_),
    .Q(\acc0.A[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1018_ (.CLK(net104),
    .D(_0116_),
    .Q(\acc0.A[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1019_ (.CLK(net105),
    .D(net207),
    .Q(\acc0.A[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1020_ (.CLK(net106),
    .D(_0118_),
    .Q(\acc0.A[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1021_ (.CLK(net107),
    .D(_0119_),
    .Q(\acc0.A[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1022_ (.CLK(net108),
    .D(net151),
    .Q(\acc0.A[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1023_ (.CLK(net109),
    .D(net177),
    .Q(\acc0.A[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1024_ (.CLK(net110),
    .D(_0122_),
    .Q(\acc0.A[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1025_ (.CLK(net111),
    .D(net200),
    .Q(\acc0.A[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1026_ (.CLK(net112),
    .D(_0124_),
    .Q(\acc0.A[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1027_ (.CLK(net113),
    .D(net156),
    .Q(\acc0.A[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1028_ (.CLK(net114),
    .D(_0126_),
    .Q(\acc0.A[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1029_ (.CLK(net115),
    .D(net191),
    .Q(\acc0.A[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1030_ (.CLK(net116),
    .D(net209),
    .Q(\acc0.A[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1031_ (.CLK(net117),
    .D(net163),
    .Q(\acc0.A[31] ));
 sky130_fd_sc_hd__dfxtp_1 _1032_ (.CLK(net118),
    .D(net202),
    .Q(\comp0.B[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1033_ (.CLK(net119),
    .D(_0131_),
    .Q(\comp0.B[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1034_ (.CLK(net120),
    .D(net186),
    .Q(\comp0.B[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1035_ (.CLK(net121),
    .D(_0133_),
    .Q(\comp0.B[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1036_ (.CLK(net122),
    .D(net161),
    .Q(\comp0.B[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1037_ (.CLK(net123),
    .D(_0135_),
    .Q(\comp0.B[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1038_ (.CLK(net124),
    .D(net172),
    .Q(\comp0.B[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1039_ (.CLK(net125),
    .D(_0137_),
    .Q(\comp0.B[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1040_ (.CLK(net126),
    .D(net174),
    .Q(\comp0.B[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1041_ (.CLK(net127),
    .D(net153),
    .Q(\comp0.B[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1042_ (.CLK(net128),
    .D(_0140_),
    .Q(\comp0.B[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1043_ (.CLK(net129),
    .D(net196),
    .Q(\comp0.B[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1044_ (.CLK(net130),
    .D(net194),
    .Q(\comp0.B[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1045_ (.CLK(net131),
    .D(net184),
    .Q(\comp0.B[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1046_ (.CLK(net132),
    .D(net158),
    .Q(\comp0.B[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1047_ (.CLK(net133),
    .D(_0145_),
    .Q(\acc0.A[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.CLK(net134),
    .D(_0146_),
    .Q(\acc0.A[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1049_ (.CLK(net135),
    .D(_0147_),
    .Q(\acc0.A[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1050_ (.CLK(net136),
    .D(_0148_),
    .Q(\acc0.A[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1051_ (.CLK(net137),
    .D(_0149_),
    .Q(\acc0.A[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1052_ (.CLK(net138),
    .D(_0150_),
    .Q(\acc0.A[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1053_ (.CLK(net139),
    .D(_0151_),
    .Q(\acc0.A[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1054_ (.CLK(net140),
    .D(net169),
    .Q(\acc0.A[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1055_ (.CLK(net141),
    .D(net179),
    .Q(\acc0.A[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1056_ (.CLK(net142),
    .D(net182),
    .Q(\acc0.A[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1057_ (.CLK(net143),
    .D(net189),
    .Q(\acc0.A[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1058_ (.CLK(net144),
    .D(_0156_),
    .Q(\acc0.A[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1059_ (.CLK(net145),
    .D(_0157_),
    .Q(\acc0.A[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1060_ (.CLK(net146),
    .D(_0158_),
    .Q(\acc0.A[14] ));
 sky130_fd_sc_hd__dfxtp_2 _1061_ (.CLK(net147),
    .D(_0159_),
    .Q(\acc0.A[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1062_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0160_),
    .Q(\control0.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1063_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0161_),
    .Q(\control0.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1064_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0162_),
    .Q(\control0.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1065_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0163_),
    .Q(\control0.reset ));
 sky130_fd_sc_hd__dfxtp_1 _1066_ (.CLK(clknet_1_1__leaf_clk),
    .D(net232),
    .Q(\control0.sh ));
 sky130_fd_sc_hd__dfxtp_1 _1067_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0165_),
    .Q(\control0.add ));
 sky130_fd_sc_hd__dfxtp_1 _1068_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0166_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _1069_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0167_),
    .Q(\control0.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1070_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0168_),
    .Q(\control0.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1071_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0169_),
    .Q(\control0.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1072_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0170_),
    .Q(\control0.count[3] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0457_ (.A(_0457_),
    .X(clknet_0__0457_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0458_ (.A(_0458_),
    .X(clknet_0__0458_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0459_ (.A(_0459_),
    .X(clknet_0__0459_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0460_ (.A(_0460_),
    .X(clknet_0__0460_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0461_ (.A(_0461_),
    .X(clknet_0__0461_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0462_ (.A(_0462_),
    .X(clknet_0__0462_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0463_ (.A(_0463_),
    .X(clknet_0__0463_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0464_ (.A(_0464_),
    .X(clknet_0__0464_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0465_ (.A(_0465_),
    .X(clknet_0__0465_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0457_ (.A(clknet_0__0457_),
    .X(clknet_1_0__leaf__0457_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0458_ (.A(clknet_0__0458_),
    .X(clknet_1_0__leaf__0458_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0459_ (.A(clknet_0__0459_),
    .X(clknet_1_0__leaf__0459_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0460_ (.A(clknet_0__0460_),
    .X(clknet_1_0__leaf__0460_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0461_ (.A(clknet_0__0461_),
    .X(clknet_1_0__leaf__0461_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0462_ (.A(clknet_0__0462_),
    .X(clknet_1_0__leaf__0462_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0463_ (.A(clknet_0__0463_),
    .X(clknet_1_0__leaf__0463_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0464_ (.A(clknet_0__0464_),
    .X(clknet_1_0__leaf__0464_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0465_ (.A(clknet_0__0465_),
    .X(clknet_1_0__leaf__0465_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0457_ (.A(clknet_0__0457_),
    .X(clknet_1_1__leaf__0457_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0458_ (.A(clknet_0__0458_),
    .X(clknet_1_1__leaf__0458_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0459_ (.A(clknet_0__0459_),
    .X(clknet_1_1__leaf__0459_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0460_ (.A(clknet_0__0460_),
    .X(clknet_1_1__leaf__0460_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0461_ (.A(clknet_0__0461_),
    .X(clknet_1_1__leaf__0461_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0462_ (.A(clknet_0__0462_),
    .X(clknet_1_1__leaf__0462_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0463_ (.A(clknet_0__0463_),
    .X(clknet_1_1__leaf__0463_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0464_ (.A(clknet_0__0464_),
    .X(clknet_1_1__leaf__0464_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0465_ (.A(clknet_0__0465_),
    .X(clknet_1_1__leaf__0465_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload0 (.A(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_1_0__leaf__0465_));
 sky130_fd_sc_hd__clkinvlp_4 clkload2 (.A(clknet_1_0__leaf__0464_));
 sky130_fd_sc_hd__clkinvlp_4 clkload3 (.A(clknet_1_1__leaf__0461_));
 sky130_fd_sc_hd__clkinvlp_4 clkload4 (.A(clknet_1_0__leaf__0459_));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\acc0.A[5] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\comp0.B[15] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\acc0.A[14] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net63),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0144_),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net35),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\comp0.B[5] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0134_),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\acc0.A[31] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0129_),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\control0.count[2] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\acc0.A[15] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0114_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\acc0.A[0] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\control0.count[3] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\acc0.A[7] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0152_),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\acc0.A[3] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\comp0.B[7] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0136_),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\comp0.B[9] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0138_),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\acc0.A[2] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\acc0.A[22] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\acc0.A[21] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0121_),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\acc0.A[8] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0153_),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\comp0.B[8] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\acc0.A[9] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_0154_),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\comp0.B[14] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0143_),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\comp0.B[3] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0132_),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0120_),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\acc0.A[20] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\acc0.A[10] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0155_),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\acc0.A[28] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0127_),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\acc0.A[11] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\comp0.B[13] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0142_),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\comp0.B[12] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0141_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\comp0.B[10] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\acc0.A[27] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\comp0.B[11] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\acc0.A[24] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0123_),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\comp0.B[1] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0130_),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\comp0.B[2] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\comp0.B[6] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\comp0.B[4] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\acc0.A[18] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0139_),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0117_),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\acc0.A[30] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0128_),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\acc0.A[25] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\acc0.A[19] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net65),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net49),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net66),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\acc0.A[23] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net52),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\acc0.A[4] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net37),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\acc0.A[1] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\acc0.A[17] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net48),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\acc0.A[16] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net58),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net46),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net55),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net60),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\control0.count[1] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\acc0.A[26] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net57),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\acc0.A[12] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\acc0.A[13] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\acc0.A[6] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\control0.sh ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_0164_),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net61),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net36),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net64),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\control0.state[2] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0125_),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net53),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net41),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net59),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\control0.state[1] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net51),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net56),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net50),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net54),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net40),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net38),
    .X(net246));
 sky130_fd_sc_hd__buf_1 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(A[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(A[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(A[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(A[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(A[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(A[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(A[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(B[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(B[10]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(B[11]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(B[12]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(B[13]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(B[14]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(B[15]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(B[1]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(B[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(B[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(B[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(B[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(B[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(B[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(B[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(B[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(init),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(rst),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(A[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(A[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(done));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(pp[0]));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net37),
    .X(pp[10]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(pp[11]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(pp[12]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(pp[13]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(pp[14]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(pp[15]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(pp[16]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(pp[17]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(pp[18]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(pp[19]));
 sky130_fd_sc_hd__clkbuf_4 output47 (.A(net47),
    .X(pp[1]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(pp[20]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(pp[21]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(pp[22]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(pp[23]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(pp[24]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(pp[25]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(pp[26]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(pp[27]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(pp[28]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(pp[29]));
 sky130_fd_sc_hd__clkbuf_4 output58 (.A(net58),
    .X(pp[2]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(pp[30]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(pp[31]));
 sky130_fd_sc_hd__clkbuf_4 output61 (.A(net61),
    .X(pp[3]));
 sky130_fd_sc_hd__clkbuf_4 output62 (.A(net62),
    .X(pp[4]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .X(pp[5]));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net64),
    .X(pp[6]));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(pp[7]));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(pp[8]));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(pp[9]));
endmodule

