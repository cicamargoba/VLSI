* SPICE3 file created from mult_32.ext - technology: sky130A

X0 net101 clknet_1_0__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND clknet_1_0__leaf__0461_ net101 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 net101 clknet_1_0__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR clknet_1_0__leaf__0461_ net101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 net61 _0985_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 _0985_/a_891_413# _0985_/a_193_47# _0985_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6 _0985_/a_561_413# _0985_/a_27_47# _0985_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7 VPWR net71 _0985_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 net61 _0985_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 _0985_/a_381_47# _0083_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND _0985_/a_634_159# _0985_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11 VPWR _0985_/a_891_413# _0985_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12 _0985_/a_466_413# _0985_/a_193_47# _0985_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13 VPWR _0985_/a_634_159# _0985_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14 _0985_/a_634_159# _0985_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15 _0985_/a_634_159# _0985_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X16 _0985_/a_975_413# _0985_/a_193_47# _0985_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VGND _0985_/a_1059_315# _0985_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X18 _0985_/a_193_47# _0985_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 _0985_/a_891_413# _0985_/a_27_47# _0985_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X20 _0985_/a_592_47# _0985_/a_193_47# _0985_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X21 VPWR _0985_/a_1059_315# _0985_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X22 _0985_/a_1017_47# _0985_/a_27_47# _0985_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X23 _0985_/a_193_47# _0985_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 _0985_/a_466_413# _0985_/a_27_47# _0985_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X25 VGND _0985_/a_891_413# _0985_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X26 _0985_/a_381_47# _0083_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 VGND net71 _0985_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X28 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=707.2962 ps=6.62772k w=0.87 l=1.05
X29 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=450.85931 ps=4.80461k w=0.55 l=1.05
X30 VPWR _0243_ _0770_/a_382_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X31 _0770_/a_297_47# control0.add _0770_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X32 _0770_/a_297_47# _0243_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VGND _0389_ _0770_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X34 VPWR _0770_/a_79_21# _0390_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X35 _0770_/a_79_21# control0.add VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X36 _0770_/a_382_297# _0389_ _0770_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X37 VGND _0770_/a_79_21# _0390_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X38 net82 clknet_1_0__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X39 VGND clknet_1_0__leaf__0459_ net82 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X40 net82 clknet_1_0__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X41 VPWR clknet_1_0__leaf__0459_ net82 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X42 VPWR net34 _0968_/a_193_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X43 _0968_/a_193_297# control0.state\[1\] _0968_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X44 _0486_ control0.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X45 VGND net34 _0486_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X46 _0968_/a_109_297# control0.state\[0\] _0486_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X47 VGND control0.state\[0\] _0486_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X48 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X49 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X50 VPWR acc0.A\[6\] _0822_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X51 VGND acc0.A\[6\] _0430_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 _0822_/a_109_297# net64 _0430_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X53 _0430_ net64 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X54 _0753_/a_465_47# _0233_ _0753_/a_381_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 VGND _0375_ _0753_/a_561_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X56 VPWR _0231_ _0753_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X57 _0753_/a_297_297# _0233_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X58 _0753_/a_297_297# _0375_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X59 VPWR _0222_ _0753_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X60 _0753_/a_381_47# _0222_ _0753_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18362 ps=1.215 w=0.65 l=0.15
X61 _0753_/a_297_297# _0343_ _0753_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X62 VPWR _0753_/a_79_21# _0377_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X63 _0753_/a_79_21# _0343_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.18362 pd=1.215 as=0.16087 ps=1.145 w=0.65 l=0.15
X64 VGND _0753_/a_79_21# _0377_ VGND sky130_fd_pr__nfet_01v8 ad=0.16087 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X65 _0753_/a_561_47# _0231_ _0753_/a_465_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X66 VPWR net55 _0684_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X67 _0316_ _0684_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X68 VGND net55 _0684_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X69 _0684_/a_59_75# acc0.A\[27\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X70 _0316_ _0684_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X71 _0684_/a_145_75# acc0.A\[27\] _0684_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X72 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X73 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X74 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X75 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X76 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X77 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X78 acc0.A\[21\] _1021_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X79 _1021_/a_891_413# _1021_/a_193_47# _1021_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X80 _1021_/a_561_413# _1021_/a_27_47# _1021_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X81 VPWR net107 _1021_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X82 acc0.A\[21\] _1021_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X83 _1021_/a_381_47# _0119_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X84 VGND _1021_/a_634_159# _1021_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X85 VPWR _1021_/a_891_413# _1021_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X86 _1021_/a_466_413# _1021_/a_193_47# _1021_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X87 VPWR _1021_/a_634_159# _1021_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X88 _1021_/a_634_159# _1021_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X89 _1021_/a_634_159# _1021_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X90 _1021_/a_975_413# _1021_/a_193_47# _1021_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X91 VGND _1021_/a_1059_315# _1021_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X92 _1021_/a_193_47# _1021_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X93 _1021_/a_891_413# _1021_/a_27_47# _1021_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X94 _1021_/a_592_47# _1021_/a_193_47# _1021_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X95 VPWR _1021_/a_1059_315# _1021_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X96 _1021_/a_1017_47# _1021_/a_27_47# _1021_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X97 _1021_/a_193_47# _1021_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X98 _1021_/a_466_413# _1021_/a_27_47# _1021_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X99 VGND _1021_/a_891_413# _1021_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X100 _1021_/a_381_47# _0119_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X101 VGND net107 _1021_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X102 VPWR _0281_ _0805_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X103 VPWR _0402_ _0805_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X104 _0805_/a_181_47# _0286_ _0805_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X105 VGND _0402_ _0805_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X106 _0805_/a_27_47# _0286_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X107 _0417_ _0805_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X108 _0417_ _0805_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X109 _0805_/a_109_47# _0281_ _0805_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X110 _0736_/a_56_297# _0219_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X111 VPWR _0362_ _0736_/a_56_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X112 _0107_ _0181_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X113 _0736_/a_139_47# _0362_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2665 ps=2.12 w=0.65 l=0.15
X114 _0736_/a_311_297# _0363_ _0736_/a_56_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X115 _0107_ _0181_ _0736_/a_311_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X116 VGND _0363_ _0107_ VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X117 _0107_ _0219_ _0736_/a_139_47# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X118 VPWR _0226_ _0598_/a_382_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.305 ps=2.61 w=1 l=0.15
X119 _0598_/a_297_47# _0229_ _0598_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.3705 pd=3.74 as=0.169 ps=1.82 w=0.65 l=0.15
X120 _0598_/a_297_47# _0226_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X121 VGND _0227_ _0598_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X122 VPWR _0598_/a_79_21# _0230_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X123 _0598_/a_79_21# _0229_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.15
X124 _0598_/a_382_297# _0227_ _0598_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X125 VGND _0598_/a_79_21# _0230_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X126 VPWR acc0.A\[13\] _0299_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X127 _0299_ acc0.A\[13\] _0667_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X128 _0667_/a_113_47# net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X129 _0299_ net40 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X130 VPWR clknet_0__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X131 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X132 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X133 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X134 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X135 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X136 clkbuf_1_0__f__0459_/a_110_47# clknet_0__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X137 clkbuf_1_0__f__0459_/a_110_47# clknet_0__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X138 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X139 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X140 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X141 clkbuf_1_0__f__0459_/a_110_47# clknet_0__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X142 VGND clknet_0__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X143 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X144 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X145 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X146 VGND clknet_0__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X147 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X148 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X149 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X150 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X151 clkbuf_1_0__f__0459_/a_110_47# clknet_0__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X152 VPWR clknet_0__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X153 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X154 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X155 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X156 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X157 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X158 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X159 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X160 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X161 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X162 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X163 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X164 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X165 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X166 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X167 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X168 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X169 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X170 VPWR _0121_ hold30/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X171 VGND hold30/a_285_47# hold30/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X172 net177 hold30/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X173 VGND _0121_ hold30/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X174 VPWR hold30/a_285_47# hold30/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X175 hold30/a_285_47# hold30/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X176 hold30/a_285_47# hold30/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X177 net177 hold30/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X178 VPWR acc0.A\[10\] hold41/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X179 VGND hold41/a_285_47# hold41/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X180 net188 hold41/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X181 VGND acc0.A\[10\] hold41/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X182 VPWR hold41/a_285_47# hold41/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X183 hold41/a_285_47# hold41/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X184 hold41/a_285_47# hold41/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X185 net188 hold41/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X186 VPWR acc0.A\[24\] hold52/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X187 VGND hold52/a_285_47# hold52/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X188 net199 hold52/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X189 VGND acc0.A\[24\] hold52/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X190 VPWR hold52/a_285_47# hold52/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X191 hold52/a_285_47# hold52/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X192 hold52/a_285_47# hold52/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X193 net199 hold52/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X194 VPWR acc0.A\[25\] hold63/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X195 VGND hold63/a_285_47# hold63/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X196 net210 hold63/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X197 VGND acc0.A\[25\] hold63/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X198 VPWR hold63/a_285_47# hold63/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X199 hold63/a_285_47# hold63/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X200 hold63/a_285_47# hold63/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X201 net210 hold63/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X202 VPWR acc0.A\[16\] hold74/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X203 VGND hold74/a_285_47# hold74/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X204 net221 hold74/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X205 VGND acc0.A\[16\] hold74/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X206 VPWR hold74/a_285_47# hold74/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X207 hold74/a_285_47# hold74/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X208 hold74/a_285_47# hold74/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X209 net221 hold74/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X212 VPWR _0164_ hold85/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X213 VGND hold85/a_285_47# hold85/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X214 net232 hold85/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X215 VGND _0164_ hold85/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X216 VPWR hold85/a_285_47# hold85/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X217 hold85/a_285_47# hold85/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X218 hold85/a_285_47# hold85/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X219 net232 hold85/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X220 VPWR net50 hold96/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X221 VGND hold96/a_285_47# hold96/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X222 net243 hold96/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X223 VGND net50 hold96/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X224 VPWR hold96/a_285_47# hold96/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X225 hold96/a_285_47# hold96/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X226 hold96/a_285_47# hold96/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X227 net243 hold96/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X232 _0521_/a_81_21# _0192_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08937 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X233 _0521_/a_299_297# _0192_ _0521_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X234 VPWR _0521_/a_81_21# _0151_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X235 VPWR net230 _0521_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X236 VGND _0521_/a_81_21# _0151_ VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X237 VGND _0179_ _0521_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X238 _0521_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X239 _0521_/a_384_47# net230 _0521_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08937 ps=0.925 w=0.65 l=0.15
X240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X242 net50 _1004_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X243 _1004_/a_891_413# _1004_/a_193_47# _1004_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X244 _1004_/a_561_413# _1004_/a_27_47# _1004_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X245 VPWR net90 _1004_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X246 net50 _1004_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X247 _1004_/a_381_47# _0102_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X248 VGND _1004_/a_634_159# _1004_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X249 VPWR _1004_/a_891_413# _1004_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X250 _1004_/a_466_413# _1004_/a_193_47# _1004_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X251 VPWR _1004_/a_634_159# _1004_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X252 _1004_/a_634_159# _1004_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X253 _1004_/a_634_159# _1004_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X254 _1004_/a_975_413# _1004_/a_193_47# _1004_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X255 VGND _1004_/a_1059_315# _1004_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X256 _1004_/a_193_47# _1004_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X257 _1004_/a_891_413# _1004_/a_27_47# _1004_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X258 _1004_/a_592_47# _1004_/a_193_47# _1004_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X259 VPWR _1004_/a_1059_315# _1004_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X260 _1004_/a_1017_47# _1004_/a_27_47# _1004_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X261 _1004_/a_193_47# _1004_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X262 _1004_/a_466_413# _1004_/a_27_47# _1004_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X263 VGND _1004_/a_891_413# _1004_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X264 _1004_/a_381_47# _0102_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X265 VGND net90 _1004_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X266 VPWR _0719_/a_27_47# _0350_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X267 _0350_ _0719_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X268 VPWR control0.add _0719_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X269 _0350_ _0719_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X270 VGND _0719_/a_27_47# _0350_ VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X271 VGND control0.add _0719_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X274 VPWR output53/a_27_47# pp[25] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X275 pp[25] output53/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X276 VPWR net53 output53/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X277 pp[25] output53/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X278 VGND output53/a_27_47# pp[25] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X279 VGND net53 output53/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X280 VPWR output42/a_27_47# pp[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X281 pp[15] output42/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X282 VPWR net42 output42/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X283 pp[15] output42/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X284 VGND output42/a_27_47# pp[15] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X285 VGND net42 output42/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X286 VPWR net64 output64/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X287 VGND output64/a_27_47# pp[6] VGND sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X288 VGND output64/a_27_47# pp[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X289 pp[6] output64/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X290 pp[6] output64/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X291 VGND net64 output64/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X292 VPWR output64/a_27_47# pp[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X293 pp[6] output64/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X294 pp[6] output64/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X295 VPWR output64/a_27_47# pp[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X298 VPWR _0182_ _0504_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X299 VGND _0504_/a_27_47# _0183_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X300 VGND _0504_/a_27_47# _0183_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X301 _0183_ _0504_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X302 _0183_ _0504_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X303 VGND _0182_ _0504_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X304 VPWR _0504_/a_27_47# _0183_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X305 _0183_ _0504_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X306 _0183_ _0504_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X307 VPWR _0504_/a_27_47# _0183_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X316 net58 _0984_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X317 _0984_/a_891_413# _0984_/a_193_47# _0984_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X318 _0984_/a_561_413# _0984_/a_27_47# _0984_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X319 VPWR net70 _0984_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X320 net58 _0984_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X321 _0984_/a_381_47# _0082_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X322 VGND _0984_/a_634_159# _0984_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X323 VPWR _0984_/a_891_413# _0984_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X324 _0984_/a_466_413# _0984_/a_193_47# _0984_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X325 VPWR _0984_/a_634_159# _0984_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X326 _0984_/a_634_159# _0984_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X327 _0984_/a_634_159# _0984_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X328 _0984_/a_975_413# _0984_/a_193_47# _0984_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X329 VGND _0984_/a_1059_315# _0984_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X330 _0984_/a_193_47# _0984_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X331 _0984_/a_891_413# _0984_/a_27_47# _0984_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X332 _0984_/a_592_47# _0984_/a_193_47# _0984_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X333 VPWR _0984_/a_1059_315# _0984_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X334 _0984_/a_1017_47# _0984_/a_27_47# _0984_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X335 _0984_/a_193_47# _0984_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X336 _0984_/a_466_413# _0984_/a_27_47# _0984_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X337 VGND _0984_/a_891_413# _0984_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X338 _0984_/a_381_47# _0082_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X339 VGND net70 _0984_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X344 _0485_ _0967_/a_215_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X345 VGND _0967_/a_215_297# _0485_ VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X346 VPWR _0967_/a_215_297# _0485_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X347 _0967_/a_109_93# control0.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X348 _0967_/a_215_297# _0967_/a_109_93# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X349 VGND _0476_ _0967_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X350 VGND control0.state\[0\] _0967_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X351 _0485_ _0967_/a_215_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X352 _0967_/a_215_297# control0.state\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X353 _0967_/a_109_93# control0.state\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X354 VPWR control0.state\[0\] _0967_/a_487_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X355 VGND _0967_/a_215_297# _0485_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X356 _0967_/a_487_297# control0.state\[2\] _0967_/a_403_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X357 _0967_/a_403_297# _0476_ _0967_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X358 VPWR _0967_/a_215_297# _0485_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X359 _0485_ _0967_/a_215_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X360 _0485_ _0967_/a_215_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X361 _0967_/a_297_297# _0967_/a_109_93# _0967_/a_215_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X362 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X363 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X364 net139 clknet_1_0__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X365 VGND clknet_1_0__leaf__0465_ net139 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X366 net139 clknet_1_0__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X367 VPWR clknet_1_0__leaf__0465_ net139 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X372 _0752_/a_300_297# _0752_/a_27_413# _0376_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X373 VGND _0375_ _0752_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X374 VPWR _0234_ _0752_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X375 _0376_ _0752_/a_27_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.10187 ps=0.99 w=0.65 l=0.15
X376 VPWR _0222_ _0752_/a_300_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X377 _0752_/a_384_47# _0222_ _0376_ VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X378 VGND _0234_ _0752_/a_27_413# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.1113 ps=1.37 w=0.42 l=0.15
X379 _0752_/a_300_297# _0375_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X380 VPWR _0251_ _0429_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X381 _0429_ _0251_ _0821_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X382 _0821_/a_113_47# _0252_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X383 _0429_ _0252_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X384 VPWR _0313_ _0315_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X385 _0315_ _0313_ _0683_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X386 _0683_/a_113_47# _0314_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X387 _0315_ _0314_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X392 net120 clknet_1_1__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X393 VGND clknet_1_1__leaf__0463_ net120 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X394 net120 clknet_1_1__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X395 VPWR clknet_1_1__leaf__0463_ net120 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X396 acc0.A\[20\] _1020_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X397 _1020_/a_891_413# _1020_/a_193_47# _1020_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X398 _1020_/a_561_413# _1020_/a_27_47# _1020_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X399 VPWR net106 _1020_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X400 acc0.A\[20\] _1020_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X401 _1020_/a_381_47# _0118_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X402 VGND _1020_/a_634_159# _1020_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X403 VPWR _1020_/a_891_413# _1020_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X404 _1020_/a_466_413# _1020_/a_193_47# _1020_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X405 VPWR _1020_/a_634_159# _1020_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X406 _1020_/a_634_159# _1020_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X407 _1020_/a_634_159# _1020_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X408 _1020_/a_975_413# _1020_/a_193_47# _1020_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X409 VGND _1020_/a_1059_315# _1020_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X410 _1020_/a_193_47# _1020_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X411 _1020_/a_891_413# _1020_/a_27_47# _1020_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X412 _1020_/a_592_47# _1020_/a_193_47# _1020_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X413 VPWR _1020_/a_1059_315# _1020_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X414 _1020_/a_1017_47# _1020_/a_27_47# _1020_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X415 _1020_/a_193_47# _1020_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X416 _1020_/a_466_413# _1020_/a_27_47# _1020_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X417 VGND _1020_/a_891_413# _1020_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X418 _1020_/a_381_47# _0118_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X419 VGND net106 _1020_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X420 net134 clknet_1_0__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X421 VGND clknet_1_0__leaf__0464_ net134 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X422 net134 clknet_1_0__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X423 VPWR clknet_1_0__leaf__0464_ net134 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X424 VPWR clknet_0__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X425 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X426 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X427 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X428 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X429 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X430 clkbuf_1_0__f__0458_/a_110_47# clknet_0__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X431 clkbuf_1_0__f__0458_/a_110_47# clknet_0__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X432 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X433 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X434 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X435 clkbuf_1_0__f__0458_/a_110_47# clknet_0__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X436 VGND clknet_0__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X437 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X438 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X439 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X440 VGND clknet_0__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X441 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X442 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X443 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X444 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X445 clkbuf_1_0__f__0458_/a_110_47# clknet_0__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X446 VPWR clknet_0__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X447 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X448 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X449 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X450 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X451 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X452 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X453 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X454 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X455 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X456 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X457 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X458 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X459 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X460 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X461 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X462 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X463 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X464 VPWR _0350_ _0735_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X465 VGND _0350_ _0363_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X466 _0735_/a_109_297# net224 _0363_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X467 _0363_ net224 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X468 VGND _0347_ _0804_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X469 _0804_/a_510_47# _0416_ _0804_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X470 _0804_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X471 VPWR _0416_ _0804_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X472 _0804_/a_79_21# _0415_ _0804_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X473 _0804_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X474 _0804_/a_79_21# _0399_ _0804_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X475 VPWR _0804_/a_79_21# _0092_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X476 VGND _0804_/a_79_21# _0092_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X477 _0804_/a_215_47# _0415_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.10563 ps=0.975 w=0.65 l=0.15
X478 VPWR acc0.A\[12\] _0298_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X479 _0298_ acc0.A\[12\] _0666_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X480 _0666_/a_113_47# net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X481 _0298_ net39 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X482 _0229_ _0228_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X483 VGND _0228_ _0229_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X484 _0229_ _0228_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X485 VPWR _0228_ _0229_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X486 VPWR control0.count\[3\] hold20/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X487 VGND hold20/a_285_47# hold20/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X488 net167 hold20/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X489 VGND control0.count\[3\] hold20/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X490 VPWR hold20/a_285_47# hold20/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X491 hold20/a_285_47# hold20/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X492 hold20/a_285_47# hold20/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X493 net167 hold20/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X494 VPWR acc0.A\[8\] hold31/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X495 VGND hold31/a_285_47# hold31/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X496 net178 hold31/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X497 VGND acc0.A\[8\] hold31/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X498 VPWR hold31/a_285_47# hold31/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X499 hold31/a_285_47# hold31/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X500 hold31/a_285_47# hold31/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X501 net178 hold31/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X502 VPWR _0155_ hold42/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X503 VGND hold42/a_285_47# hold42/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X504 net189 hold42/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X505 VGND _0155_ hold42/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X506 VPWR hold42/a_285_47# hold42/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X507 hold42/a_285_47# hold42/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X508 hold42/a_285_47# hold42/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X509 net189 hold42/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X510 VPWR _0123_ hold53/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X511 VGND hold53/a_285_47# hold53/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X512 net200 hold53/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X513 VGND _0123_ hold53/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X514 VPWR hold53/a_285_47# hold53/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X515 hold53/a_285_47# hold53/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X516 hold53/a_285_47# hold53/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X517 net200 hold53/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X518 VPWR acc0.A\[19\] hold64/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X519 VGND hold64/a_285_47# hold64/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X520 net211 hold64/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X521 VGND acc0.A\[19\] hold64/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X522 VPWR hold64/a_285_47# hold64/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X523 hold64/a_285_47# hold64/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X524 hold64/a_285_47# hold64/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X525 net211 hold64/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X526 VPWR net58 hold75/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X527 VGND hold75/a_285_47# hold75/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X528 net222 hold75/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X529 VGND net58 hold75/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X530 VPWR hold75/a_285_47# hold75/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X531 hold75/a_285_47# hold75/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X532 hold75/a_285_47# hold75/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X533 net222 hold75/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X534 VPWR net61 hold86/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X535 VGND hold86/a_285_47# hold86/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X536 net233 hold86/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X537 VGND net61 hold86/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X538 VPWR hold86/a_285_47# hold86/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X539 hold86/a_285_47# hold86/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X540 hold86/a_285_47# hold86/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X541 net233 hold86/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X542 VPWR net54 hold97/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X543 VGND hold97/a_285_47# hold97/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X544 net244 hold97/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X545 VGND net54 hold97/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X546 VPWR hold97/a_285_47# hold97/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X547 hold97/a_285_47# hold97/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X548 hold97/a_285_47# hold97/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X549 net244 hold97/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X552 VPWR net14 _0520_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X553 _0520_/a_27_297# _0186_ _0520_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X554 VGND net14 _0520_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X555 _0192_ _0520_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X556 _0520_/a_27_297# _0186_ _0520_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X557 _0520_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X558 _0520_/a_373_47# _0180_ _0520_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X559 _0192_ _0520_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X560 _0520_/a_109_297# net168 _0520_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X561 _0520_/a_109_47# net168 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X562 net49 _1003_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X563 _1003_/a_891_413# _1003_/a_193_47# _1003_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X564 _1003_/a_561_413# _1003_/a_27_47# _1003_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X565 VPWR net89 _1003_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X566 net49 _1003_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X567 _1003_/a_381_47# _0101_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X568 VGND _1003_/a_634_159# _1003_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X569 VPWR _1003_/a_891_413# _1003_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X570 _1003_/a_466_413# _1003_/a_193_47# _1003_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X571 VPWR _1003_/a_634_159# _1003_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X572 _1003_/a_634_159# _1003_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X573 _1003_/a_634_159# _1003_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X574 _1003_/a_975_413# _1003_/a_193_47# _1003_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X575 VGND _1003_/a_1059_315# _1003_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X576 _1003_/a_193_47# _1003_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X577 _1003_/a_891_413# _1003_/a_27_47# _1003_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X578 _1003_/a_592_47# _1003_/a_193_47# _1003_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X579 VPWR _1003_/a_1059_315# _1003_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X580 _1003_/a_1017_47# _1003_/a_27_47# _1003_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X581 _1003_/a_193_47# _1003_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X582 _1003_/a_466_413# _1003_/a_27_47# _1003_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X583 VGND _1003_/a_891_413# _1003_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X584 _1003_/a_381_47# _0101_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X585 VGND net89 _1003_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X588 _0718_/a_377_297# _0337_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X589 _0718_/a_47_47# _0348_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X590 _0718_/a_129_47# _0348_ _0718_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X591 _0718_/a_285_47# _0348_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X592 _0349_ _0718_/a_47_47# _0718_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X593 VGND _0337_ _0718_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X594 VPWR _0337_ _0718_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X595 VPWR _0718_/a_47_47# _0349_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X596 _0349_ _0348_ _0718_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X597 _0718_/a_285_47# _0337_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X598 VPWR acc0.A\[10\] _0281_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X599 _0281_ acc0.A\[10\] _0649_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X600 _0649_/a_113_47# net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X601 _0281_ net37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X604 net115 clknet_1_1__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X605 VGND clknet_1_1__leaf__0462_ net115 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X606 net115 clknet_1_1__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X607 VPWR clknet_1_1__leaf__0462_ net115 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X608 VPWR output54/a_27_47# pp[26] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X609 pp[26] output54/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X610 VPWR net54 output54/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X611 pp[26] output54/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X612 VGND output54/a_27_47# pp[26] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X613 VGND net54 output54/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X614 VPWR output43/a_27_47# pp[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X615 pp[16] output43/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X616 VPWR net43 output43/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X617 pp[16] output43/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X618 VGND output43/a_27_47# pp[16] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X619 VGND net43 output43/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X620 VPWR net65 output65/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X621 VGND output65/a_27_47# pp[7] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X622 VGND output65/a_27_47# pp[7] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X623 pp[7] output65/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X624 pp[7] output65/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X625 VGND net65 output65/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X626 VPWR output65/a_27_47# pp[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X627 pp[7] output65/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X628 pp[7] output65/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X629 VPWR output65/a_27_47# pp[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X630 VPWR _0180_ _0503_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X631 VGND _0180_ _0182_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X632 _0503_/a_109_297# control0.sh _0182_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X633 _0182_ control0.sh VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X634 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X635 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X636 net47 _0983_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X637 _0983_/a_891_413# _0983_/a_193_47# _0983_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X638 _0983_/a_561_413# _0983_/a_27_47# _0983_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X639 VPWR net69 _0983_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X640 net47 _0983_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X641 _0983_/a_381_47# _0081_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X642 VGND _0983_/a_634_159# _0983_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X643 VPWR _0983_/a_891_413# _0983_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X644 _0983_/a_466_413# _0983_/a_193_47# _0983_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X645 VPWR _0983_/a_634_159# _0983_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X646 _0983_/a_634_159# _0983_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X647 _0983_/a_634_159# _0983_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X648 _0983_/a_975_413# _0983_/a_193_47# _0983_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X649 VGND _0983_/a_1059_315# _0983_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X650 _0983_/a_193_47# _0983_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X651 _0983_/a_891_413# _0983_/a_27_47# _0983_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X652 _0983_/a_592_47# _0983_/a_193_47# _0983_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X653 VPWR _0983_/a_1059_315# _0983_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X654 _0983_/a_1017_47# _0983_/a_27_47# _0983_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X655 _0983_/a_193_47# _0983_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X656 _0983_/a_466_413# _0983_/a_27_47# _0983_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X657 VGND _0983_/a_891_413# _0983_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X658 _0983_/a_381_47# _0081_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X659 VGND net69 _0983_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X660 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X662 _0484_ _0483_ _0966_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X663 VPWR net236 _0484_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X664 _0966_/a_27_47# _0483_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X665 _0484_ net236 _0966_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X666 _0966_/a_109_297# _0482_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X667 VGND _0482_ _0966_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X668 _0375_ _0751_/a_29_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X669 _0751_/a_111_297# _0374_ _0751_/a_29_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X670 _0375_ _0751_/a_29_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.10187 ps=0.99 w=0.65 l=0.15
X671 _0751_/a_183_297# _0227_ _0751_/a_111_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X672 VPWR _0225_ _0751_/a_183_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X673 _0751_/a_29_53# _0227_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X674 VGND _0374_ _0751_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X675 VGND _0225_ _0751_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X676 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X677 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X678 VGND _0369_ _0820_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X679 _0820_/a_510_47# _0428_ _0820_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X680 _0820_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X681 VPWR _0428_ _0820_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X682 _0820_/a_79_21# net214 _0820_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X683 _0820_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X684 _0820_/a_79_21# _0399_ _0820_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X685 VPWR _0820_/a_79_21# _0088_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X686 VGND _0820_/a_79_21# _0088_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X687 _0820_/a_215_47# net214 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X690 VGND acc0.A\[25\] _0682_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X691 _0682_/a_68_297# net53 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X692 _0314_ _0682_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X693 VPWR acc0.A\[25\] _0682_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X694 _0314_ _0682_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X695 _0682_/a_150_297# net53 _0682_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X698 VPWR _0468_ _0949_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X699 _0469_ _0949_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X700 VGND _0468_ _0949_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X701 _0949_/a_59_75# control0.state\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X702 _0469_ _0949_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X703 _0949_/a_145_75# control0.state\[0\] _0949_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X706 VGND _0218_ _0803_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X707 _0803_/a_68_297# net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X708 _0416_ _0803_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X709 VPWR _0218_ _0803_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X710 _0416_ _0803_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X711 _0803_/a_150_297# net39 _0803_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X714 VPWR clknet_0__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X715 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X716 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X717 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X718 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X719 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X720 clkbuf_1_0__f__0457_/a_110_47# clknet_0__0457_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X721 clkbuf_1_0__f__0457_/a_110_47# clknet_0__0457_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X722 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X723 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X724 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X725 clkbuf_1_0__f__0457_/a_110_47# clknet_0__0457_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X726 VGND clknet_0__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X727 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X728 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X729 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X730 VGND clknet_0__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X731 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X732 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X733 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X734 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X735 clkbuf_1_0__f__0457_/a_110_47# clknet_0__0457_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X736 VPWR clknet_0__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X737 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X738 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X739 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X740 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X741 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X742 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X743 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X744 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X745 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X746 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X747 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X748 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X749 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X750 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X751 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X752 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X753 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X754 VPWR acc0.A\[13\] _0665_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X755 VGND acc0.A\[13\] _0297_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X756 _0665_/a_109_297# net40 _0297_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X757 _0297_ net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X758 _0734_/a_377_297# _0318_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X759 _0734_/a_47_47# _0361_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X760 _0734_/a_129_47# _0361_ _0734_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X761 _0734_/a_285_47# _0361_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X762 _0362_ _0734_/a_47_47# _0734_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X763 VGND _0318_ _0734_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X764 VPWR _0318_ _0734_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X765 VPWR _0734_/a_47_47# _0362_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X766 _0362_ _0361_ _0734_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X767 _0734_/a_285_47# _0318_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X768 VPWR net49 _0596_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X769 _0228_ _0596_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X770 VGND net49 _0596_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X771 _0596_/a_59_75# acc0.A\[21\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X772 _0228_ _0596_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X773 _0596_/a_145_75# acc0.A\[21\] _0596_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X776 VPWR comp0.B\[15\] hold10/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X777 VGND hold10/a_285_47# hold10/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X778 net157 hold10/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X779 VGND comp0.B\[15\] hold10/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X780 VPWR hold10/a_285_47# hold10/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X781 hold10/a_285_47# hold10/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X782 hold10/a_285_47# hold10/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X783 net157 hold10/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X784 VPWR acc0.A\[7\] hold21/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X785 VGND hold21/a_285_47# hold21/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X786 net168 hold21/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X787 VGND acc0.A\[7\] hold21/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X788 VPWR hold21/a_285_47# hold21/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X789 hold21/a_285_47# hold21/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X790 hold21/a_285_47# hold21/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X791 net168 hold21/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X792 VPWR _0153_ hold32/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X793 VGND hold32/a_285_47# hold32/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X794 net179 hold32/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X795 VGND _0153_ hold32/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X796 VPWR hold32/a_285_47# hold32/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X797 hold32/a_285_47# hold32/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X798 hold32/a_285_47# hold32/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X799 net179 hold32/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X800 VPWR acc0.A\[28\] hold43/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X801 VGND hold43/a_285_47# hold43/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X802 net190 hold43/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X803 VGND acc0.A\[28\] hold43/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X804 VPWR hold43/a_285_47# hold43/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X805 hold43/a_285_47# hold43/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X806 hold43/a_285_47# hold43/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X807 net190 hold43/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X808 VPWR comp0.B\[1\] hold54/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X809 VGND hold54/a_285_47# hold54/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X810 net201 hold54/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X811 VGND comp0.B\[1\] hold54/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X812 VPWR hold54/a_285_47# hold54/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X813 hold54/a_285_47# hold54/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X814 hold54/a_285_47# hold54/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X815 net201 hold54/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X816 VPWR net65 hold65/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X817 VGND hold65/a_285_47# hold65/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X818 net212 hold65/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X819 VGND net65 hold65/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X820 VPWR hold65/a_285_47# hold65/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X821 hold65/a_285_47# hold65/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X822 hold65/a_285_47# hold65/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X823 net212 hold65/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X824 VPWR net46 hold76/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X825 VGND hold76/a_285_47# hold76/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X826 net223 hold76/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X827 VGND net46 hold76/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X828 VPWR hold76/a_285_47# hold76/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X829 hold76/a_285_47# hold76/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X830 hold76/a_285_47# hold76/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X831 net223 hold76/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X832 VPWR net36 hold87/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X833 VGND hold87/a_285_47# hold87/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X834 net234 hold87/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X835 VGND net36 hold87/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X836 VPWR hold87/a_285_47# hold87/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X837 hold87/a_285_47# hold87/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X838 hold87/a_285_47# hold87/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X839 net234 hold87/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X840 VPWR net40 hold98/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X841 VGND hold98/a_285_47# hold98/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X842 net245 hold98/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X843 VGND net40 hold98/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X844 VPWR hold98/a_285_47# hold98/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X845 hold98/a_285_47# hold98/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X846 hold98/a_285_47# hold98/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X847 net245 hold98/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X848 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X849 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X850 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X851 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X852 net48 _1002_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X853 _1002_/a_891_413# _1002_/a_193_47# _1002_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X854 _1002_/a_561_413# _1002_/a_27_47# _1002_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X855 VPWR net88 _1002_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X856 net48 _1002_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X857 _1002_/a_381_47# _0100_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X858 VGND _1002_/a_634_159# _1002_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X859 VPWR _1002_/a_891_413# _1002_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X860 _1002_/a_466_413# _1002_/a_193_47# _1002_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X861 VPWR _1002_/a_634_159# _1002_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X862 _1002_/a_634_159# _1002_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X863 _1002_/a_634_159# _1002_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X864 _1002_/a_975_413# _1002_/a_193_47# _1002_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X865 VGND _1002_/a_1059_315# _1002_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X866 _1002_/a_193_47# _1002_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X867 _1002_/a_891_413# _1002_/a_27_47# _1002_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X868 _1002_/a_592_47# _1002_/a_193_47# _1002_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X869 VPWR _1002_/a_1059_315# _1002_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X870 _1002_/a_1017_47# _1002_/a_27_47# _1002_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X871 _1002_/a_193_47# _1002_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X872 _1002_/a_466_413# _1002_/a_27_47# _1002_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X873 VGND _1002_/a_891_413# _1002_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X874 _1002_/a_381_47# _0100_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X875 VGND net88 _1002_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X876 _0648_/a_27_297# _0277_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X877 _0648_/a_27_297# _0279_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X878 _0648_/a_277_297# _0277_ _0648_/a_205_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X879 VPWR _0276_ _0648_/a_277_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X880 _0280_ _0648_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10187 ps=0.99 w=0.65 l=0.15
X881 _0648_/a_205_297# _0278_ _0648_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X882 _0280_ _0648_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X883 VGND _0278_ _0648_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X884 _0648_/a_109_297# _0279_ _0648_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X885 VGND _0276_ _0648_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X886 VPWR _0717_/a_80_21# _0348_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X887 _0717_/a_209_297# _0334_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X888 _0717_/a_303_47# _0333_ _0717_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X889 _0717_/a_209_47# _0334_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.11213 ps=0.995 w=0.65 l=0.15
X890 VGND _0717_/a_80_21# _0348_ VGND sky130_fd_pr__nfet_01v8 ad=0.11213 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X891 VGND _0335_ _0717_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X892 _0717_/a_80_21# _0221_ _0717_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X893 VPWR _0333_ _0717_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X894 _0717_/a_80_21# _0335_ _0717_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X895 _0717_/a_209_297# _0221_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X896 VPWR _0183_ _0579_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X897 _0579_/a_27_297# _0217_ _0579_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X898 VGND _0183_ _0579_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X899 _0118_ _0579_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X900 _0579_/a_27_297# _0217_ _0579_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X901 _0579_/a_109_297# net187 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X902 _0579_/a_373_47# net187 _0579_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X903 _0118_ _0579_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X904 _0579_/a_109_297# net211 _0579_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X905 _0579_/a_109_47# net211 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X906 VPWR output55/a_27_47# pp[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X907 pp[27] output55/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X908 VPWR net55 output55/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X909 pp[27] output55/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X910 VGND output55/a_27_47# pp[27] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X911 VGND net55 output55/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X912 VPWR output44/a_27_47# pp[17] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X913 pp[17] output44/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X914 VPWR net44 output44/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X915 pp[17] output44/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X916 VGND output44/a_27_47# pp[17] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X917 VGND net44 output44/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X918 VPWR net66 output66/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X919 VGND output66/a_27_47# pp[8] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X920 VGND output66/a_27_47# pp[8] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X921 pp[8] output66/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X922 pp[8] output66/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X923 VGND net66 output66/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X924 VPWR output66/a_27_47# pp[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X925 pp[8] output66/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X926 pp[8] output66/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X927 VPWR output66/a_27_47# pp[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X928 net68 clknet_1_0__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X929 VGND clknet_1_0__leaf__0458_ net68 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X930 net68 clknet_1_0__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X931 VPWR clknet_1_0__leaf__0458_ net68 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X934 VPWR _0180_ _0502_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X935 VGND _0502_/a_27_47# _0181_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X936 VGND _0502_/a_27_47# _0181_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X937 _0181_ _0502_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X938 _0181_ _0502_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X939 VGND _0180_ _0502_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X940 VPWR _0502_/a_27_47# _0181_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X941 _0181_ _0502_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X942 _0181_ _0502_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X943 VPWR _0502_/a_27_47# _0181_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X944 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X945 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X946 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X947 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X948 net93 clknet_1_1__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X949 VGND clknet_1_1__leaf__0460_ net93 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X950 net93 clknet_1_1__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X951 VPWR clknet_1_1__leaf__0460_ net93 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X952 net36 _0982_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X953 _0982_/a_891_413# _0982_/a_193_47# _0982_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X954 _0982_/a_561_413# _0982_/a_27_47# _0982_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X955 VPWR net68 _0982_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X956 net36 _0982_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X957 _0982_/a_381_47# _0080_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X958 VGND _0982_/a_634_159# _0982_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X959 VPWR _0982_/a_891_413# _0982_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X960 _0982_/a_466_413# _0982_/a_193_47# _0982_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X961 VPWR _0982_/a_634_159# _0982_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X962 _0982_/a_634_159# _0982_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X963 _0982_/a_634_159# _0982_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X964 _0982_/a_975_413# _0982_/a_193_47# _0982_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X965 VGND _0982_/a_1059_315# _0982_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X966 _0982_/a_193_47# _0982_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X967 _0982_/a_891_413# _0982_/a_27_47# _0982_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X968 _0982_/a_592_47# _0982_/a_193_47# _0982_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X969 VPWR _0982_/a_1059_315# _0982_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X970 _0982_/a_1017_47# _0982_/a_27_47# _0982_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X971 _0982_/a_193_47# _0982_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X972 _0982_/a_466_413# _0982_/a_27_47# _0982_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X973 VGND _0982_/a_891_413# _0982_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X974 _0982_/a_381_47# _0080_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X975 VGND net68 _0982_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X977 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X978 _0965_/a_377_297# control0.count\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X979 _0965_/a_47_47# _0478_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X980 _0965_/a_129_47# _0478_ _0965_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X981 _0965_/a_285_47# _0478_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X982 _0483_ _0965_/a_47_47# _0965_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X983 VGND control0.count\[3\] _0965_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X984 VPWR control0.count\[3\] _0965_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X985 VPWR _0965_/a_47_47# _0483_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X986 _0483_ _0478_ _0965_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X987 _0965_/a_285_47# control0.count\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X988 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X989 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X990 VPWR acc0.A\[25\] _0313_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X991 _0313_ acc0.A\[25\] _0681_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X992 _0681_/a_113_47# net53 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X993 _0313_ net53 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X996 VPWR _0226_ _0750_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2415 ps=2.83 w=0.42 l=0.15
X997 VPWR _0373_ _0750_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X998 _0750_/a_181_47# _0229_ _0750_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0882 pd=1.26 as=0.0882 ps=1.26 w=0.42 l=0.15
X999 VGND _0373_ _0750_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1000 _0750_/a_27_47# _0229_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1001 _0374_ _0750_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1002 _0374_ _0750_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1003 _0750_/a_109_47# _0226_ _0750_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1006 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1007 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1008 VPWR net34 _0948_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1009 VGND net34 _0468_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1010 _0948_/a_109_297# control0.state\[2\] _0468_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1011 _0468_ control0.state\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1012 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1013 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1016 VPWR _0414_ _0802_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1017 _0415_ _0802_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X1018 VGND _0414_ _0802_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1019 _0802_/a_59_75# _0404_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1020 _0415_ _0802_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X1021 _0802_/a_145_75# _0404_ _0802_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X1022 VPWR _0281_ _0664_/a_382_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.305 ps=2.61 w=1 l=0.15
X1023 _0664_/a_297_47# _0285_ _0664_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.3705 pd=3.74 as=0.169 ps=1.82 w=0.65 l=0.15
X1024 _0664_/a_297_47# _0281_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1025 VGND _0284_ _0664_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1026 VPWR _0664_/a_79_21# _0296_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X1027 _0664_/a_79_21# _0285_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.15
X1028 _0664_/a_382_297# _0284_ _0664_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1029 VGND _0664_/a_79_21# _0296_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1030 _0733_/a_222_93# _0319_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1031 VPWR _0321_ _0733_/a_544_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X1032 VGND _0733_/a_79_199# _0361_ VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1033 _0733_/a_222_93# _0319_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X1034 VGND _0360_ _0733_/a_448_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1035 _0733_/a_448_47# _0733_/a_222_93# _0733_/a_79_199# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1036 _0733_/a_79_199# _0733_/a_222_93# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X1037 _0733_/a_544_297# _0360_ _0733_/a_79_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1038 _0733_/a_448_47# _0321_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1039 VPWR _0733_/a_79_199# _0361_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
X1040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1042 VPWR acc0.A\[21\] _0595_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1043 VGND acc0.A\[21\] _0227_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1044 _0595_/a_109_297# net49 _0227_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1045 _0227_ net49 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1046 VPWR _0144_ hold11/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1047 VGND hold11/a_285_47# hold11/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1048 net158 hold11/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1049 VGND _0144_ hold11/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1050 VPWR hold11/a_285_47# hold11/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1051 hold11/a_285_47# hold11/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1052 hold11/a_285_47# hold11/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1053 net158 hold11/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1054 VPWR _0152_ hold22/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1055 VGND hold22/a_285_47# hold22/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1056 net169 hold22/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1057 VGND _0152_ hold22/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1058 VPWR hold22/a_285_47# hold22/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1059 hold22/a_285_47# hold22/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1060 hold22/a_285_47# hold22/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1061 net169 hold22/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1062 VPWR comp0.B\[8\] hold33/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1063 VGND hold33/a_285_47# hold33/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1064 net180 hold33/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1065 VGND comp0.B\[8\] hold33/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1066 VPWR hold33/a_285_47# hold33/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1067 hold33/a_285_47# hold33/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1068 hold33/a_285_47# hold33/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1069 net180 hold33/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1070 VPWR _0127_ hold44/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1071 VGND hold44/a_285_47# hold44/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1072 net191 hold44/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1073 VGND _0127_ hold44/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1074 VPWR hold44/a_285_47# hold44/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1075 hold44/a_285_47# hold44/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1076 hold44/a_285_47# hold44/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1077 net191 hold44/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1078 VPWR _0130_ hold55/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1079 VGND hold55/a_285_47# hold55/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1080 net202 hold55/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1081 VGND _0130_ hold55/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1082 VPWR hold55/a_285_47# hold55/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1083 hold55/a_285_47# hold55/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1084 hold55/a_285_47# hold55/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1085 net202 hold55/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1086 VPWR net49 hold66/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1087 VGND hold66/a_285_47# hold66/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1088 net213 hold66/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1089 VGND net49 hold66/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1090 VPWR hold66/a_285_47# hold66/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1091 hold66/a_285_47# hold66/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1092 hold66/a_285_47# hold66/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1093 net213 hold66/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1094 VPWR net55 hold77/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1095 VGND hold77/a_285_47# hold77/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1096 net224 hold77/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1097 VGND net55 hold77/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1098 VPWR hold77/a_285_47# hold77/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1099 hold77/a_285_47# hold77/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1100 hold77/a_285_47# hold77/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1101 net224 hold77/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1102 VPWR net64 hold88/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1103 VGND hold88/a_285_47# hold88/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1104 net235 hold88/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1105 VGND net64 hold88/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1106 VPWR hold88/a_285_47# hold88/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1107 hold88/a_285_47# hold88/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1108 hold88/a_285_47# hold88/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1109 net235 hold88/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1110 VPWR net38 hold99/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1111 VGND hold99/a_285_47# hold99/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1112 net246 hold99/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1113 VGND net38 hold99/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1114 VPWR hold99/a_285_47# hold99/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1115 hold99/a_285_47# hold99/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1116 hold99/a_285_47# hold99/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1117 net246 hold99/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1120 net46 _1001_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1121 _1001_/a_891_413# _1001_/a_193_47# _1001_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1122 _1001_/a_561_413# _1001_/a_27_47# _1001_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1123 VPWR net87 _1001_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1124 net46 _1001_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1125 _1001_/a_381_47# _0099_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1126 VGND _1001_/a_634_159# _1001_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1127 VPWR _1001_/a_891_413# _1001_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1128 _1001_/a_466_413# _1001_/a_193_47# _1001_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1129 VPWR _1001_/a_634_159# _1001_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1130 _1001_/a_634_159# _1001_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1131 _1001_/a_634_159# _1001_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1132 _1001_/a_975_413# _1001_/a_193_47# _1001_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1133 VGND _1001_/a_1059_315# _1001_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1134 _1001_/a_193_47# _1001_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1135 _1001_/a_891_413# _1001_/a_27_47# _1001_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1136 _1001_/a_592_47# _1001_/a_193_47# _1001_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1137 VPWR _1001_/a_1059_315# _1001_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1138 _1001_/a_1017_47# _1001_/a_27_47# _1001_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1139 _1001_/a_193_47# _1001_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1140 _1001_/a_466_413# _1001_/a_27_47# _1001_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1141 VGND _1001_/a_891_413# _1001_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1142 _1001_/a_381_47# _0099_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1143 VGND net87 _1001_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1144 VPWR _0346_ _0716_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1145 VGND _0716_/a_27_47# _0347_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1146 VGND _0716_/a_27_47# _0347_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1147 _0347_ _0716_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1148 _0347_ _0716_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1149 VGND _0346_ _0716_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1150 VPWR _0716_/a_27_47# _0347_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1151 _0347_ _0716_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1152 _0347_ _0716_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1153 VPWR _0716_/a_27_47# _0347_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1158 VPWR _0183_ _0578_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1159 _0578_/a_27_297# _0217_ _0578_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1160 VGND _0183_ _0578_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1161 _0119_ _0578_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1162 _0578_/a_27_297# _0217_ _0578_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1163 _0578_/a_109_297# net150 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1164 _0578_/a_373_47# net150 _0578_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1165 _0119_ _0578_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1166 _0578_/a_109_297# net187 _0578_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1167 _0578_/a_109_47# net187 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1168 _0647_/a_377_297# acc0.A\[12\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X1169 _0647_/a_47_47# net39 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1170 _0647_/a_129_47# net39 _0647_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X1171 _0647_/a_285_47# net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X1172 _0279_ _0647_/a_47_47# _0647_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X1173 VGND acc0.A\[12\] _0647_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1174 VPWR acc0.A\[12\] _0647_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1175 VPWR _0647_/a_47_47# _0279_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X1176 _0279_ net39 _0647_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1177 _0647_/a_285_47# acc0.A\[12\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1182 VPWR output56/a_27_47# pp[28] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1183 pp[28] output56/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1184 VPWR net56 output56/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1185 pp[28] output56/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1186 VGND output56/a_27_47# pp[28] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1187 VGND net56 output56/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1188 VPWR output45/a_27_47# pp[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1189 pp[18] output45/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1190 VPWR net45 output45/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1191 pp[18] output45/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1192 VGND output45/a_27_47# pp[18] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1193 VGND net45 output45/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1194 VPWR net67 output67/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1195 VGND output67/a_27_47# pp[9] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1196 VGND output67/a_27_47# pp[9] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1197 pp[9] output67/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1198 pp[9] output67/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1199 VGND net67 output67/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1200 VPWR output67/a_27_47# pp[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1201 pp[9] output67/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1202 pp[9] output67/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1203 VPWR output67/a_27_47# pp[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1204 VPWR _0501_/a_27_47# _0180_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1205 _0180_ _0501_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1206 VPWR control0.reset _0501_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1207 _0180_ _0501_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1208 VGND _0501_/a_27_47# _0180_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1209 VGND control0.reset _0501_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1212 net70 clknet_1_0__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1213 VGND clknet_1_0__leaf__0458_ net70 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1214 net70 clknet_1_0__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1215 VPWR clknet_1_0__leaf__0458_ net70 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1216 VPWR _0466_ _0981_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1217 _0981_/a_27_297# _0490_ _0981_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1218 VGND _0466_ _0981_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1219 _0170_ _0981_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1220 _0981_/a_27_297# _0490_ _0981_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1221 _0981_/a_109_297# net167 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1222 _0981_/a_373_47# net167 _0981_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1223 _0170_ _0981_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1224 _0981_/a_109_297# _0488_ _0981_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1225 _0981_/a_109_47# _0488_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1226 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1230 VPWR _0480_ _0964_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1231 VGND _0480_ _0482_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1232 _0964_/a_109_297# _0481_ _0482_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1233 _0482_ _0481_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1234 net131 clknet_1_1__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1235 VGND clknet_1_1__leaf__0464_ net131 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1236 net131 clknet_1_1__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1237 VPWR clknet_1_1__leaf__0464_ net131 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1238 net145 clknet_1_1__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1239 VGND clknet_1_1__leaf__0465_ net145 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1240 net145 clknet_1_1__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1241 VPWR clknet_1_1__leaf__0465_ net145 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1244 VPWR _0680_/a_80_21# _0312_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1245 _0680_/a_80_21# _0238_ _0680_/a_472_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1246 VPWR _0305_ _0680_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1247 VGND _0311_ _0680_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X1248 VGND _0680_/a_80_21# _0312_ VGND sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X1249 _0680_/a_300_47# _0305_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X1250 _0680_/a_217_297# _0294_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1251 _0680_/a_80_21# _0294_ _0680_/a_300_47# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1252 _0680_/a_472_297# _0311_ _0680_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X1253 _0680_/a_80_21# _0238_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X1254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1256 net78 clknet_1_1__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1257 VGND clknet_1_1__leaf__0459_ net78 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1258 net78 clknet_1_1__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1259 VPWR clknet_1_1__leaf__0459_ net78 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1260 VPWR control0.state\[2\] _0947_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1261 VGND control0.state\[2\] _0467_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1262 _0947_/a_109_297# _0466_ _0467_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1263 _0467_ _0466_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1264 VPWR clknet_1_0__leaf_clk clkload0/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1265 VGND clkload0/a_27_47# clkload0/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1266 VGND clkload0/a_27_47# clkload0/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1267 clkload0/X clkload0/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1268 clkload0/X clkload0/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1269 VGND clknet_1_0__leaf_clk clkload0/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1270 VPWR clkload0/a_27_47# clkload0/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1271 clkload0/X clkload0/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1272 clkload0/X clkload0/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1273 VPWR clkload0/a_27_47# clkload0/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1280 VPWR _0279_ _0414_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1281 _0414_ _0279_ _0801_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1282 _0801_/a_113_47# _0403_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1283 _0414_ _0403_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1286 VPWR _0290_ _0663_/a_207_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1287 _0295_ _0663_/a_207_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X1288 _0663_/a_297_47# _0663_/a_27_413# _0663_/a_207_413# VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X1289 _0295_ _0663_/a_207_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1290 _0663_/a_207_413# _0663_/a_27_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1291 VPWR _0288_ _0663_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1292 VGND _0290_ _0663_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1293 _0663_/a_27_413# _0288_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1294 VPWR _0732_/a_80_21# _0360_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1295 _0732_/a_209_297# _0313_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.65 pd=5.3 as=0 ps=0 w=1 l=0.15
X1296 _0732_/a_303_47# _0359_ _0732_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.208 ps=1.94 w=0.65 l=0.15
X1297 _0732_/a_209_47# _0313_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1298 VGND _0732_/a_80_21# _0360_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X1299 VGND _0328_ _0732_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X1300 _0732_/a_80_21# _0324_ _0732_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1301 VPWR _0359_ _0732_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1302 _0732_/a_80_21# _0328_ _0732_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0 ps=0 w=1 l=0.15
X1303 _0732_/a_209_297# _0324_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1304 VPWR acc0.A\[20\] _0226_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1305 _0226_ acc0.A\[20\] _0594_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1306 _0594_/a_113_47# net48 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1307 _0226_ net48 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1312 net112 clknet_1_0__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1313 VGND clknet_1_0__leaf__0462_ net112 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1314 net112 clknet_1_0__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1315 VPWR clknet_1_0__leaf__0462_ net112 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1318 net126 clknet_1_0__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1319 VGND clknet_1_0__leaf__0463_ net126 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1320 net126 clknet_1_0__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1321 VPWR clknet_1_0__leaf__0463_ net126 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1322 VPWR net35 hold12/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1323 VGND hold12/a_285_47# hold12/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1324 net159 hold12/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1325 VGND net35 hold12/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1326 VPWR hold12/a_285_47# hold12/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1327 hold12/a_285_47# hold12/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1328 hold12/a_285_47# hold12/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1329 net159 hold12/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1330 VPWR acc0.A\[3\] hold23/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1331 VGND hold23/a_285_47# hold23/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1332 net170 hold23/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1333 VGND acc0.A\[3\] hold23/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1334 VPWR hold23/a_285_47# hold23/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1335 hold23/a_285_47# hold23/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1336 hold23/a_285_47# hold23/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1337 net170 hold23/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1338 VPWR acc0.A\[9\] hold34/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1339 VGND hold34/a_285_47# hold34/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1340 net181 hold34/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1341 VGND acc0.A\[9\] hold34/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1342 VPWR hold34/a_285_47# hold34/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1343 hold34/a_285_47# hold34/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1344 hold34/a_285_47# hold34/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1345 net181 hold34/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1346 VPWR acc0.A\[11\] hold45/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1347 VGND hold45/a_285_47# hold45/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1348 net192 hold45/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1349 VGND acc0.A\[11\] hold45/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1350 VPWR hold45/a_285_47# hold45/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1351 hold45/a_285_47# hold45/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1352 hold45/a_285_47# hold45/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1353 net192 hold45/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1354 VPWR comp0.B\[2\] hold56/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1355 VGND hold56/a_285_47# hold56/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1356 net203 hold56/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1357 VGND comp0.B\[2\] hold56/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1358 VPWR hold56/a_285_47# hold56/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1359 hold56/a_285_47# hold56/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1360 hold56/a_285_47# hold56/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1361 net203 hold56/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1362 VPWR net66 hold67/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1363 VGND hold67/a_285_47# hold67/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1364 net214 hold67/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1365 VGND net66 hold67/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1366 VPWR hold67/a_285_47# hold67/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1367 hold67/a_285_47# hold67/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1368 hold67/a_285_47# hold67/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1369 net214 hold67/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1370 VPWR net60 hold78/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1371 VGND hold78/a_285_47# hold78/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1372 net225 hold78/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1373 VGND net60 hold78/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1374 VPWR hold78/a_285_47# hold78/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1375 hold78/a_285_47# hold78/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1376 hold78/a_285_47# hold78/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1377 net225 hold78/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1378 VPWR control0.state\[2\] hold89/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1379 VGND hold89/a_285_47# hold89/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1380 net236 hold89/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1381 VGND control0.state\[2\] hold89/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1382 VPWR hold89/a_285_47# hold89/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1383 hold89/a_285_47# hold89/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1384 hold89/a_285_47# hold89/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1385 net236 hold89/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1386 net45 _1000_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1387 _1000_/a_891_413# _1000_/a_193_47# _1000_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1388 _1000_/a_561_413# _1000_/a_27_47# _1000_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1389 VPWR net86 _1000_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1390 net45 _1000_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1391 _1000_/a_381_47# _0098_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1392 VGND _1000_/a_634_159# _1000_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1393 VPWR _1000_/a_891_413# _1000_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1394 _1000_/a_466_413# _1000_/a_193_47# _1000_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1395 VPWR _1000_/a_634_159# _1000_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1396 _1000_/a_634_159# _1000_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1397 _1000_/a_634_159# _1000_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1398 _1000_/a_975_413# _1000_/a_193_47# _1000_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1399 VGND _1000_/a_1059_315# _1000_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1400 _1000_/a_193_47# _1000_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1401 _1000_/a_891_413# _1000_/a_27_47# _1000_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1402 _1000_/a_592_47# _1000_/a_193_47# _1000_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1403 VPWR _1000_/a_1059_315# _1000_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1404 _1000_/a_1017_47# _1000_/a_27_47# _1000_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1405 _1000_/a_193_47# _1000_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1406 _1000_/a_466_413# _1000_/a_27_47# _1000_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1407 VGND _1000_/a_891_413# _1000_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1408 _1000_/a_381_47# _0098_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1409 VGND net86 _1000_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1410 VPWR _0343_ _0715_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1411 VGND _0715_/a_27_47# _0346_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1412 VGND _0715_/a_27_47# _0346_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1413 _0346_ _0715_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1414 _0346_ _0715_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1415 VGND _0343_ _0715_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1416 VPWR _0715_/a_27_47# _0346_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1417 _0346_ _0715_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1418 _0346_ _0715_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1419 VPWR _0715_/a_27_47# _0346_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1422 VPWR _0183_ _0577_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1423 _0577_/a_27_297# _0217_ _0577_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1424 VGND _0183_ _0577_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1425 _0120_ _0577_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1426 _0577_/a_27_297# _0217_ _0577_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1427 _0577_/a_109_297# acc0.A\[22\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1428 _0577_/a_373_47# acc0.A\[22\] _0577_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1429 _0120_ _0577_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1430 _0577_/a_109_297# net150 _0577_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1431 _0577_/a_109_47# net150 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1432 _0646_/a_377_297# acc0.A\[13\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X1433 _0646_/a_47_47# net40 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1434 _0646_/a_129_47# net40 _0646_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X1435 _0646_/a_285_47# net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X1436 _0278_ _0646_/a_47_47# _0646_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X1437 VGND acc0.A\[13\] _0646_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1438 VPWR acc0.A\[13\] _0646_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1439 VPWR _0646_/a_47_47# _0278_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X1440 _0278_ net40 _0646_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1441 _0646_/a_285_47# acc0.A\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1444 VPWR output57/a_27_47# pp[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1445 pp[29] output57/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1446 VPWR net57 output57/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1447 pp[29] output57/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1448 VGND output57/a_27_47# pp[29] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1449 VGND net57 output57/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1450 VPWR output46/a_27_47# pp[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1451 pp[19] output46/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1452 VPWR net46 output46/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1453 pp[19] output46/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1454 VGND output46/a_27_47# pp[19] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1455 VGND net46 output46/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1456 VPWR output35/a_27_47# done VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1457 done output35/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1458 VPWR net35 output35/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1459 done output35/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1460 VGND output35/a_27_47# done VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1461 VGND net35 output35/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1464 VPWR _0178_ _0500_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1465 VGND _0500_/a_27_47# _0179_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1466 VGND _0500_/a_27_47# _0179_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1467 _0179_ _0500_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1468 _0179_ _0500_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1469 VGND _0178_ _0500_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1470 VPWR _0500_/a_27_47# _0179_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1471 _0179_ _0500_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1472 _0179_ _0500_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1473 VPWR _0500_/a_27_47# _0179_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1480 VPWR net58 _0629_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1481 _0261_ _0629_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X1482 VGND net58 _0629_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1483 _0629_/a_59_75# acc0.A\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1484 _0261_ _0629_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X1485 _0629_/a_145_75# acc0.A\[2\] _0629_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X1486 _0490_ _0483_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1487 VGND _0483_ _0490_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1488 _0490_ _0483_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1489 VPWR _0483_ _0490_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1502 _0481_ _0963_/a_35_297# _0963_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1503 _0481_ control0.count\[0\] _0963_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X1504 _0963_/a_35_297# control0.count\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1505 _0963_/a_117_297# control0.count\[0\] _0963_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1506 VPWR control0.count\[0\] _0963_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1507 VGND control0.count\[1\] _0963_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1508 VGND _0963_/a_35_297# _0481_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X1509 _0963_/a_285_297# control0.count\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1510 VPWR control0.count\[1\] _0963_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1511 _0963_/a_285_47# control0.count\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1514 VPWR _0946_/a_30_53# _0466_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1515 VGND _0946_/a_30_53# _0466_ VGND sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X1516 _0466_ _0946_/a_30_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X1517 _0946_/a_112_297# control0.state\[0\] _0946_/a_30_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1518 _0466_ _0946_/a_30_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10187 ps=0.99 w=0.65 l=0.15
X1519 VGND net34 _0946_/a_30_53# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1520 _0946_/a_30_53# control0.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1521 VGND control0.state\[0\] _0946_/a_30_53# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1522 _0946_/a_184_297# control0.state\[1\] _0946_/a_112_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1523 VPWR net34 _0946_/a_184_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1526 clkload1/Y clknet_1_0__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X1527 VGND clknet_1_0__leaf__0465_ clkload1/a_268_47# VGND sky130_fd_pr__nfet_01v8 ad=0.14575 pd=1.63 as=0.05775 ps=0.76 w=0.55 l=0.15
X1528 clkload1/Y clknet_1_0__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X1529 clkload1/Y clknet_1_0__leaf__0465_ clkload1/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.077 pd=0.83 as=0.05775 ps=0.76 w=0.55 l=0.15
X1530 VPWR clknet_1_0__leaf__0465_ clkload1/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X1531 clkload1/a_110_47# clknet_1_0__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.14575 ps=1.63 w=0.55 l=0.15
X1532 clkload1/a_268_47# clknet_1_0__leaf__0465_ clkload1/Y VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.077 ps=0.83 w=0.55 l=0.15
X1533 VPWR clknet_1_0__leaf__0465_ clkload1/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X1534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1538 _0800_/a_240_47# net245 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1539 _0093_ _0800_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1540 VGND _0219_ _0800_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1541 _0800_/a_51_297# _0413_ _0800_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X1542 _0800_/a_149_47# _0345_ _0800_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.09912 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X1543 _0800_/a_240_47# _0412_ _0800_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09912 ps=0.955 w=0.65 l=0.15
X1544 VPWR _0219_ _0800_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X1545 _0093_ _0800_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X1546 _0800_/a_149_47# _0413_ _0800_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1547 _0800_/a_245_297# _0412_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1548 VPWR _0345_ _0800_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X1549 _0800_/a_512_297# net245 _0800_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
X1550 _0731_/a_81_21# _0326_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X1551 _0731_/a_299_297# _0326_ _0731_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X1552 VPWR _0731_/a_81_21# _0359_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1553 VPWR _0250_ _0731_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1554 VGND _0731_/a_81_21# _0359_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1555 VGND _0312_ _0731_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X1556 _0731_/a_299_297# _0312_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1557 _0731_/a_384_47# _0250_ _0731_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1558 VPWR _0222_ _0225_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1559 _0225_ _0222_ _0593_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1560 _0593_/a_113_47# _0224_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1561 _0225_ _0224_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1562 _0662_/a_81_21# _0293_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X1563 _0662_/a_299_297# _0293_ _0662_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X1564 VPWR _0662_/a_81_21# _0294_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1565 VPWR _0259_ _0662_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1566 VGND _0662_/a_81_21# _0294_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1567 VGND _0275_ _0662_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X1568 _0662_/a_299_297# _0275_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1569 _0662_/a_384_47# _0259_ _0662_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1574 VPWR comp0.B\[5\] hold13/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1575 VGND hold13/a_285_47# hold13/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1576 net160 hold13/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1577 VGND comp0.B\[5\] hold13/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1578 VPWR hold13/a_285_47# hold13/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1579 hold13/a_285_47# hold13/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1580 hold13/a_285_47# hold13/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1581 net160 hold13/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1582 VPWR comp0.B\[7\] hold24/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1583 VGND hold24/a_285_47# hold24/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1584 net171 hold24/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1585 VGND comp0.B\[7\] hold24/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1586 VPWR hold24/a_285_47# hold24/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1587 hold24/a_285_47# hold24/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1588 hold24/a_285_47# hold24/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1589 net171 hold24/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1590 VPWR _0154_ hold35/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1591 VGND hold35/a_285_47# hold35/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1592 net182 hold35/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1593 VGND _0154_ hold35/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1594 VPWR hold35/a_285_47# hold35/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1595 hold35/a_285_47# hold35/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1596 hold35/a_285_47# hold35/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1597 net182 hold35/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1598 VPWR comp0.B\[13\] hold46/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1599 VGND hold46/a_285_47# hold46/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1600 net193 hold46/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1601 VGND comp0.B\[13\] hold46/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1602 VPWR hold46/a_285_47# hold46/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1603 hold46/a_285_47# hold46/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1604 hold46/a_285_47# hold46/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1605 net193 hold46/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1606 VPWR comp0.B\[6\] hold57/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1607 VGND hold57/a_285_47# hold57/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1608 net204 hold57/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1609 VGND comp0.B\[6\] hold57/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1610 VPWR hold57/a_285_47# hold57/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1611 hold57/a_285_47# hold57/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1612 hold57/a_285_47# hold57/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1613 net204 hold57/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1614 VPWR acc0.A\[23\] hold68/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1615 VGND hold68/a_285_47# hold68/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1616 net215 hold68/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1617 VGND acc0.A\[23\] hold68/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1618 VPWR hold68/a_285_47# hold68/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1619 hold68/a_285_47# hold68/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1620 hold68/a_285_47# hold68/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1621 net215 hold68/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1622 VPWR control0.count\[1\] hold79/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1623 VGND hold79/a_285_47# hold79/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1624 net226 hold79/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1625 VGND control0.count\[1\] hold79/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1626 VPWR hold79/a_285_47# hold79/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1627 hold79/a_285_47# hold79/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1628 hold79/a_285_47# hold79/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1629 net226 hold79/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1632 _0714_/a_240_47# _0219_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X1633 _0111_ _0714_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X1634 VGND net225 _0714_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1635 _0714_/a_51_297# _0344_ _0714_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X1636 _0714_/a_149_47# _0345_ _0714_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X1637 _0714_/a_240_47# _0342_ _0714_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1638 VPWR net225 _0714_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1639 _0111_ _0714_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X1640 _0714_/a_149_47# _0344_ _0714_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1641 _0714_/a_245_297# _0342_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1642 VPWR _0345_ _0714_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1643 _0714_/a_512_297# _0219_ _0714_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1644 _0645_/a_377_297# acc0.A\[14\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X1645 _0645_/a_47_47# net41 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1646 _0645_/a_129_47# net41 _0645_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X1647 _0645_/a_285_47# net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X1648 _0277_ _0645_/a_47_47# _0645_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X1649 VGND acc0.A\[14\] _0645_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1650 VPWR acc0.A\[14\] _0645_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1651 VPWR _0645_/a_47_47# _0277_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X1652 _0277_ net41 _0645_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1653 _0645_/a_285_47# acc0.A\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1654 VPWR _0183_ _0576_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1655 _0576_/a_27_297# _0217_ _0576_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1656 VGND _0183_ _0576_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1657 _0121_ _0576_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1658 _0576_/a_27_297# _0217_ _0576_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1659 _0576_/a_109_297# acc0.A\[23\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1660 _0576_/a_373_47# acc0.A\[23\] _0576_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1661 _0121_ _0576_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1662 _0576_/a_109_297# net176 _0576_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1663 _0576_/a_109_47# net176 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1664 acc0.A\[13\] _1059_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1665 _1059_/a_891_413# _1059_/a_193_47# _1059_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1666 _1059_/a_561_413# _1059_/a_27_47# _1059_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1667 VPWR net145 _1059_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1668 acc0.A\[13\] _1059_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1669 _1059_/a_381_47# _0157_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1670 VGND _1059_/a_634_159# _1059_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1671 VPWR _1059_/a_891_413# _1059_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1672 _1059_/a_466_413# _1059_/a_193_47# _1059_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1673 VPWR _1059_/a_634_159# _1059_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1674 _1059_/a_634_159# _1059_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1675 _1059_/a_634_159# _1059_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1676 _1059_/a_975_413# _1059_/a_193_47# _1059_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1677 VGND _1059_/a_1059_315# _1059_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1678 _1059_/a_193_47# _1059_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1679 _1059_/a_891_413# _1059_/a_27_47# _1059_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1680 _1059_/a_592_47# _1059_/a_193_47# _1059_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1681 VPWR _1059_/a_1059_315# _1059_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1682 _1059_/a_1017_47# _1059_/a_27_47# _1059_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1683 _1059_/a_193_47# _1059_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1684 _1059_/a_466_413# _1059_/a_27_47# _1059_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1685 VGND _1059_/a_891_413# _1059_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1686 _1059_/a_381_47# _0157_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1687 VGND net145 _1059_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1690 VPWR output36/a_27_47# pp[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1691 pp[0] output36/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1692 VPWR net36 output36/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1693 pp[0] output36/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1694 VGND output36/a_27_47# pp[0] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1695 VGND net36 output36/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1696 VPWR net58 output58/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1697 VGND output58/a_27_47# pp[2] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1698 VGND output58/a_27_47# pp[2] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1699 pp[2] output58/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1700 pp[2] output58/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1701 VGND net58 output58/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1702 VPWR output58/a_27_47# pp[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1703 pp[2] output58/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1704 pp[2] output58/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1705 VPWR output58/a_27_47# pp[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1706 VPWR net47 output47/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1707 VGND output47/a_27_47# pp[1] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1708 VGND output47/a_27_47# pp[1] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1709 pp[1] output47/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1710 pp[1] output47/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1711 VGND net47 output47/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1712 VPWR output47/a_27_47# pp[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1713 pp[1] output47/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1714 pp[1] output47/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1715 VPWR output47/a_27_47# pp[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1718 net104 clknet_1_0__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1719 VGND clknet_1_0__leaf__0461_ net104 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1720 net104 clknet_1_0__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1721 VPWR clknet_1_0__leaf__0461_ net104 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1722 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1724 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1725 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1726 VPWR acc0.A\[3\] _0628_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1727 VGND acc0.A\[3\] _0260_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1728 _0628_/a_109_297# net61 _0260_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1729 _0260_ net61 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1730 _0559_/a_240_47# net26 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X1731 _0133_ _0559_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X1732 VGND _0208_ _0559_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1733 _0559_/a_51_297# net205 _0559_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X1734 _0559_/a_149_47# _0212_ _0559_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X1735 _0559_/a_240_47# _0173_ _0559_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1736 VPWR _0208_ _0559_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1737 _0133_ _0559_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X1738 _0559_/a_149_47# net205 _0559_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1739 _0559_/a_245_297# _0173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1740 VPWR _0212_ _0559_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1741 _0559_/a_512_297# net26 _0559_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1744 net85 clknet_1_1__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1745 VGND clknet_1_1__leaf__0459_ net85 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1746 net85 clknet_1_1__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1747 VPWR clknet_1_1__leaf__0459_ net85 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1750 VPWR _0478_ _0962_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1751 VGND _0478_ _0480_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1752 _0962_/a_109_297# _0479_ _0480_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1753 _0480_ _0479_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1754 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1755 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1762 clkload2/Y clknet_1_0__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.25
X1763 VGND clknet_1_0__leaf__0464_ clkload2/a_268_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1155 ps=1.52 w=0.55 l=0.15
X1764 clkload2/Y clknet_1_0__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X1765 clkload2/Y clknet_1_0__leaf__0464_ clkload2/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.154 pd=1.66 as=0.1155 ps=1.52 w=0.55 l=0.15
X1766 VPWR clknet_1_0__leaf__0464_ clkload2/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X1767 clkload2/a_110_47# clknet_1_0__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.15
X1768 clkload2/a_268_47# clknet_1_0__leaf__0464_ clkload2/Y VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.15
X1769 VPWR clknet_1_0__leaf__0464_ clkload2/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X1770 _0661_/a_27_297# _0288_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.252 pd=2.88 as=0 ps=0 w=0.42 l=0.15
X1771 _0661_/a_27_297# _0292_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1772 _0661_/a_277_297# _0288_ _0661_/a_205_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1386 pd=1.5 as=0.0882 ps=1.26 w=0.42 l=0.15
X1773 VPWR _0287_ _0661_/a_277_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1774 _0293_ _0661_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1775 _0661_/a_205_297# _0289_ _0661_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1386 ps=1.5 w=0.42 l=0.15
X1776 _0293_ _0661_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1777 VGND _0289_ _0661_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1778 _0661_/a_109_297# _0292_ _0661_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1779 VGND _0287_ _0661_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1780 VGND _0347_ _0730_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X1781 _0730_/a_510_47# _0358_ _0730_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X1782 _0730_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X1783 VPWR _0358_ _0730_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1784 _0730_/a_79_21# _0357_ _0730_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X1785 _0730_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1786 _0730_/a_79_21# _0352_ _0730_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X1787 VPWR _0730_/a_79_21# _0108_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1788 VGND _0730_/a_79_21# _0108_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1789 _0730_/a_215_47# _0357_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1790 VGND acc0.A\[22\] _0592_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1791 _0592_/a_68_297# net50 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1792 _0224_ _0592_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1793 VPWR acc0.A\[22\] _0592_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X1794 _0224_ _0592_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X1795 _0592_/a_150_297# net50 _0592_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1798 VPWR _0134_ hold14/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1799 VGND hold14/a_285_47# hold14/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1800 net161 hold14/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1801 VGND _0134_ hold14/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1802 VPWR hold14/a_285_47# hold14/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1803 hold14/a_285_47# hold14/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1804 hold14/a_285_47# hold14/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1805 net161 hold14/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1806 VPWR _0136_ hold25/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1807 VGND hold25/a_285_47# hold25/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1808 net172 hold25/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1809 VGND _0136_ hold25/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1810 VPWR hold25/a_285_47# hold25/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1811 hold25/a_285_47# hold25/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1812 hold25/a_285_47# hold25/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1813 net172 hold25/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1814 VPWR comp0.B\[14\] hold36/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1815 VGND hold36/a_285_47# hold36/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1816 net183 hold36/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1817 VGND comp0.B\[14\] hold36/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1818 VPWR hold36/a_285_47# hold36/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1819 hold36/a_285_47# hold36/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1820 hold36/a_285_47# hold36/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1821 net183 hold36/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1822 VPWR _0142_ hold47/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1823 VGND hold47/a_285_47# hold47/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1824 net194 hold47/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1825 VGND _0142_ hold47/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1826 VPWR hold47/a_285_47# hold47/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1827 hold47/a_285_47# hold47/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1828 hold47/a_285_47# hold47/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1829 net194 hold47/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1830 VPWR comp0.B\[4\] hold58/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1831 VGND hold58/a_285_47# hold58/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1832 net205 hold58/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1833 VGND comp0.B\[4\] hold58/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1834 VPWR hold58/a_285_47# hold58/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1835 hold58/a_285_47# hold58/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1836 hold58/a_285_47# hold58/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1837 net205 hold58/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1838 VPWR net52 hold69/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1839 VGND hold69/a_285_47# hold69/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1840 net216 hold69/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1841 VGND net52 hold69/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1842 VPWR hold69/a_285_47# hold69/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1843 hold69/a_285_47# hold69/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1844 hold69/a_285_47# hold69/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1845 net216 hold69/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1846 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1847 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1848 net117 clknet_1_1__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1849 VGND clknet_1_1__leaf__0462_ net117 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1850 net117 clknet_1_1__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1851 VPWR clknet_1_1__leaf__0462_ net117 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1852 VPWR _0208_ _0713_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1853 VGND _0713_/a_27_47# _0345_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1854 VGND _0713_/a_27_47# _0345_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1855 _0345_ _0713_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1856 _0345_ _0713_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1857 VGND _0208_ _0713_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1858 VPWR _0713_/a_27_47# _0345_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1859 _0345_ _0713_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1860 _0345_ _0713_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1861 VPWR _0713_/a_27_47# _0345_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1862 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1863 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1864 _0644_/a_377_297# acc0.A\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X1865 _0644_/a_47_47# net42 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1866 _0644_/a_129_47# net42 _0644_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X1867 _0644_/a_285_47# net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X1868 _0276_ _0644_/a_47_47# _0644_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X1869 VGND acc0.A\[15\] _0644_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1870 VPWR acc0.A\[15\] _0644_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1871 VPWR _0644_/a_47_47# _0276_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X1872 _0276_ net42 _0644_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1873 _0644_/a_285_47# acc0.A\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1874 VPWR _0216_ _0575_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1875 _0575_/a_27_297# _0217_ _0575_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1876 VGND _0216_ _0575_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1877 _0122_ _0575_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1878 _0575_/a_27_297# _0217_ _0575_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1879 _0575_/a_109_297# net199 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1880 _0575_/a_373_47# net199 _0575_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1881 _0122_ _0575_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1882 _0575_/a_109_297# net215 _0575_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1883 _0575_/a_109_47# net215 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1884 acc0.A\[12\] _1058_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1885 _1058_/a_891_413# _1058_/a_193_47# _1058_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1886 _1058_/a_561_413# _1058_/a_27_47# _1058_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1887 VPWR net144 _1058_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1888 acc0.A\[12\] _1058_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1889 _1058_/a_381_47# _0156_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1890 VGND _1058_/a_634_159# _1058_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1891 VPWR _1058_/a_891_413# _1058_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1892 _1058_/a_466_413# _1058_/a_193_47# _1058_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1893 VPWR _1058_/a_634_159# _1058_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1894 _1058_/a_634_159# _1058_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1895 _1058_/a_634_159# _1058_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1896 _1058_/a_975_413# _1058_/a_193_47# _1058_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1897 VGND _1058_/a_1059_315# _1058_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1898 _1058_/a_193_47# _1058_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1899 _1058_/a_891_413# _1058_/a_27_47# _1058_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1900 _1058_/a_592_47# _1058_/a_193_47# _1058_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1901 VPWR _1058_/a_1059_315# _1058_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1902 _1058_/a_1017_47# _1058_/a_27_47# _1058_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1903 _1058_/a_193_47# _1058_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1904 _1058_/a_466_413# _1058_/a_27_47# _1058_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1905 VGND _1058_/a_891_413# _1058_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1906 _1058_/a_381_47# _0156_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1907 VGND net144 _1058_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1908 VPWR output59/a_27_47# pp[30] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1909 pp[30] output59/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1910 VPWR net59 output59/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1911 pp[30] output59/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1912 VGND output59/a_27_47# pp[30] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1913 VGND net59 output59/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1914 VPWR output48/a_27_47# pp[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1915 pp[20] output48/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1916 VPWR net48 output48/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1917 pp[20] output48/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1918 VGND output48/a_27_47# pp[20] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1919 VGND net48 output48/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1920 VPWR net37 output37/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1921 VGND output37/a_27_47# pp[10] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1922 VGND output37/a_27_47# pp[10] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1923 pp[10] output37/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1924 pp[10] output37/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1925 VGND net37 output37/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1926 VPWR output37/a_27_47# pp[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1927 pp[10] output37/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1928 pp[10] output37/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1929 VPWR output37/a_27_47# pp[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1934 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1935 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1936 _0627_/a_109_93# _0258_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1937 _0627_/a_215_53# _0255_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1938 VGND _0627_/a_109_93# _0627_/a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1939 VGND _0254_ _0627_/a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1940 VPWR _0254_ _0627_/a_369_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1941 _0627_/a_369_297# _0255_ _0627_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X1942 _0259_ _0627_/a_215_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1943 _0627_/a_297_297# _0627_/a_109_93# _0627_/a_215_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1944 _0627_/a_109_93# _0258_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1945 _0259_ _0627_/a_215_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X1946 VGND net185 _0558_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1947 _0558_/a_68_297# _0175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1948 _0212_ _0558_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1949 VPWR net185 _0558_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X1950 _0212_ _0558_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X1951 _0558_/a_150_297# _0175_ _0558_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1954 VPWR acc0.A\[14\] hold100/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1955 VGND hold100/a_285_47# hold100/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1956 net247 hold100/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1957 VGND acc0.A\[14\] hold100/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1958 VPWR hold100/a_285_47# hold100/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1959 hold100/a_285_47# hold100/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1960 hold100/a_285_47# hold100/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1961 net247 hold100/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1964 net89 clknet_1_0__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1965 VGND clknet_1_0__leaf__0460_ net89 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1966 net89 clknet_1_0__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1967 VPWR clknet_1_0__leaf__0460_ net89 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1968 _0961_/a_199_47# control0.count\[1\] _0479_ VGND sky130_fd_pr__nfet_01v8 ad=0.09588 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1969 _0961_/a_113_297# control0.count\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X1970 _0479_ control0.count\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1971 VPWR control0.count\[1\] _0961_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X1972 _0961_/a_113_297# control0.count\[2\] _0479_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1973 VGND control0.count\[0\] _0961_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.09588 ps=0.945 w=0.65 l=0.15
X1974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1976 net123 clknet_1_0__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1977 VGND clknet_1_0__leaf__0463_ net123 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1978 net123 clknet_1_0__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1979 VPWR clknet_1_0__leaf__0463_ net123 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1984 clkload3/Y clknet_1_1__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.25
X1985 VGND clknet_1_1__leaf__0461_ clkload3/a_268_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1155 ps=1.52 w=0.55 l=0.15
X1986 clkload3/Y clknet_1_1__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X1987 clkload3/Y clknet_1_1__leaf__0461_ clkload3/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.154 pd=1.66 as=0.1155 ps=1.52 w=0.55 l=0.15
X1988 VPWR clknet_1_1__leaf__0461_ clkload3/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X1989 clkload3/a_110_47# clknet_1_1__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.15
X1990 clkload3/a_268_47# clknet_1_1__leaf__0461_ clkload3/Y VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.15
X1991 VPWR clknet_1_1__leaf__0461_ clkload3/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X1992 VPWR _0290_ _0292_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1993 _0292_ _0290_ _0660_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1994 _0660_/a_113_47# _0291_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1995 _0292_ _0291_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1996 VPWR acc0.A\[23\] _0591_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1997 VGND acc0.A\[23\] _0223_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1998 _0591_/a_109_297# net51 _0223_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1999 _0223_ net51 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2002 _0789_/a_75_199# _0277_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13487 ps=1.065 w=0.65 l=0.15
X2003 _0789_/a_208_47# _0404_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12513 pd=1.035 as=0.11213 ps=0.995 w=0.65 l=0.15
X2004 _0789_/a_315_47# _0298_ _0789_/a_208_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.12513 ps=1.035 w=0.65 l=0.15
X2005 VGND _0297_ _0789_/a_75_199# VGND sky130_fd_pr__nfet_01v8 ad=0.13487 pd=1.065 as=0.10563 ps=0.975 w=0.65 l=0.15
X2006 _0789_/a_75_199# _0299_ _0789_/a_315_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X2007 _0789_/a_75_199# _0277_ _0789_/a_544_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=1.415 w=1 l=0.15
X2008 _0789_/a_544_297# _0297_ _0789_/a_201_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.415 as=0.1625 ps=1.325 w=1 l=0.15
X2009 VPWR _0789_/a_75_199# _0405_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.285 ps=2.57 w=1 l=0.15
X2010 _0789_/a_201_297# _0404_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1425 ps=1.285 w=1 l=0.15
X2011 VPWR _0298_ _0789_/a_201_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X2012 _0789_/a_201_297# _0299_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.305 ps=1.61 w=1 l=0.15
X2013 VGND _0789_/a_75_199# _0405_ VGND sky130_fd_pr__nfet_01v8 ad=0.11213 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
X2014 VPWR clknet_1_1__leaf__0457_ _0858_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2015 _0458_ _0858_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2016 _0458_ _0858_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2017 VGND clknet_1_1__leaf__0457_ _0858_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2018 VPWR acc0.A\[31\] hold15/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2019 VGND hold15/a_285_47# hold15/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2020 net162 hold15/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2021 VGND acc0.A\[31\] hold15/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2022 VPWR hold15/a_285_47# hold15/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2023 hold15/a_285_47# hold15/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2024 hold15/a_285_47# hold15/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2025 net162 hold15/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2026 VPWR comp0.B\[9\] hold26/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2027 VGND hold26/a_285_47# hold26/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2028 net173 hold26/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2029 VGND comp0.B\[9\] hold26/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2030 VPWR hold26/a_285_47# hold26/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2031 hold26/a_285_47# hold26/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2032 hold26/a_285_47# hold26/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2033 net173 hold26/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2034 VPWR _0143_ hold37/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2035 VGND hold37/a_285_47# hold37/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2036 net184 hold37/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2037 VGND _0143_ hold37/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2038 VPWR hold37/a_285_47# hold37/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2039 hold37/a_285_47# hold37/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2040 hold37/a_285_47# hold37/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2041 net184 hold37/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2042 VPWR comp0.B\[12\] hold48/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2043 VGND hold48/a_285_47# hold48/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2044 net195 hold48/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2045 VGND comp0.B\[12\] hold48/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2046 VPWR hold48/a_285_47# hold48/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2047 hold48/a_285_47# hold48/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2048 hold48/a_285_47# hold48/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2049 net195 hold48/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2050 VPWR acc0.A\[18\] hold59/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2051 VGND hold59/a_285_47# hold59/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2052 net206 hold59/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2053 VGND acc0.A\[18\] hold59/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2054 VPWR hold59/a_285_47# hold59/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2055 hold59/a_285_47# hold59/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2056 hold59/a_285_47# hold59/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2057 net206 hold59/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2058 net73 clknet_1_1__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2059 VGND clknet_1_1__leaf__0458_ net73 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2060 net73 clknet_1_1__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2061 VPWR clknet_1_1__leaf__0458_ net73 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2062 _0643_/a_103_199# _0274_ _0643_/a_253_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2063 VPWR _0643_/a_103_199# _0275_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2064 _0643_/a_337_297# _0269_ _0643_/a_253_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2065 _0643_/a_103_199# _0272_ _0643_/a_337_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X2066 _0643_/a_253_297# _0260_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X2067 VPWR _0274_ _0643_/a_103_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X2068 VGND _0643_/a_103_199# _0275_ VGND sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X2069 _0643_/a_253_47# _0260_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X2070 _0643_/a_253_47# _0272_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2071 VGND _0269_ _0643_/a_253_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2072 _0712_/a_465_47# _0339_ _0712_/a_381_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1755 ps=1.84 w=0.65 l=0.15
X2073 VGND _0341_ _0712_/a_561_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X2074 VPWR _0340_ _0712_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.86 ps=7.72 w=1 l=0.15
X2075 _0712_/a_297_297# _0339_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2076 _0712_/a_297_297# _0341_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2077 VPWR _0220_ _0712_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2078 _0712_/a_381_47# _0220_ _0712_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.36725 ps=2.43 w=0.65 l=0.15
X2079 _0712_/a_297_297# _0343_ _0712_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2080 VPWR _0712_/a_79_21# _0344_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2081 _0712_/a_79_21# _0343_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2082 VGND _0712_/a_79_21# _0344_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2083 _0712_/a_561_47# _0340_ _0712_/a_465_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2084 VPWR _0216_ _0574_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2085 _0574_/a_27_297# _0217_ _0574_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2086 VGND _0216_ _0574_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2087 _0123_ _0574_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2088 _0574_/a_27_297# _0217_ _0574_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2089 _0574_/a_109_297# acc0.A\[25\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2090 _0574_/a_373_47# acc0.A\[25\] _0574_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2091 _0123_ _0574_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2092 _0574_/a_109_297# net199 _0574_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2093 _0574_/a_109_47# net199 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2094 acc0.A\[11\] _1057_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2095 _1057_/a_891_413# _1057_/a_193_47# _1057_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2096 _1057_/a_561_413# _1057_/a_27_47# _1057_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2097 VPWR net143 _1057_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2098 acc0.A\[11\] _1057_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2099 _1057_/a_381_47# net189 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2100 VGND _1057_/a_634_159# _1057_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2101 VPWR _1057_/a_891_413# _1057_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2102 _1057_/a_466_413# _1057_/a_193_47# _1057_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2103 VPWR _1057_/a_634_159# _1057_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2104 _1057_/a_634_159# _1057_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2105 _1057_/a_634_159# _1057_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2106 _1057_/a_975_413# _1057_/a_193_47# _1057_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2107 VGND _1057_/a_1059_315# _1057_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2108 _1057_/a_193_47# _1057_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2109 _1057_/a_891_413# _1057_/a_27_47# _1057_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2110 _1057_/a_592_47# _1057_/a_193_47# _1057_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2111 VPWR _1057_/a_1059_315# _1057_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2112 _1057_/a_1017_47# _1057_/a_27_47# _1057_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2113 _1057_/a_193_47# _1057_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2114 _1057_/a_466_413# _1057_/a_27_47# _1057_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2115 VGND _1057_/a_891_413# _1057_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2116 _1057_/a_381_47# net189 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2117 VGND net143 _1057_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2118 VPWR output49/a_27_47# pp[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2119 pp[21] output49/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2120 VPWR net49 output49/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2121 pp[21] output49/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X2122 VGND output49/a_27_47# pp[21] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2123 VGND net49 output49/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2124 VPWR output38/a_27_47# pp[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2125 pp[11] output38/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2126 VPWR net38 output38/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2127 pp[11] output38/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X2128 VGND output38/a_27_47# pp[11] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2129 VGND net38 output38/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2132 VPWR clk clkbuf_0_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X2133 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X2134 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2135 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2136 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2137 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2138 clkbuf_0_clk/a_110_47# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2139 clkbuf_0_clk/a_110_47# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X2140 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X2141 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2142 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2143 clkbuf_0_clk/a_110_47# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2144 VGND clk clkbuf_0_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2145 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2146 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2147 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2148 VGND clk clkbuf_0_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2149 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2150 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2151 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2152 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2153 clkbuf_0_clk/a_110_47# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2154 VPWR clk clkbuf_0_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2155 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2156 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2157 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2158 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2159 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2160 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2161 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2162 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2163 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2164 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2165 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2166 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2167 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2168 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2169 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2170 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2171 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2172 _0557_/a_240_47# net27 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X2173 _0134_ _0557_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2174 VGND _0208_ _0557_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2175 _0557_/a_51_297# net160 _0557_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X2176 _0557_/a_149_47# _0211_ _0557_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X2177 _0557_/a_240_47# _0173_ _0557_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2178 VPWR _0208_ _0557_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2179 _0134_ _0557_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X2180 _0557_/a_149_47# net160 _0557_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2181 _0557_/a_245_297# _0173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2182 VPWR _0211_ _0557_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2183 _0557_/a_512_297# net27 _0557_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2186 VGND _0256_ _0626_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2187 _0626_/a_68_297# _0257_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2188 _0258_ _0626_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2189 VPWR _0256_ _0626_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2190 _0258_ _0626_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2191 _0626_/a_150_297# _0257_ _0626_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2202 VPWR net63 hold101/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2203 VGND hold101/a_285_47# hold101/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2204 net248 hold101/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2205 VGND net63 hold101/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2206 VPWR hold101/a_285_47# hold101/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2207 hold101/a_285_47# hold101/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2208 hold101/a_285_47# hold101/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2209 net248 hold101/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2212 VPWR acc0.A\[19\] _0609_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2213 VGND acc0.A\[19\] _0241_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2214 _0609_/a_109_297# net46 _0241_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2215 _0241_ net46 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2216 VPWR control0.count\[1\] _0960_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2415 ps=2.83 w=0.42 l=0.15
X2217 VPWR control0.count\[2\] _0960_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2218 _0960_/a_181_47# control0.count\[0\] _0960_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0882 pd=1.26 as=0.0882 ps=1.26 w=0.42 l=0.15
X2219 VGND control0.count\[2\] _0960_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2220 _0960_/a_27_47# control0.count\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2221 _0478_ _0960_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2222 _0478_ _0960_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2223 _0960_/a_109_47# control0.count\[1\] _0960_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2224 VPWR clknet_1_0__leaf__0457_ _0891_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X2225 _0461_ _0891_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X2226 _0461_ _0891_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X2227 VGND clknet_1_0__leaf__0457_ _0891_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X2228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2230 clkload4/Y clknet_1_0__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.25
X2231 VGND clknet_1_0__leaf__0459_ clkload4/a_268_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1155 ps=1.52 w=0.55 l=0.15
X2232 clkload4/Y clknet_1_0__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X2233 clkload4/Y clknet_1_0__leaf__0459_ clkload4/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.154 pd=1.66 as=0.1155 ps=1.52 w=0.55 l=0.15
X2234 VPWR clknet_1_0__leaf__0459_ clkload4/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X2235 clkload4/a_110_47# clknet_1_0__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.15
X2236 clkload4/a_268_47# clknet_1_0__leaf__0459_ clkload4/Y VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.15
X2237 VPWR clknet_1_0__leaf__0459_ clkload4/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X2238 VPWR acc0.A\[22\] _0222_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2239 _0222_ acc0.A\[22\] _0590_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X2240 _0590_/a_113_47# net50 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2241 _0222_ net50 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2244 VPWR clknet_1_1__leaf_clk _0857_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X2245 _0457_ _0857_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X2246 _0457_ _0857_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X2247 VGND clknet_1_1__leaf_clk _0857_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X2248 VGND _0279_ _0788_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2249 _0788_/a_68_297# _0403_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2250 _0404_ _0788_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2251 VPWR _0279_ _0788_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2252 _0404_ _0788_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2253 _0788_/a_150_297# _0403_ _0788_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2254 VPWR _0129_ hold16/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2255 VGND hold16/a_285_47# hold16/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2256 net163 hold16/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2257 VGND _0129_ hold16/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2258 VPWR hold16/a_285_47# hold16/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2259 hold16/a_285_47# hold16/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2260 hold16/a_285_47# hold16/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2261 net163 hold16/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2262 VPWR _0138_ hold27/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2263 VGND hold27/a_285_47# hold27/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2264 net174 hold27/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2265 VGND _0138_ hold27/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2266 VPWR hold27/a_285_47# hold27/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2267 hold27/a_285_47# hold27/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2268 hold27/a_285_47# hold27/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2269 net174 hold27/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2270 VPWR comp0.B\[3\] hold38/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2271 VGND hold38/a_285_47# hold38/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2272 net185 hold38/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2273 VGND comp0.B\[3\] hold38/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2274 VPWR hold38/a_285_47# hold38/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2275 hold38/a_285_47# hold38/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2276 hold38/a_285_47# hold38/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2277 net185 hold38/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2278 VPWR _0141_ hold49/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2279 VGND hold49/a_285_47# hold49/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2280 net196 hold49/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2281 VGND _0141_ hold49/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2282 VPWR hold49/a_285_47# hold49/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2283 hold49/a_285_47# hold49/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2284 hold49/a_285_47# hold49/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2285 net196 hold49/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2290 _0343_ control0.add VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2291 VGND control0.add _0343_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2292 _0343_ control0.add VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2293 VPWR control0.add _0343_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2294 _0642_/a_298_297# _0642_/a_27_413# _0642_/a_215_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2295 _0642_/a_215_297# _0642_/a_27_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X2296 _0642_/a_298_297# _0273_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2297 _0274_ _0642_/a_215_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25837 ps=1.445 w=0.65 l=0.15
X2298 VPWR _0251_ _0642_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2299 _0274_ _0642_/a_215_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2300 _0642_/a_382_47# _0252_ _0642_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X2301 VGND _0251_ _0642_/a_27_413# VGND sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X2302 VPWR _0252_ _0642_/a_298_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X2303 VGND _0273_ _0642_/a_382_47# VGND sky130_fd_pr__nfet_01v8 ad=0.25837 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
X2304 VPWR _0178_ _0573_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X2305 VGND _0573_/a_27_47# _0217_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X2306 VGND _0573_/a_27_47# _0217_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2307 _0217_ _0573_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X2308 _0217_ _0573_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2309 VGND _0178_ _0573_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X2310 VPWR _0573_/a_27_47# _0217_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2311 _0217_ _0573_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2312 _0217_ _0573_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2313 VPWR _0573_/a_27_47# _0217_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2314 net108 clknet_1_0__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2315 VGND clknet_1_0__leaf__0462_ net108 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2316 net108 clknet_1_0__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2317 VPWR clknet_1_0__leaf__0462_ net108 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2318 acc0.A\[10\] _1056_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2319 _1056_/a_891_413# _1056_/a_193_47# _1056_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2320 _1056_/a_561_413# _1056_/a_27_47# _1056_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2321 VPWR net142 _1056_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2322 acc0.A\[10\] _1056_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2323 _1056_/a_381_47# net182 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2324 VGND _1056_/a_634_159# _1056_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2325 VPWR _1056_/a_891_413# _1056_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2326 _1056_/a_466_413# _1056_/a_193_47# _1056_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2327 VPWR _1056_/a_634_159# _1056_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2328 _1056_/a_634_159# _1056_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2329 _1056_/a_634_159# _1056_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2330 _1056_/a_975_413# _1056_/a_193_47# _1056_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2331 VGND _1056_/a_1059_315# _1056_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2332 _1056_/a_193_47# _1056_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2333 _1056_/a_891_413# _1056_/a_27_47# _1056_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2334 _1056_/a_592_47# _1056_/a_193_47# _1056_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2335 VPWR _1056_/a_1059_315# _1056_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2336 _1056_/a_1017_47# _1056_/a_27_47# _1056_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2337 _1056_/a_193_47# _1056_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2338 _1056_/a_466_413# _1056_/a_27_47# _1056_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2339 VGND _1056_/a_891_413# _1056_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2340 _1056_/a_381_47# net182 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2341 VGND net142 _1056_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2342 VPWR output39/a_27_47# pp[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2343 pp[12] output39/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2344 VPWR net39 output39/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2345 pp[12] output39/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X2346 VGND output39/a_27_47# pp[12] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2347 VGND net39 output39/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2348 net96 clknet_1_1__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2349 VGND clknet_1_1__leaf__0460_ net96 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2350 net96 clknet_1_1__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2351 VPWR clknet_1_1__leaf__0460_ net96 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2352 VPWR net63 _0625_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2353 _0257_ _0625_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X2354 VGND net63 _0625_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2355 _0625_/a_59_75# acc0.A\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2356 _0257_ _0625_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2357 _0625_/a_145_75# acc0.A\[5\] _0625_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X2358 VGND comp0.B\[4\] _0556_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2359 _0556_/a_68_297# _0175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2360 _0211_ _0556_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2361 VPWR comp0.B\[4\] _0556_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2362 _0211_ _0556_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2363 _0556_/a_150_297# _0175_ _0556_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2364 comp0.B\[7\] _1039_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2365 _1039_/a_891_413# _1039_/a_193_47# _1039_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2366 _1039_/a_561_413# _1039_/a_27_47# _1039_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2367 VPWR net125 _1039_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2368 comp0.B\[7\] _1039_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2369 _1039_/a_381_47# _0137_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2370 VGND _1039_/a_634_159# _1039_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2371 VPWR _1039_/a_891_413# _1039_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2372 _1039_/a_466_413# _1039_/a_193_47# _1039_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2373 VPWR _1039_/a_634_159# _1039_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2374 _1039_/a_634_159# _1039_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2375 _1039_/a_634_159# _1039_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2376 _1039_/a_975_413# _1039_/a_193_47# _1039_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2377 VGND _1039_/a_1059_315# _1039_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2378 _1039_/a_193_47# _1039_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2379 _1039_/a_891_413# _1039_/a_27_47# _1039_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2380 _1039_/a_592_47# _1039_/a_193_47# _1039_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2381 VPWR _1039_/a_1059_315# _1039_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2382 _1039_/a_1017_47# _1039_/a_27_47# _1039_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2383 _1039_/a_193_47# _1039_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2384 _1039_/a_466_413# _1039_/a_27_47# _1039_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2385 VGND _1039_/a_891_413# _1039_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2386 _1039_/a_381_47# _0137_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2387 VGND net125 _1039_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2392 _0240_ net44 _0608_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X2393 VPWR _0239_ _0240_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X2394 _0608_/a_27_47# net44 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X2395 _0240_ _0239_ _0608_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2396 _0608_/a_109_297# acc0.A\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2397 VGND acc0.A\[17\] _0608_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2398 VGND comp0.B\[12\] _0539_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2399 _0539_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2400 _0202_ _0539_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2401 VPWR comp0.B\[12\] _0539_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2402 _0202_ _0539_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2403 _0539_/a_150_297# _0176_ _0539_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2410 net147 clknet_1_0__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2411 VGND clknet_1_0__leaf__0465_ net147 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2412 net147 clknet_1_0__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2413 VPWR clknet_1_0__leaf__0465_ net147 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2418 control0.count\[3\] _1072_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2419 _1072_/a_891_413# _1072_/a_193_47# _1072_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2420 _1072_/a_561_413# _1072_/a_27_47# _1072_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2421 VPWR clknet_1_0__leaf_clk _1072_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2422 control0.count\[3\] _1072_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2423 _1072_/a_381_47# _0170_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2424 VGND _1072_/a_634_159# _1072_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2425 VPWR _1072_/a_891_413# _1072_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2426 _1072_/a_466_413# _1072_/a_193_47# _1072_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2427 VPWR _1072_/a_634_159# _1072_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2428 _1072_/a_634_159# _1072_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2429 _1072_/a_634_159# _1072_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2430 _1072_/a_975_413# _1072_/a_193_47# _1072_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2431 VGND _1072_/a_1059_315# _1072_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2432 _1072_/a_193_47# _1072_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2433 _1072_/a_891_413# _1072_/a_27_47# _1072_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2434 _1072_/a_592_47# _1072_/a_193_47# _1072_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2435 VPWR _1072_/a_1059_315# _1072_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2436 _1072_/a_1017_47# _1072_/a_27_47# _1072_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2437 _1072_/a_193_47# _1072_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2438 _1072_/a_466_413# _1072_/a_27_47# _1072_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2439 VGND _1072_/a_891_413# _1072_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2440 _1072_/a_381_47# _0170_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2441 VGND clknet_1_0__leaf_clk _1072_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2444 VPWR _0787_/a_80_21# _0403_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X2445 _0787_/a_209_297# _0402_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.65 pd=5.3 as=0 ps=0 w=1 l=0.15
X2446 _0787_/a_303_47# _0285_ _0787_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.208 ps=1.94 w=0.65 l=0.15
X2447 _0787_/a_209_47# _0402_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2448 VGND _0787_/a_80_21# _0403_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X2449 VGND _0284_ _0787_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X2450 _0787_/a_80_21# _0281_ _0787_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2451 VPWR _0285_ _0787_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2452 _0787_/a_80_21# _0284_ _0787_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0 ps=0 w=1 l=0.15
X2453 _0787_/a_209_297# _0281_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2454 VGND _0346_ _0856_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X2455 _0856_/a_510_47# _0456_ _0856_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X2456 _0856_/a_79_21# _0345_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X2457 VPWR _0456_ _0856_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2458 _0856_/a_79_21# _0264_ _0856_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X2459 _0856_/a_297_297# _0346_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2460 _0856_/a_79_21# _0345_ _0856_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X2461 VPWR _0856_/a_79_21# _0080_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2462 VGND _0856_/a_79_21# _0080_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2463 _0856_/a_215_47# _0264_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2464 VPWR control0.count\[2\] hold17/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2465 VGND hold17/a_285_47# hold17/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2466 net164 hold17/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2467 VGND control0.count\[2\] hold17/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2468 VPWR hold17/a_285_47# hold17/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2469 hold17/a_285_47# hold17/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2470 hold17/a_285_47# hold17/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2471 net164 hold17/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2472 VPWR acc0.A\[2\] hold28/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2473 VGND hold28/a_285_47# hold28/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2474 net175 hold28/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2475 VGND acc0.A\[2\] hold28/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2476 VPWR hold28/a_285_47# hold28/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2477 hold28/a_285_47# hold28/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2478 hold28/a_285_47# hold28/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2479 net175 hold28/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2480 VPWR _0132_ hold39/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2481 VGND hold39/a_285_47# hold39/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2482 net186 hold39/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2483 VGND _0132_ hold39/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2484 VPWR hold39/a_285_47# hold39/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2485 hold39/a_285_47# hold39/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2486 hold39/a_285_47# hold39/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2487 net186 hold39/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2490 _0342_ _0340_ _0710_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2491 _0342_ _0340_ _0710_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2492 VPWR _0339_ _0710_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X2493 _0710_/a_109_297# _0220_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2494 _0710_/a_381_47# _0220_ _0342_ VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X2495 _0710_/a_109_297# _0341_ _0342_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2496 _0710_/a_109_47# _0341_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2497 VGND _0339_ _0710_/a_381_47# VGND sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.06825 ps=0.86 w=0.65 l=0.15
X2498 VPWR acc0.A\[6\] _0273_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2499 _0273_ acc0.A\[6\] _0641_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X2500 _0641_/a_113_47# net64 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2501 _0273_ net64 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2502 VPWR _0216_ _0572_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2503 _0572_/a_27_297# _0195_ _0572_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2504 VGND _0216_ _0572_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2505 _0124_ _0572_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2506 _0572_/a_27_297# _0195_ _0572_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2507 _0572_/a_109_297# net155 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2508 _0572_/a_373_47# net155 _0572_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2509 _0124_ _0572_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2510 _0572_/a_109_297# net210 _0572_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2511 _0572_/a_109_47# net210 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2512 acc0.A\[9\] _1055_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2513 _1055_/a_891_413# _1055_/a_193_47# _1055_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2514 _1055_/a_561_413# _1055_/a_27_47# _1055_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2515 VPWR net141 _1055_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2516 acc0.A\[9\] _1055_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2517 _1055_/a_381_47# net179 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2518 VGND _1055_/a_634_159# _1055_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2519 VPWR _1055_/a_891_413# _1055_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2520 _1055_/a_466_413# _1055_/a_193_47# _1055_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2521 VPWR _1055_/a_634_159# _1055_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2522 _1055_/a_634_159# _1055_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2523 _1055_/a_634_159# _1055_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2524 _1055_/a_975_413# _1055_/a_193_47# _1055_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2525 VGND _1055_/a_1059_315# _1055_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2526 _1055_/a_193_47# _1055_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2527 _1055_/a_891_413# _1055_/a_27_47# _1055_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2528 _1055_/a_592_47# _1055_/a_193_47# _1055_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2529 VPWR _1055_/a_1059_315# _1055_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2530 _1055_/a_1017_47# _1055_/a_27_47# _1055_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2531 _1055_/a_193_47# _1055_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2532 _1055_/a_466_413# _1055_/a_27_47# _1055_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2533 VGND _1055_/a_891_413# _1055_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2534 _1055_/a_381_47# net179 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2535 VGND net141 _1055_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2536 VPWR _0432_ _0839_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2537 VGND _0432_ _0444_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2538 _0839_/a_109_297# _0443_ _0444_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2539 _0444_ _0443_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2542 VPWR net62 _0624_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2543 _0256_ _0624_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X2544 VGND net62 _0624_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2545 _0624_/a_59_75# acc0.A\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2546 _0256_ _0624_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2547 _0624_/a_145_75# acc0.A\[4\] _0624_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X2548 _0555_/a_240_47# net28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X2549 _0135_ _0555_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2550 VGND _0208_ _0555_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2551 _0555_/a_51_297# net204 _0555_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X2552 _0555_/a_149_47# _0210_ _0555_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X2553 _0555_/a_240_47# _0173_ _0555_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2554 VPWR _0208_ _0555_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2555 _0135_ _0555_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X2556 _0555_/a_149_47# net204 _0555_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2557 _0555_/a_245_297# _0173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2558 VPWR _0210_ _0555_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2559 _0555_/a_512_297# net28 _0555_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2562 comp0.B\[6\] _1038_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2563 _1038_/a_891_413# _1038_/a_193_47# _1038_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2564 _1038_/a_561_413# _1038_/a_27_47# _1038_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2565 VPWR net124 _1038_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2566 comp0.B\[6\] _1038_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2567 _1038_/a_381_47# net172 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2568 VGND _1038_/a_634_159# _1038_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2569 VPWR _1038_/a_891_413# _1038_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2570 _1038_/a_466_413# _1038_/a_193_47# _1038_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2571 VPWR _1038_/a_634_159# _1038_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2572 _1038_/a_634_159# _1038_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2573 _1038_/a_634_159# _1038_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2574 _1038_/a_975_413# _1038_/a_193_47# _1038_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2575 VGND _1038_/a_1059_315# _1038_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2576 _1038_/a_193_47# _1038_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2577 _1038_/a_891_413# _1038_/a_27_47# _1038_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2578 _1038_/a_592_47# _1038_/a_193_47# _1038_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2579 VPWR _1038_/a_1059_315# _1038_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2580 _1038_/a_1017_47# _1038_/a_27_47# _1038_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2581 _1038_/a_193_47# _1038_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2582 _1038_/a_466_413# _1038_/a_27_47# _1038_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2583 VGND _1038_/a_891_413# _1038_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2584 _1038_/a_381_47# net172 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2585 VGND net124 _1038_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2586 net100 clknet_1_0__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2587 VGND clknet_1_0__leaf__0461_ net100 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2588 net100 clknet_1_0__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2589 VPWR clknet_1_0__leaf__0461_ net100 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2590 _0538_/a_240_47# net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X2591 _0143_ _0538_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2592 VGND _0172_ _0538_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2593 _0538_/a_51_297# net183 _0538_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X2594 _0538_/a_149_47# _0201_ _0538_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X2595 _0538_/a_240_47# _0174_ _0538_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2596 VPWR _0172_ _0538_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2597 _0143_ _0538_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X2598 _0538_/a_149_47# net183 _0538_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2599 _0538_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2600 VPWR _0201_ _0538_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2601 _0538_/a_512_297# net21 _0538_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2602 VPWR net44 _0607_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2603 _0607_/a_27_297# net43 _0607_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2604 VGND net44 _0607_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2605 _0239_ _0607_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2606 _0607_/a_27_297# net43 _0607_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2607 _0607_/a_109_297# acc0.A\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2608 _0607_/a_373_47# acc0.A\[17\] _0607_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2609 _0239_ _0607_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2610 _0607_/a_109_297# acc0.A\[16\] _0607_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2611 _0607_/a_109_47# acc0.A\[16\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2612 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2616 net81 clknet_1_1__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2617 VGND clknet_1_1__leaf__0459_ net81 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2618 net81 clknet_1_1__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2619 VPWR clknet_1_1__leaf__0459_ net81 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2620 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2621 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2624 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2627 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2628 control0.count\[2\] _1071_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2629 _1071_/a_891_413# _1071_/a_193_47# _1071_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2630 _1071_/a_561_413# _1071_/a_27_47# _1071_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2631 VPWR clknet_1_0__leaf_clk _1071_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2632 control0.count\[2\] _1071_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2633 _1071_/a_381_47# _0169_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2634 VGND _1071_/a_634_159# _1071_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2635 VPWR _1071_/a_891_413# _1071_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2636 _1071_/a_466_413# _1071_/a_193_47# _1071_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2637 VPWR _1071_/a_634_159# _1071_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2638 _1071_/a_634_159# _1071_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2639 _1071_/a_634_159# _1071_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2640 _1071_/a_975_413# _1071_/a_193_47# _1071_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2641 VGND _1071_/a_1059_315# _1071_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2642 _1071_/a_193_47# _1071_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2643 _1071_/a_891_413# _1071_/a_27_47# _1071_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2644 _1071_/a_592_47# _1071_/a_193_47# _1071_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2645 VPWR _1071_/a_1059_315# _1071_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2646 _1071_/a_1017_47# _1071_/a_27_47# _1071_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2647 _1071_/a_193_47# _1071_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2648 _1071_/a_466_413# _1071_/a_27_47# _1071_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2649 VGND _1071_/a_891_413# _1071_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2650 _1071_/a_381_47# _0169_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2651 VGND clknet_1_0__leaf_clk _1071_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2652 VPWR clknet_1_1__leaf__0457_ _0924_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X2653 _0464_ _0924_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X2654 _0464_ _0924_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X2655 VGND clknet_1_1__leaf__0457_ _0924_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X2656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2659 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2660 _0855_/a_81_21# net234 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2661 _0855_/a_299_297# net234 _0855_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X2662 VPWR _0855_/a_81_21# _0456_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2663 VPWR net149 _0855_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2664 VGND _0855_/a_81_21# _0456_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2665 VGND _0350_ _0855_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X2666 _0855_/a_299_297# _0350_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2667 _0855_/a_384_47# net149 _0855_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2668 VPWR _0786_/a_80_21# _0402_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X2669 _0786_/a_80_21# _0289_ _0786_/a_472_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.31 ps=2.62 w=1 l=0.15
X2670 VPWR _0401_ _0786_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.545 ps=5.09 w=1 l=0.15
X2671 VGND _0283_ _0786_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.35425 ps=3.69 w=0.65 l=0.15
X2672 VGND _0786_/a_80_21# _0402_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X2673 _0786_/a_300_47# _0401_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2674 _0786_/a_217_297# _0295_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2675 _0786_/a_80_21# _0295_ _0786_/a_300_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2676 _0786_/a_472_297# _0283_ _0786_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2677 _0786_/a_80_21# _0289_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2678 VPWR acc0.A\[15\] hold18/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2679 VGND hold18/a_285_47# hold18/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2680 net165 hold18/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2681 VGND acc0.A\[15\] hold18/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2682 VPWR hold18/a_285_47# hold18/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2683 hold18/a_285_47# hold18/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2684 hold18/a_285_47# hold18/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2685 net165 hold18/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2686 VPWR acc0.A\[22\] hold29/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2687 VGND hold29/a_285_47# hold29/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2688 net176 hold29/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2689 VGND acc0.A\[22\] hold29/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2690 VPWR hold29/a_285_47# hold29/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2691 hold29/a_285_47# hold29/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2692 hold29/a_285_47# hold29/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2693 net176 hold29/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2698 _0272_ _0640_/a_215_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2699 _0640_/a_109_53# _0271_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2700 _0640_/a_215_297# _0640_/a_109_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2701 _0272_ _0640_/a_215_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10187 ps=0.99 w=0.65 l=0.15
X2702 _0640_/a_392_297# _0255_ _0640_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X2703 _0640_/a_465_297# _0257_ _0640_/a_392_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X2704 _0640_/a_215_297# _0257_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2705 VPWR _0254_ _0640_/a_465_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X2706 _0640_/a_297_297# _0640_/a_109_53# _0640_/a_215_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X2707 _0640_/a_109_53# _0271_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2708 VGND _0255_ _0640_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X2709 VGND _0254_ _0640_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X2710 VPWR _0216_ _0571_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2711 _0571_/a_27_297# _0195_ _0571_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2712 VGND _0216_ _0571_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2713 _0125_ _0571_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2714 _0571_/a_27_297# _0195_ _0571_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2715 _0571_/a_109_297# acc0.A\[27\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2716 _0571_/a_373_47# acc0.A\[27\] _0571_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2717 _0125_ _0571_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2718 _0571_/a_109_297# net155 _0571_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2719 _0571_/a_109_47# net155 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2720 acc0.A\[8\] _1054_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2721 _1054_/a_891_413# _1054_/a_193_47# _1054_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2722 _1054_/a_561_413# _1054_/a_27_47# _1054_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2723 VPWR net140 _1054_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2724 acc0.A\[8\] _1054_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2725 _1054_/a_381_47# net169 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2726 VGND _1054_/a_634_159# _1054_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2727 VPWR _1054_/a_891_413# _1054_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2728 _1054_/a_466_413# _1054_/a_193_47# _1054_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2729 VPWR _1054_/a_634_159# _1054_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2730 _1054_/a_634_159# _1054_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2731 _1054_/a_634_159# _1054_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2732 _1054_/a_975_413# _1054_/a_193_47# _1054_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2733 VGND _1054_/a_1059_315# _1054_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2734 _1054_/a_193_47# _1054_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2735 _1054_/a_891_413# _1054_/a_27_47# _1054_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2736 _1054_/a_592_47# _1054_/a_193_47# _1054_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2737 VPWR _1054_/a_1059_315# _1054_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2738 _1054_/a_1017_47# _1054_/a_27_47# _1054_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2739 _1054_/a_193_47# _1054_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2740 _1054_/a_466_413# _1054_/a_27_47# _1054_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2741 VGND _1054_/a_891_413# _1054_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2742 _1054_/a_381_47# net169 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2743 VGND net140 _1054_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2744 _0769_/a_81_21# _0244_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2745 _0769_/a_299_297# _0244_ _0769_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X2746 VPWR _0769_/a_81_21# _0389_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2747 VPWR _0386_ _0769_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2748 VGND _0769_/a_81_21# _0389_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2749 VGND _0388_ _0769_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X2750 _0769_/a_299_297# _0388_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2751 _0769_/a_384_47# _0386_ _0769_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2752 VPWR _0431_ _0838_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2753 VGND _0431_ _0443_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2754 _0838_/a_109_297# _0271_ _0443_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2755 _0443_ _0271_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2756 VPWR acc0.A\[5\] _0623_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2757 VGND acc0.A\[5\] _0255_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2758 _0623_/a_109_297# net63 _0255_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2759 _0255_ net63 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2760 VGND net160 _0554_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2761 _0554_/a_68_297# _0175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2762 _0210_ _0554_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2763 VPWR net160 _0554_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2764 _0210_ _0554_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2765 _0554_/a_150_297# _0175_ _0554_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2768 comp0.B\[5\] _1037_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2769 _1037_/a_891_413# _1037_/a_193_47# _1037_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2770 _1037_/a_561_413# _1037_/a_27_47# _1037_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2771 VPWR net123 _1037_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2772 comp0.B\[5\] _1037_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2773 _1037_/a_381_47# _0135_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2774 VGND _1037_/a_634_159# _1037_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2775 VPWR _1037_/a_891_413# _1037_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2776 _1037_/a_466_413# _1037_/a_193_47# _1037_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2777 VPWR _1037_/a_634_159# _1037_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2778 _1037_/a_634_159# _1037_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2779 _1037_/a_634_159# _1037_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2780 _1037_/a_975_413# _1037_/a_193_47# _1037_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2781 VGND _1037_/a_1059_315# _1037_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2782 _1037_/a_193_47# _1037_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2783 _1037_/a_891_413# _1037_/a_27_47# _1037_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2784 _1037_/a_592_47# _1037_/a_193_47# _1037_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2785 VPWR _1037_/a_1059_315# _1037_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2786 _1037_/a_1017_47# _1037_/a_27_47# _1037_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2787 _1037_/a_193_47# _1037_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2788 _1037_/a_466_413# _1037_/a_27_47# _1037_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2789 VGND _1037_/a_891_413# _1037_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2790 _1037_/a_381_47# _0135_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2791 VGND net123 _1037_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2792 net87 clknet_1_0__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2793 VGND clknet_1_0__leaf__0459_ net87 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2794 net87 clknet_1_0__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2795 VPWR clknet_1_0__leaf__0459_ net87 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2798 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2799 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2802 _0238_ _0606_/a_215_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0 ps=0 w=1 l=0.15
X2803 _0606_/a_109_53# _0237_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2804 _0606_/a_215_297# _0606_/a_109_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2415 pd=2.83 as=0 ps=0 w=0.42 l=0.15
X2805 _0238_ _0606_/a_215_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2806 _0606_/a_392_297# _0236_ _0606_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0903 pd=1.27 as=0.1365 ps=1.49 w=0.42 l=0.15
X2807 _0606_/a_465_297# _0234_ _0606_/a_392_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.45 as=0 ps=0 w=0.42 l=0.15
X2808 _0606_/a_215_297# _0234_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2809 VPWR _0225_ _0606_/a_465_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2810 _0606_/a_297_297# _0606_/a_109_53# _0606_/a_215_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2811 _0606_/a_109_53# _0237_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2812 VGND _0236_ _0606_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2813 VGND _0225_ _0606_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2814 VGND comp0.B\[13\] _0537_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2815 _0537_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2816 _0201_ _0537_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2817 VPWR comp0.B\[13\] _0537_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2818 _0201_ _0537_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2819 _0537_/a_150_297# _0176_ _0537_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2820 net76 clknet_1_1__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2821 VGND clknet_1_1__leaf__0458_ net76 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2822 net76 clknet_1_1__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2823 VPWR clknet_1_1__leaf__0458_ net76 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2824 net138 clknet_1_0__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2825 VGND clknet_1_0__leaf__0465_ net138 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2826 net138 clknet_1_0__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2827 VPWR clknet_1_0__leaf__0465_ net138 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2834 net119 clknet_1_1__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2835 VGND clknet_1_1__leaf__0463_ net119 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2836 net119 clknet_1_1__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2837 VPWR clknet_1_1__leaf__0463_ net119 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2838 control0.count\[1\] _1070_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2839 _1070_/a_891_413# _1070_/a_193_47# _1070_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2840 _1070_/a_561_413# _1070_/a_27_47# _1070_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2841 VPWR clknet_1_0__leaf_clk _1070_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2842 control0.count\[1\] _1070_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2843 _1070_/a_381_47# _0168_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2844 VGND _1070_/a_634_159# _1070_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2845 VPWR _1070_/a_891_413# _1070_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2846 _1070_/a_466_413# _1070_/a_193_47# _1070_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2847 VPWR _1070_/a_634_159# _1070_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2848 _1070_/a_634_159# _1070_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2849 _1070_/a_634_159# _1070_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2850 _1070_/a_975_413# _1070_/a_193_47# _1070_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2851 VGND _1070_/a_1059_315# _1070_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2852 _1070_/a_193_47# _1070_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2853 _1070_/a_891_413# _1070_/a_27_47# _1070_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2854 _1070_/a_592_47# _1070_/a_193_47# _1070_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2855 VPWR _1070_/a_1059_315# _1070_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2856 _1070_/a_1017_47# _1070_/a_27_47# _1070_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2857 _1070_/a_193_47# _1070_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2858 _1070_/a_466_413# _1070_/a_27_47# _1070_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2859 VGND _1070_/a_891_413# _1070_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2860 _1070_/a_381_47# _0168_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2861 VGND clknet_1_0__leaf_clk _1070_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2862 net133 clknet_1_0__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2863 VGND clknet_1_0__leaf__0464_ net133 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2864 net133 clknet_1_0__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2865 VPWR clknet_1_0__leaf__0464_ net133 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2866 VGND _0347_ _0854_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X2867 _0854_/a_510_47# _0455_ _0854_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X2868 _0854_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X2869 VPWR _0455_ _0854_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2870 _0854_/a_79_21# _0454_ _0854_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X2871 _0854_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2872 _0854_/a_79_21# _0399_ _0854_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X2873 VPWR _0854_/a_79_21# _0081_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2874 VGND _0854_/a_79_21# _0081_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2875 _0854_/a_215_47# _0454_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2876 _0785_/a_81_21# _0292_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2877 _0785_/a_299_297# _0292_ _0785_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X2878 VPWR _0785_/a_81_21# _0401_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2879 VPWR _0259_ _0785_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2880 VGND _0785_/a_81_21# _0401_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2881 VGND _0275_ _0785_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X2882 _0785_/a_299_297# _0275_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2883 _0785_/a_384_47# _0259_ _0785_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2884 VPWR _0114_ hold19/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2885 VGND hold19/a_285_47# hold19/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2886 net166 hold19/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2887 VGND _0114_ hold19/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2888 VPWR hold19/a_285_47# hold19/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2889 hold19/a_285_47# hold19/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2890 hold19/a_285_47# hold19/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2891 net166 hold19/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2892 VPWR _0216_ _0570_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2893 _0570_/a_27_297# _0195_ _0570_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2894 VGND _0216_ _0570_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2895 _0126_ _0570_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2896 _0570_/a_27_297# _0195_ _0570_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2897 _0570_/a_109_297# net190 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2898 _0570_/a_373_47# net190 _0570_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2899 _0126_ _0570_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2900 _0570_/a_109_297# net197 _0570_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2901 _0570_/a_109_47# net197 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2902 acc0.A\[7\] _1053_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2903 _1053_/a_891_413# _1053_/a_193_47# _1053_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2904 _1053_/a_561_413# _1053_/a_27_47# _1053_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2905 VPWR net139 _1053_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2906 acc0.A\[7\] _1053_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2907 _1053_/a_381_47# _0151_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2908 VGND _1053_/a_634_159# _1053_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2909 VPWR _1053_/a_891_413# _1053_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2910 _1053_/a_466_413# _1053_/a_193_47# _1053_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2911 VPWR _1053_/a_634_159# _1053_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2912 _1053_/a_634_159# _1053_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2913 _1053_/a_634_159# _1053_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2914 _1053_/a_975_413# _1053_/a_193_47# _1053_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2915 VGND _1053_/a_1059_315# _1053_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2916 _1053_/a_193_47# _1053_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2917 _1053_/a_891_413# _1053_/a_27_47# _1053_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2918 _1053_/a_592_47# _1053_/a_193_47# _1053_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2919 VPWR _1053_/a_1059_315# _1053_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2920 _1053_/a_1017_47# _1053_/a_27_47# _1053_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2921 _1053_/a_193_47# _1053_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2922 _1053_/a_466_413# _1053_/a_27_47# _1053_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2923 VGND _1053_/a_891_413# _1053_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2924 _1053_/a_381_47# _0151_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2925 VGND net139 _1053_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2926 _0837_/a_585_47# _0442_ _0837_/a_266_47# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.11863 ps=1.015 w=0.65 l=0.15
X2927 VGND _0440_ _0837_/a_266_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2928 VPWR _0837_/a_81_21# _0085_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.26 ps=2.52 w=1 l=0.15
X2929 _0837_/a_81_21# _0172_ _0837_/a_585_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2930 VGND _0837_/a_81_21# _0085_ VGND sky130_fd_pr__nfet_01v8 ad=0.20312 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
X2931 _0837_/a_266_297# _0346_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.3125 ps=1.625 w=1 l=0.15
X2932 _0837_/a_368_297# _0440_ _0837_/a_266_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X2933 _0837_/a_266_47# _0441_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.11863 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X2934 _0837_/a_266_47# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.20312 ps=1.275 w=0.65 l=0.15
X2935 _0837_/a_81_21# _0441_ _0837_/a_368_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X2936 _0837_/a_81_21# _0172_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X2937 VPWR _0442_ _0837_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X2938 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2939 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2940 _0388_ _0310_ _0768_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X2941 VPWR _0240_ _0388_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X2942 _0768_/a_27_47# _0310_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X2943 _0388_ _0240_ _0768_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2944 _0768_/a_109_297# _0387_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2945 VGND _0387_ _0768_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2946 VGND acc0.A\[28\] _0699_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2947 _0699_/a_68_297# net56 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2948 _0331_ _0699_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2949 VPWR acc0.A\[28\] _0699_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2950 _0331_ _0699_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2951 _0699_/a_150_297# net56 _0699_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2954 VPWR _0252_ _0254_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2955 _0254_ _0251_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2956 _0622_/a_193_47# _0252_ _0622_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2957 _0254_ _0251_ _0622_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2958 _0254_ _0253_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2959 _0622_/a_109_47# _0253_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2960 _0553_/a_240_47# net29 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X2961 _0136_ _0553_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2962 VGND _0208_ _0553_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2963 _0553_/a_51_297# net171 _0553_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X2964 _0553_/a_149_47# _0209_ _0553_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X2965 _0553_/a_240_47# _0174_ _0553_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2966 VPWR _0208_ _0553_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2967 _0136_ _0553_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X2968 _0553_/a_149_47# net171 _0553_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2969 _0553_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2970 VPWR _0209_ _0553_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2971 _0553_/a_512_297# net29 _0553_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2974 comp0.B\[4\] _1036_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2975 _1036_/a_891_413# _1036_/a_193_47# _1036_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2976 _1036_/a_561_413# _1036_/a_27_47# _1036_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2977 VPWR net122 _1036_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2978 comp0.B\[4\] _1036_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2979 _1036_/a_381_47# net161 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2980 VGND _1036_/a_634_159# _1036_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2981 VPWR _1036_/a_891_413# _1036_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2982 _1036_/a_466_413# _1036_/a_193_47# _1036_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2983 VPWR _1036_/a_634_159# _1036_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2984 _1036_/a_634_159# _1036_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2985 _1036_/a_634_159# _1036_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2986 _1036_/a_975_413# _1036_/a_193_47# _1036_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2987 VGND _1036_/a_1059_315# _1036_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2988 _1036_/a_193_47# _1036_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2989 _1036_/a_891_413# _1036_/a_27_47# _1036_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2990 _1036_/a_592_47# _1036_/a_193_47# _1036_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2991 VPWR _1036_/a_1059_315# _1036_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2992 _1036_/a_1017_47# _1036_/a_27_47# _1036_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2993 _1036_/a_193_47# _1036_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2994 _1036_/a_466_413# _1036_/a_27_47# _1036_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2995 VGND _1036_/a_891_413# _1036_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2996 _1036_/a_381_47# net161 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2997 VGND net122 _1036_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2999 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3002 _0536_/a_240_47# net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X3003 _0144_ _0536_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X3004 VGND _0172_ _0536_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3005 _0536_/a_51_297# net157 _0536_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X3006 _0536_/a_149_47# _0200_ _0536_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X3007 _0536_/a_240_47# _0174_ _0536_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3008 VPWR _0172_ _0536_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3009 _0144_ _0536_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X3010 _0536_/a_149_47# net157 _0536_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3011 _0536_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3012 VPWR _0200_ _0536_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3013 _0536_/a_512_297# net22 _0536_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3016 VPWR _0228_ _0605_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3017 VGND _0228_ _0237_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3018 _0605_/a_109_297# _0227_ _0237_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3019 _0237_ _0227_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3020 acc0.A\[19\] _1019_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3021 _1019_/a_891_413# _1019_/a_193_47# _1019_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3022 _1019_/a_561_413# _1019_/a_27_47# _1019_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3023 VPWR net105 _1019_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3024 acc0.A\[19\] _1019_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3025 _1019_/a_381_47# net207 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3026 VGND _1019_/a_634_159# _1019_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3027 VPWR _1019_/a_891_413# _1019_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3028 _1019_/a_466_413# _1019_/a_193_47# _1019_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3029 VPWR _1019_/a_634_159# _1019_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3030 _1019_/a_634_159# _1019_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3031 _1019_/a_634_159# _1019_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3032 _1019_/a_975_413# _1019_/a_193_47# _1019_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3033 VGND _1019_/a_1059_315# _1019_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3034 _1019_/a_193_47# _1019_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3035 _1019_/a_891_413# _1019_/a_27_47# _1019_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3036 _1019_/a_592_47# _1019_/a_193_47# _1019_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3037 VPWR _1019_/a_1059_315# _1019_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3038 _1019_/a_1017_47# _1019_/a_27_47# _1019_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3039 _1019_/a_193_47# _1019_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3040 _1019_/a_466_413# _1019_/a_27_47# _1019_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3041 VGND _1019_/a_891_413# _1019_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3042 _1019_/a_381_47# net207 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3043 VGND net105 _1019_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3044 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3045 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3048 VPWR clknet_0__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3049 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3050 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3051 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3052 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3053 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3054 clkbuf_1_1__f__0465_/a_110_47# clknet_0__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3055 clkbuf_1_1__f__0465_/a_110_47# clknet_0__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3056 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3057 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3058 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3059 clkbuf_1_1__f__0465_/a_110_47# clknet_0__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3060 VGND clknet_0__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3061 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3062 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3063 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3064 VGND clknet_0__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3065 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3066 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3067 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3068 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3069 clkbuf_1_1__f__0465_/a_110_47# clknet_0__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3070 VPWR clknet_0__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3071 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3072 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3073 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3074 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3075 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3076 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3077 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3078 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3079 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3080 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3081 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3082 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3083 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3084 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3085 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3086 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3087 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3088 _0519_/a_81_21# _0191_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X3089 _0519_/a_299_297# _0191_ _0519_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X3090 VPWR _0519_/a_81_21# _0152_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3091 VPWR net168 _0519_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3092 VGND _0519_/a_81_21# _0152_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3093 VGND _0179_ _0519_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X3094 _0519_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3095 _0519_/a_384_47# net168 _0519_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X3099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X3100 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3101 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3102 net44 _0999_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3103 _0999_/a_891_413# _0999_/a_193_47# _0999_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3104 _0999_/a_561_413# _0999_/a_27_47# _0999_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3105 VPWR net85 _0999_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3106 net44 _0999_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3107 _0999_/a_381_47# _0097_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3108 VGND _0999_/a_634_159# _0999_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3109 VPWR _0999_/a_891_413# _0999_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3110 _0999_/a_466_413# _0999_/a_193_47# _0999_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3111 VPWR _0999_/a_634_159# _0999_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3112 _0999_/a_634_159# _0999_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3113 _0999_/a_634_159# _0999_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3114 _0999_/a_975_413# _0999_/a_193_47# _0999_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3115 VGND _0999_/a_1059_315# _0999_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3116 _0999_/a_193_47# _0999_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3117 _0999_/a_891_413# _0999_/a_27_47# _0999_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3118 _0999_/a_592_47# _0999_/a_193_47# _0999_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3119 VPWR _0999_/a_1059_315# _0999_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3120 _0999_/a_1017_47# _0999_/a_27_47# _0999_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3121 _0999_/a_193_47# _0999_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3122 _0999_/a_466_413# _0999_/a_27_47# _0999_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3123 VGND _0999_/a_891_413# _0999_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3124 _0999_/a_381_47# _0097_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3125 VGND net85 _0999_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3126 VGND _0218_ _0853_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3127 _0853_/a_68_297# net47 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3128 _0455_ _0853_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3129 VPWR _0218_ _0853_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3130 _0455_ _0853_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3131 _0853_/a_150_297# net47 _0853_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3132 VPWR acc0.A\[14\] _0400_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3133 _0400_ acc0.A\[14\] _0784_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X3134 _0784_/a_113_47# net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3135 _0400_ net41 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3136 VPWR A[0] input1/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X3137 net1 input1/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X3138 net1 input1/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X3139 VGND A[0] input1/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X3140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X3145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X3146 acc0.A\[6\] _1052_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3147 _1052_/a_891_413# _1052_/a_193_47# _1052_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3148 _1052_/a_561_413# _1052_/a_27_47# _1052_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3149 VPWR net138 _1052_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3150 acc0.A\[6\] _1052_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3151 _1052_/a_381_47# _0150_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3152 VGND _1052_/a_634_159# _1052_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3153 VPWR _1052_/a_891_413# _1052_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3154 _1052_/a_466_413# _1052_/a_193_47# _1052_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3155 VPWR _1052_/a_634_159# _1052_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3156 _1052_/a_634_159# _1052_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3157 _1052_/a_634_159# _1052_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3158 _1052_/a_975_413# _1052_/a_193_47# _1052_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3159 VGND _1052_/a_1059_315# _1052_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3160 _1052_/a_193_47# _1052_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3161 _1052_/a_891_413# _1052_/a_27_47# _1052_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3162 _1052_/a_592_47# _1052_/a_193_47# _1052_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3163 VPWR _1052_/a_1059_315# _1052_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3164 _1052_/a_1017_47# _1052_/a_27_47# _1052_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3165 _1052_/a_193_47# _1052_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3166 _1052_/a_466_413# _1052_/a_27_47# _1052_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3167 VGND _1052_/a_891_413# _1052_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3168 _1052_/a_381_47# _0150_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3169 VGND net138 _1052_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3170 VGND _0218_ _0836_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3171 _0836_/a_68_297# net248 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3172 _0442_ _0836_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3173 VPWR _0218_ _0836_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3174 _0442_ _0836_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3175 _0836_/a_150_297# net248 _0836_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3176 VPWR _0305_ _0767_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3177 _0387_ _0767_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X3178 VGND _0305_ _0767_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3179 _0767_/a_59_75# _0294_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3180 _0387_ _0767_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X3181 _0767_/a_145_75# _0294_ _0767_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X3182 _0698_/a_199_47# _0317_ _0330_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X3183 _0698_/a_113_297# _0319_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X3184 _0330_ _0316_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3185 VPWR _0317_ _0698_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3186 _0698_/a_113_297# _0316_ _0330_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X3187 VGND _0319_ _0698_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3190 _0253_ _0621_/a_35_297# _0621_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X3191 _0253_ net64 _0621_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X3192 _0621_/a_35_297# net64 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X3193 _0621_/a_117_297# net64 _0621_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X3194 VPWR net64 _0621_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3195 VGND acc0.A\[6\] _0621_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3196 VGND _0621_/a_35_297# _0253_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3197 _0621_/a_285_297# acc0.A\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3198 VPWR acc0.A\[6\] _0621_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3199 _0621_/a_285_47# acc0.A\[6\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3200 VGND comp0.B\[6\] _0552_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3201 _0552_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3202 _0209_ _0552_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3203 VPWR comp0.B\[6\] _0552_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3204 _0209_ _0552_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3205 _0552_/a_150_297# _0176_ _0552_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3206 comp0.B\[3\] _1035_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3207 _1035_/a_891_413# _1035_/a_193_47# _1035_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3208 _1035_/a_561_413# _1035_/a_27_47# _1035_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3209 VPWR net121 _1035_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3210 comp0.B\[3\] _1035_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3211 _1035_/a_381_47# _0133_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3212 VGND _1035_/a_634_159# _1035_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3213 VPWR _1035_/a_891_413# _1035_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3214 _1035_/a_466_413# _1035_/a_193_47# _1035_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3215 VPWR _1035_/a_634_159# _1035_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3216 _1035_/a_634_159# _1035_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3217 _1035_/a_634_159# _1035_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3218 _1035_/a_975_413# _1035_/a_193_47# _1035_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3219 VGND _1035_/a_1059_315# _1035_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3220 _1035_/a_193_47# _1035_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3221 _1035_/a_891_413# _1035_/a_27_47# _1035_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3222 _1035_/a_592_47# _1035_/a_193_47# _1035_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3223 VPWR _1035_/a_1059_315# _1035_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3224 _1035_/a_1017_47# _1035_/a_27_47# _1035_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3225 _1035_/a_193_47# _1035_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3226 _1035_/a_466_413# _1035_/a_27_47# _1035_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3227 VGND _1035_/a_891_413# _1035_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3228 _1035_/a_381_47# _0133_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3229 VGND net121 _1035_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3232 _0819_/a_81_21# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X3233 _0819_/a_299_297# _0346_ _0819_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X3234 VPWR _0819_/a_81_21# _0428_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3235 VPWR _0401_ _0819_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3236 VGND _0819_/a_81_21# _0428_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3237 VGND _0427_ _0819_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X3238 _0819_/a_299_297# _0427_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3239 _0819_/a_384_47# _0401_ _0819_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3240 net92 clknet_1_0__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3241 VGND clknet_1_0__leaf__0460_ net92 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3242 net92 clknet_1_0__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3243 VPWR clknet_1_0__leaf__0460_ net92 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3244 VPWR _0226_ _0236_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3245 _0236_ _0226_ _0604_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X3246 _0604_/a_113_47# _0235_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3247 _0236_ _0235_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3249 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3250 VGND comp0.B\[14\] _0535_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3251 _0535_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3252 _0200_ _0535_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3253 VPWR comp0.B\[14\] _0535_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3254 _0200_ _0535_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3255 _0535_/a_150_297# _0176_ _0535_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3258 acc0.A\[18\] _1018_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3259 _1018_/a_891_413# _1018_/a_193_47# _1018_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3260 _1018_/a_561_413# _1018_/a_27_47# _1018_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3261 VPWR net104 _1018_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3262 acc0.A\[18\] _1018_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3263 _1018_/a_381_47# _0116_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3264 VGND _1018_/a_634_159# _1018_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3265 VPWR _1018_/a_891_413# _1018_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3266 _1018_/a_466_413# _1018_/a_193_47# _1018_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3267 VPWR _1018_/a_634_159# _1018_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3268 _1018_/a_634_159# _1018_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3269 _1018_/a_634_159# _1018_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3270 _1018_/a_975_413# _1018_/a_193_47# _1018_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3271 VGND _1018_/a_1059_315# _1018_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3272 _1018_/a_193_47# _1018_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3273 _1018_/a_891_413# _1018_/a_27_47# _1018_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3274 _1018_/a_592_47# _1018_/a_193_47# _1018_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3275 VPWR _1018_/a_1059_315# _1018_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3276 _1018_/a_1017_47# _1018_/a_27_47# _1018_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3277 _1018_/a_193_47# _1018_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3278 _1018_/a_466_413# _1018_/a_27_47# _1018_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3279 VGND _1018_/a_891_413# _1018_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3280 _1018_/a_381_47# _0116_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3281 VGND net104 _1018_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3282 VPWR clknet_0__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3283 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3284 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3285 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3286 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3287 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3288 clkbuf_1_1__f__0464_/a_110_47# clknet_0__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3289 clkbuf_1_1__f__0464_/a_110_47# clknet_0__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3290 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3291 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3292 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3293 clkbuf_1_1__f__0464_/a_110_47# clknet_0__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3294 VGND clknet_0__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3295 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3296 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3297 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3298 VGND clknet_0__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3299 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3300 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3301 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3302 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3303 clkbuf_1_1__f__0464_/a_110_47# clknet_0__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3304 VPWR clknet_0__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3305 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3306 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3307 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3308 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3309 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3310 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3311 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3312 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3313 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3314 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3315 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3316 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3317 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3318 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3319 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3320 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3321 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3322 VPWR net15 _0518_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X3323 _0518_/a_27_297# _0186_ _0518_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X3324 VGND net15 _0518_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X3325 _0191_ _0518_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3326 _0518_/a_27_297# _0186_ _0518_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X3327 _0518_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3328 _0518_/a_373_47# _0180_ _0518_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3329 _0191_ _0518_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3330 _0518_/a_109_297# acc0.A\[8\] _0518_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3331 _0518_/a_109_47# acc0.A\[8\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3334 net43 _0998_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3335 _0998_/a_891_413# _0998_/a_193_47# _0998_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3336 _0998_/a_561_413# _0998_/a_27_47# _0998_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3337 VPWR net84 _0998_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3338 net43 _0998_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3339 _0998_/a_381_47# _0096_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3340 VGND _0998_/a_634_159# _0998_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3341 VPWR _0998_/a_891_413# _0998_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3342 _0998_/a_466_413# _0998_/a_193_47# _0998_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3343 VPWR _0998_/a_634_159# _0998_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3344 _0998_/a_634_159# _0998_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3345 _0998_/a_634_159# _0998_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3346 _0998_/a_975_413# _0998_/a_193_47# _0998_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3347 VGND _0998_/a_1059_315# _0998_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3348 _0998_/a_193_47# _0998_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3349 _0998_/a_891_413# _0998_/a_27_47# _0998_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3350 _0998_/a_592_47# _0998_/a_193_47# _0998_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3351 VPWR _0998_/a_1059_315# _0998_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3352 _0998_/a_1017_47# _0998_/a_27_47# _0998_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3353 _0998_/a_193_47# _0998_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3354 _0998_/a_466_413# _0998_/a_27_47# _0998_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3355 VGND _0998_/a_891_413# _0998_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3356 _0998_/a_381_47# _0096_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3357 VGND net84 _0998_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3358 _0454_ _0852_/a_35_297# _0852_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X3359 _0454_ _0453_ _0852_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X3360 _0852_/a_35_297# _0453_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X3361 _0852_/a_117_297# _0453_ _0852_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X3362 VPWR _0453_ _0852_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3363 VGND _0264_ _0852_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3364 VGND _0852_/a_35_297# _0454_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3365 _0852_/a_285_297# _0264_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3366 VPWR _0264_ _0852_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3367 _0852_/a_285_47# _0264_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3368 VGND _0347_ _0783_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X3369 _0783_/a_510_47# _0398_ _0783_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X3370 _0783_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X3371 VPWR _0398_ _0783_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3372 _0783_/a_79_21# _0397_ _0783_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X3373 _0783_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3374 _0783_/a_79_21# _0399_ _0783_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X3375 VPWR _0783_/a_79_21# _0096_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3376 VGND _0783_/a_79_21# _0096_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3377 _0783_/a_215_47# _0397_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3378 VPWR input2/a_75_212# net2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3379 input2/a_75_212# A[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3380 input2/a_75_212# A[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3381 VGND input2/a_75_212# net2 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X3383 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X3384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X3385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X3386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3388 acc0.A\[5\] _1051_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3389 _1051_/a_891_413# _1051_/a_193_47# _1051_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3390 _1051_/a_561_413# _1051_/a_27_47# _1051_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3391 VPWR net137 _1051_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3392 acc0.A\[5\] _1051_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3393 _1051_/a_381_47# _0149_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3394 VGND _1051_/a_634_159# _1051_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3395 VPWR _1051_/a_891_413# _1051_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3396 _1051_/a_466_413# _1051_/a_193_47# _1051_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3397 VPWR _1051_/a_634_159# _1051_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3398 _1051_/a_634_159# _1051_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3399 _1051_/a_634_159# _1051_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3400 _1051_/a_975_413# _1051_/a_193_47# _1051_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3401 VGND _1051_/a_1059_315# _1051_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3402 _1051_/a_193_47# _1051_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3403 _1051_/a_891_413# _1051_/a_27_47# _1051_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3404 _1051_/a_592_47# _1051_/a_193_47# _1051_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3405 VPWR _1051_/a_1059_315# _1051_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3406 _1051_/a_1017_47# _1051_/a_27_47# _1051_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3407 _1051_/a_193_47# _1051_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3408 _1051_/a_466_413# _1051_/a_27_47# _1051_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3409 VGND _1051_/a_891_413# _1051_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3410 _1051_/a_381_47# _0149_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3411 VGND net137 _1051_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3412 _0835_/a_78_199# _0432_ _0835_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3413 VPWR _0257_ _0835_/a_493_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3414 _0835_/a_493_297# _0255_ _0835_/a_78_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3415 VPWR _0835_/a_78_199# _0441_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X3416 VGND _0255_ _0835_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X3417 _0835_/a_78_199# _0256_ _0835_/a_292_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X3418 _0835_/a_215_47# _0257_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3419 _0835_/a_215_47# _0256_ _0835_/a_78_199# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X3420 _0835_/a_292_297# _0432_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X3421 VGND _0835_/a_78_199# _0441_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3422 VPWR _0244_ _0766_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3423 VGND _0244_ _0386_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3424 _0766_/a_109_297# _0245_ _0386_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3425 _0386_ _0245_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3426 VPWR _0697_/a_80_21# _0329_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X3427 _0697_/a_80_21# _0322_ _0697_/a_472_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.31 ps=2.62 w=1 l=0.15
X3428 VPWR _0313_ _0697_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.545 ps=5.09 w=1 l=0.15
X3429 VGND _0328_ _0697_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.35425 ps=3.69 w=0.65 l=0.15
X3430 VGND _0697_/a_80_21# _0329_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X3431 _0697_/a_300_47# _0313_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X3432 _0697_/a_217_297# _0324_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3433 _0697_/a_80_21# _0324_ _0697_/a_300_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3434 _0697_/a_472_297# _0328_ _0697_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3435 _0697_/a_80_21# _0322_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3440 VPWR acc0.A\[7\] _0252_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3441 _0252_ acc0.A\[7\] _0620_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X3442 _0620_/a_113_47# net65 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3443 _0252_ net65 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3444 VPWR _0551_/a_27_47# _0208_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3445 _0208_ _0551_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3446 VPWR _0171_ _0551_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3447 _0208_ _0551_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X3448 VGND _0551_/a_27_47# _0208_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3449 VGND _0171_ _0551_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3450 comp0.B\[2\] _1034_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3451 _1034_/a_891_413# _1034_/a_193_47# _1034_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3452 _1034_/a_561_413# _1034_/a_27_47# _1034_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3453 VPWR net120 _1034_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3454 comp0.B\[2\] _1034_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3455 _1034_/a_381_47# net186 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3456 VGND _1034_/a_634_159# _1034_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3457 VPWR _1034_/a_891_413# _1034_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3458 _1034_/a_466_413# _1034_/a_193_47# _1034_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3459 VPWR _1034_/a_634_159# _1034_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3460 _1034_/a_634_159# _1034_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3461 _1034_/a_634_159# _1034_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3462 _1034_/a_975_413# _1034_/a_193_47# _1034_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3463 VGND _1034_/a_1059_315# _1034_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3464 _1034_/a_193_47# _1034_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3465 _1034_/a_891_413# _1034_/a_27_47# _1034_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3466 _1034_/a_592_47# _1034_/a_193_47# _1034_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3467 VPWR _1034_/a_1059_315# _1034_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3468 _1034_/a_1017_47# _1034_/a_27_47# _1034_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3469 _1034_/a_193_47# _1034_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3470 _1034_/a_466_413# _1034_/a_27_47# _1034_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3471 VGND _1034_/a_891_413# _1034_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3472 _1034_/a_381_47# net186 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3473 VGND net120 _1034_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3474 VPWR _0275_ _0427_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.53 ps=5.06 w=1 l=0.15
X3475 _0427_ _0259_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3476 _0818_/a_193_47# _0275_ _0818_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1755 ps=1.84 w=0.65 l=0.15
X3477 _0427_ _0259_ _0818_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3478 _0427_ _0292_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3479 _0818_/a_109_47# _0292_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3482 _0749_/a_81_21# _0236_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X3483 _0749_/a_299_297# _0236_ _0749_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X3484 VPWR _0749_/a_81_21# _0373_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3485 VPWR _0248_ _0749_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3486 VGND _0749_/a_81_21# _0373_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3487 VGND _0372_ _0749_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X3488 _0749_/a_299_297# _0372_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3489 _0749_/a_384_47# _0248_ _0749_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3494 _0534_/a_81_21# _0199_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X3495 _0534_/a_299_297# _0199_ _0534_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X3496 VPWR _0534_/a_81_21# _0145_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3497 VPWR net149 _0534_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3498 VGND _0534_/a_81_21# _0145_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3499 VGND _0195_ _0534_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X3500 _0534_/a_299_297# _0195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3501 _0534_/a_384_47# net149 _0534_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3502 VGND acc0.A\[20\] _0603_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3503 _0603_/a_68_297# net48 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3504 _0235_ _0603_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3505 VPWR acc0.A\[20\] _0603_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3506 _0235_ _0603_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3507 _0603_/a_150_297# net48 _0603_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3508 acc0.A\[17\] _1017_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3509 _1017_/a_891_413# _1017_/a_193_47# _1017_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3510 _1017_/a_561_413# _1017_/a_27_47# _1017_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3511 VPWR net103 _1017_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3512 acc0.A\[17\] _1017_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3513 _1017_/a_381_47# _0115_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3514 VGND _1017_/a_634_159# _1017_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3515 VPWR _1017_/a_891_413# _1017_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3516 _1017_/a_466_413# _1017_/a_193_47# _1017_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3517 VPWR _1017_/a_634_159# _1017_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3518 _1017_/a_634_159# _1017_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3519 _1017_/a_634_159# _1017_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3520 _1017_/a_975_413# _1017_/a_193_47# _1017_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3521 VGND _1017_/a_1059_315# _1017_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3522 _1017_/a_193_47# _1017_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3523 _1017_/a_891_413# _1017_/a_27_47# _1017_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3524 _1017_/a_592_47# _1017_/a_193_47# _1017_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3525 VPWR _1017_/a_1059_315# _1017_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3526 _1017_/a_1017_47# _1017_/a_27_47# _1017_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3527 _1017_/a_193_47# _1017_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3528 _1017_/a_466_413# _1017_/a_27_47# _1017_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3529 VGND _1017_/a_891_413# _1017_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3530 _1017_/a_381_47# _0115_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3531 VGND net103 _1017_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3532 VPWR clknet_0__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3533 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3534 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3535 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3536 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3537 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3538 clkbuf_1_1__f__0463_/a_110_47# clknet_0__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3539 clkbuf_1_1__f__0463_/a_110_47# clknet_0__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3540 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3541 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3542 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3543 clkbuf_1_1__f__0463_/a_110_47# clknet_0__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3544 VGND clknet_0__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3545 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3546 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3547 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3548 VGND clknet_0__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3549 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3550 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3551 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3552 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3553 clkbuf_1_1__f__0463_/a_110_47# clknet_0__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3554 VPWR clknet_0__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3555 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3556 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3557 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3558 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3559 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3560 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3561 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3562 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3563 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3564 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3565 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3566 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3567 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3568 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3569 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3570 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3571 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3576 _0517_/a_81_21# _0190_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X3577 _0517_/a_299_297# _0190_ _0517_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X3578 VPWR _0517_/a_81_21# _0153_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3579 VPWR net178 _0517_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3580 VGND _0517_/a_81_21# _0153_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3581 VGND _0179_ _0517_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X3582 _0517_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3583 _0517_/a_384_47# net178 _0517_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3584 net130 clknet_1_1__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3585 VGND clknet_1_1__leaf__0464_ net130 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3586 net130 clknet_1_1__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3587 VPWR clknet_1_1__leaf__0464_ net130 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3588 net144 clknet_1_1__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3589 VGND clknet_1_1__leaf__0465_ net144 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3590 net144 clknet_1_1__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3591 VPWR clknet_1_1__leaf__0465_ net144 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3592 net42 _0997_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3593 _0997_/a_891_413# _0997_/a_193_47# _0997_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3594 _0997_/a_561_413# _0997_/a_27_47# _0997_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3595 VPWR net83 _0997_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3596 net42 _0997_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3597 _0997_/a_381_47# _0095_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3598 VGND _0997_/a_634_159# _0997_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3599 VPWR _0997_/a_891_413# _0997_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3600 _0997_/a_466_413# _0997_/a_193_47# _0997_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3601 VPWR _0997_/a_634_159# _0997_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3602 _0997_/a_634_159# _0997_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3603 _0997_/a_634_159# _0997_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3604 _0997_/a_975_413# _0997_/a_193_47# _0997_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3605 VGND _0997_/a_1059_315# _0997_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3606 _0997_/a_193_47# _0997_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3607 _0997_/a_891_413# _0997_/a_27_47# _0997_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3608 _0997_/a_592_47# _0997_/a_193_47# _0997_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3609 VPWR _0997_/a_1059_315# _0997_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3610 _0997_/a_1017_47# _0997_/a_27_47# _0997_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3611 _0997_/a_193_47# _0997_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3612 _0997_/a_466_413# _0997_/a_27_47# _0997_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3613 VGND _0997_/a_891_413# _0997_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3614 _0997_/a_381_47# _0095_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3615 VGND net83 _0997_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3616 VPWR _0465_ clkbuf_0__0465_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3617 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3618 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3619 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3620 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3621 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3622 clkbuf_0__0465_/a_110_47# _0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3623 clkbuf_0__0465_/a_110_47# _0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3624 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3625 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3626 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3627 clkbuf_0__0465_/a_110_47# _0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3628 VGND _0465_ clkbuf_0__0465_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3629 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3630 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3631 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3632 VGND _0465_ clkbuf_0__0465_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3633 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3634 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3635 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3636 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3637 clkbuf_0__0465_/a_110_47# _0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3638 VPWR _0465_ clkbuf_0__0465_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3639 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3640 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3641 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3642 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3643 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3644 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3645 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3646 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3647 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3648 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3649 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3650 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3651 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3652 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3653 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3654 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3655 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3658 VPWR _0266_ _0453_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3659 _0453_ _0266_ _0851_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X3660 _0851_/a_113_47# _0452_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3661 _0453_ _0452_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3662 VPWR _0208_ _0782_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X3663 VGND _0782_/a_27_47# _0399_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X3664 VGND _0782_/a_27_47# _0399_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3665 _0399_ _0782_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X3666 _0399_ _0782_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3667 VGND _0208_ _0782_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X3668 VPWR _0782_/a_27_47# _0399_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3669 _0399_ _0782_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3670 _0399_ _0782_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3671 VPWR _0782_/a_27_47# _0399_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3672 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3673 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3674 net111 clknet_1_0__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3675 VGND clknet_1_0__leaf__0462_ net111 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3676 net111 clknet_1_0__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3677 VPWR clknet_1_0__leaf__0462_ net111 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3678 net125 clknet_1_0__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3679 VGND clknet_1_0__leaf__0463_ net125 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3680 net125 clknet_1_0__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3681 VPWR clknet_1_0__leaf__0463_ net125 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3682 VPWR input3/a_75_212# net3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X3683 input3/a_75_212# A[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X3684 input3/a_75_212# A[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X3685 VGND input3/a_75_212# net3 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X3686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3687 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3690 acc0.A\[4\] _1050_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3691 _1050_/a_891_413# _1050_/a_193_47# _1050_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3692 _1050_/a_561_413# _1050_/a_27_47# _1050_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3693 VPWR net136 _1050_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3694 acc0.A\[4\] _1050_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3695 _1050_/a_381_47# _0148_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3696 VGND _1050_/a_634_159# _1050_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3697 VPWR _1050_/a_891_413# _1050_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3698 _1050_/a_466_413# _1050_/a_193_47# _1050_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3699 VPWR _1050_/a_634_159# _1050_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3700 _1050_/a_634_159# _1050_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3701 _1050_/a_634_159# _1050_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3702 _1050_/a_975_413# _1050_/a_193_47# _1050_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3703 VGND _1050_/a_1059_315# _1050_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3704 _1050_/a_193_47# _1050_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3705 _1050_/a_891_413# _1050_/a_27_47# _1050_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3706 _1050_/a_592_47# _1050_/a_193_47# _1050_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3707 VPWR _1050_/a_1059_315# _1050_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3708 _1050_/a_1017_47# _1050_/a_27_47# _1050_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3709 _1050_/a_193_47# _1050_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3710 _1050_/a_466_413# _1050_/a_27_47# _1050_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3711 VGND _1050_/a_891_413# _1050_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3712 _1050_/a_381_47# _0148_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3713 VGND net136 _1050_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3714 VPWR _0255_ _0834_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3715 VGND _0255_ _0440_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3716 _0834_/a_109_297# _0433_ _0440_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3717 _0440_ _0433_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3718 VPWR acc0.A\[25\] _0696_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3719 VGND acc0.A\[25\] _0328_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3720 _0696_/a_109_297# net53 _0328_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3721 _0328_ net53 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3722 VGND _0369_ _0765_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X3723 _0765_/a_510_47# _0385_ _0765_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X3724 _0765_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X3725 VPWR _0385_ _0765_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3726 _0765_/a_79_21# net220 _0765_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X3727 _0765_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3728 _0765_/a_79_21# _0352_ _0765_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X3729 VPWR _0765_/a_79_21# _0100_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3730 VGND _0765_/a_79_21# _0100_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3731 _0765_/a_215_47# net220 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3732 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3734 net106 clknet_1_0__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3735 VGND clknet_1_0__leaf__0461_ net106 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3736 net106 clknet_1_0__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3737 VPWR clknet_1_0__leaf__0461_ net106 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3738 _0550_/a_240_47# net30 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X3739 _0137_ _0550_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X3740 VGND _0172_ _0550_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3741 _0550_/a_51_297# net180 _0550_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X3742 _0550_/a_149_47# _0207_ _0550_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X3743 _0550_/a_240_47# _0174_ _0550_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3744 VPWR _0172_ _0550_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3745 _0137_ _0550_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X3746 _0550_/a_149_47# net180 _0550_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3747 _0550_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3748 VPWR _0207_ _0550_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3749 _0550_/a_512_297# net30 _0550_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3750 comp0.B\[1\] _1033_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3751 _1033_/a_891_413# _1033_/a_193_47# _1033_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3752 _1033_/a_561_413# _1033_/a_27_47# _1033_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3753 VPWR net119 _1033_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3754 comp0.B\[1\] _1033_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3755 _1033_/a_381_47# _0131_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3756 VGND _1033_/a_634_159# _1033_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3757 VPWR _1033_/a_891_413# _1033_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3758 _1033_/a_466_413# _1033_/a_193_47# _1033_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3759 VPWR _1033_/a_634_159# _1033_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3760 _1033_/a_634_159# _1033_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3761 _1033_/a_634_159# _1033_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3762 _1033_/a_975_413# _1033_/a_193_47# _1033_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3763 VGND _1033_/a_1059_315# _1033_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3764 _1033_/a_193_47# _1033_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3765 _1033_/a_891_413# _1033_/a_27_47# _1033_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3766 _1033_/a_592_47# _1033_/a_193_47# _1033_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3767 VPWR _1033_/a_1059_315# _1033_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3768 _1033_/a_1017_47# _1033_/a_27_47# _1033_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3769 _1033_/a_193_47# _1033_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3770 _1033_/a_466_413# _1033_/a_27_47# _1033_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3771 VGND _1033_/a_891_413# _1033_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3772 _1033_/a_381_47# _0131_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3773 VGND net119 _1033_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3774 _0817_/a_585_47# _0426_ _0817_/a_266_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.47125 ps=4.05 w=0.65 l=0.15
X3775 VGND _0424_ _0817_/a_266_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3776 VPWR _0817_/a_81_21# _0089_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3777 _0817_/a_81_21# _0345_ _0817_/a_585_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3778 VGND _0817_/a_81_21# _0089_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3779 _0817_/a_266_297# _0346_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0 ps=0 w=1 l=0.15
X3780 _0817_/a_368_297# _0424_ _0817_/a_266_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0 ps=0 w=1 l=0.15
X3781 _0817_/a_266_47# _0425_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3782 _0817_/a_266_47# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3783 _0817_/a_81_21# _0425_ _0817_/a_368_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.535 pd=5.07 as=0 ps=0 w=1 l=0.15
X3784 _0817_/a_81_21# _0345_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3785 VPWR _0426_ _0817_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3786 _0748_/a_81_21# _0311_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X3787 _0748_/a_299_297# _0311_ _0748_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X3788 VPWR _0748_/a_81_21# _0372_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3789 VPWR _0294_ _0748_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3790 VGND _0748_/a_81_21# _0372_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3791 VGND _0305_ _0748_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X3792 _0748_/a_299_297# _0305_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3793 _0748_/a_384_47# _0294_ _0748_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3794 VGND _0246_ _0679_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3795 _0679_/a_68_297# _0310_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3796 _0311_ _0679_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3797 VPWR _0246_ _0679_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3798 _0311_ _0679_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3799 _0679_/a_150_297# _0310_ _0679_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3802 VPWR _0233_ _0234_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3803 _0234_ _0233_ _0602_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X3804 _0602_/a_113_47# _0231_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3805 _0234_ _0231_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3806 VPWR net8 _0533_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X3807 _0533_/a_27_297# _0182_ _0533_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X3808 VGND net8 _0533_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X3809 _0199_ _0533_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3810 _0533_/a_27_297# _0182_ _0533_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X3811 _0533_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3812 _0533_/a_373_47# _0180_ _0533_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3813 _0199_ _0533_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3814 _0533_/a_109_297# acc0.A\[1\] _0533_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3815 _0533_/a_109_47# acc0.A\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X3817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X3818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3820 acc0.A\[16\] _1016_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3821 _1016_/a_891_413# _1016_/a_193_47# _1016_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3822 _1016_/a_561_413# _1016_/a_27_47# _1016_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3823 VPWR net102 _1016_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3824 acc0.A\[16\] _1016_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3825 _1016_/a_381_47# net166 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3826 VGND _1016_/a_634_159# _1016_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3827 VPWR _1016_/a_891_413# _1016_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3828 _1016_/a_466_413# _1016_/a_193_47# _1016_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3829 VPWR _1016_/a_634_159# _1016_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3830 _1016_/a_634_159# _1016_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3831 _1016_/a_634_159# _1016_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3832 _1016_/a_975_413# _1016_/a_193_47# _1016_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3833 VGND _1016_/a_1059_315# _1016_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3834 _1016_/a_193_47# _1016_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3835 _1016_/a_891_413# _1016_/a_27_47# _1016_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3836 _1016_/a_592_47# _1016_/a_193_47# _1016_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3837 VPWR _1016_/a_1059_315# _1016_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3838 _1016_/a_1017_47# _1016_/a_27_47# _1016_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3839 _1016_/a_193_47# _1016_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3840 _1016_/a_466_413# _1016_/a_27_47# _1016_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3841 VGND _1016_/a_891_413# _1016_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3842 _1016_/a_381_47# net166 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3843 VGND net102 _1016_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3844 VPWR clknet_0__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3845 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3846 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3847 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3848 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3849 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3850 clkbuf_1_1__f__0462_/a_110_47# clknet_0__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3851 clkbuf_1_1__f__0462_/a_110_47# clknet_0__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3852 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3853 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3854 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3855 clkbuf_1_1__f__0462_/a_110_47# clknet_0__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3856 VGND clknet_0__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3857 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3858 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3859 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3860 VGND clknet_0__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3861 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3862 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3863 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3864 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3865 clkbuf_1_1__f__0462_/a_110_47# clknet_0__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3866 VPWR clknet_0__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3867 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3868 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3869 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3870 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3871 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3872 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3873 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3874 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3875 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3876 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3877 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3878 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3879 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3880 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3881 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3882 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3883 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3884 net97 clknet_1_1__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3885 VGND clknet_1_1__leaf__0460_ net97 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3886 net97 clknet_1_1__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3887 VPWR clknet_1_1__leaf__0460_ net97 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3888 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3889 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3890 VPWR net16 _0516_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X3891 _0516_/a_27_297# _0186_ _0516_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X3892 VGND net16 _0516_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X3893 _0190_ _0516_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3894 _0516_/a_27_297# _0186_ _0516_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X3895 _0516_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3896 _0516_/a_373_47# _0181_ _0516_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3897 _0190_ _0516_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3898 _0516_/a_109_297# acc0.A\[9\] _0516_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3899 _0516_/a_109_47# acc0.A\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3904 net41 _0996_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3905 _0996_/a_891_413# _0996_/a_193_47# _0996_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3906 _0996_/a_561_413# _0996_/a_27_47# _0996_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3907 VPWR net82 _0996_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3908 net41 _0996_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3909 _0996_/a_381_47# _0094_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3910 VGND _0996_/a_634_159# _0996_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3911 VPWR _0996_/a_891_413# _0996_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3912 _0996_/a_466_413# _0996_/a_193_47# _0996_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3913 VPWR _0996_/a_634_159# _0996_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3914 _0996_/a_634_159# _0996_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3915 _0996_/a_634_159# _0996_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3916 _0996_/a_975_413# _0996_/a_193_47# _0996_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3917 VGND _0996_/a_1059_315# _0996_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3918 _0996_/a_193_47# _0996_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3919 _0996_/a_891_413# _0996_/a_27_47# _0996_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3920 _0996_/a_592_47# _0996_/a_193_47# _0996_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3921 VPWR _0996_/a_1059_315# _0996_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3922 _0996_/a_1017_47# _0996_/a_27_47# _0996_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3923 _0996_/a_193_47# _0996_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3924 _0996_/a_466_413# _0996_/a_27_47# _0996_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3925 VGND _0996_/a_891_413# _0996_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3926 _0996_/a_381_47# _0094_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3927 VGND net82 _0996_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3928 VPWR _0464_ clkbuf_0__0464_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3929 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3930 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3931 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3932 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3933 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3934 clkbuf_0__0464_/a_110_47# _0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3935 clkbuf_0__0464_/a_110_47# _0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3936 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3937 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3938 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3939 clkbuf_0__0464_/a_110_47# _0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3940 VGND _0464_ clkbuf_0__0464_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3941 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3942 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3943 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3944 VGND _0464_ clkbuf_0__0464_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3945 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3946 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3947 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3948 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3949 clkbuf_0__0464_/a_110_47# _0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3950 VPWR _0464_ clkbuf_0__0464_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3951 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3952 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3953 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3954 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3955 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3956 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3957 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3958 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3959 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3960 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3961 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3962 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3963 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3964 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3965 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3966 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3967 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3976 VGND acc0.A\[1\] _0850_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3977 _0850_/a_68_297# net47 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3978 _0452_ _0850_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3979 VPWR acc0.A\[1\] _0850_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3980 _0452_ _0850_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3981 _0850_/a_150_297# net47 _0850_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3982 VGND _0218_ _0781_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3983 _0781_/a_68_297# net43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3984 _0398_ _0781_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3985 VPWR _0218_ _0781_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3986 _0398_ _0781_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3987 _0781_/a_150_297# net43 _0781_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3988 VPWR input4/a_75_212# net4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X3989 input4/a_75_212# A[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X3990 input4/a_75_212# A[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X3991 VGND input4/a_75_212# net4 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X3992 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3993 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3996 VPWR _0466_ _0979_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X3997 _0979_/a_27_297# _0480_ _0979_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X3998 VGND _0466_ _0979_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X3999 _0169_ _0979_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4000 _0979_/a_27_297# _0480_ _0979_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X4001 _0979_/a_109_297# net164 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4002 _0979_/a_373_47# net164 _0979_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4003 _0169_ _0979_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4004 _0979_/a_109_297# _0488_ _0979_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4005 _0979_/a_109_47# _0488_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4006 VPWR clknet_1_0__leaf__0457_ _0902_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4007 _0462_ _0902_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4008 _0462_ _0902_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4009 VGND clknet_1_0__leaf__0457_ _0902_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4010 VGND _0369_ _0833_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X4011 _0833_/a_510_47# _0439_ _0833_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X4012 _0833_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X4013 VPWR _0439_ _0833_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4014 _0833_/a_79_21# net235 _0833_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X4015 _0833_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4016 _0833_/a_79_21# _0399_ _0833_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X4017 VPWR _0833_/a_79_21# _0086_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4018 VGND _0833_/a_79_21# _0086_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4019 _0833_/a_215_47# net235 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4020 _0764_/a_81_21# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4021 _0764_/a_299_297# _0346_ _0764_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4022 VPWR _0764_/a_81_21# _0385_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4023 VPWR _0373_ _0764_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4024 VGND _0764_/a_81_21# _0385_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4025 VGND _0384_ _0764_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4026 _0764_/a_299_297# _0384_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4027 _0764_/a_384_47# _0373_ _0764_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4028 VPWR _0695_/a_80_21# _0327_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X4029 _0695_/a_80_21# _0326_ _0695_/a_472_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.31 ps=2.62 w=1 l=0.15
X4030 VPWR _0312_ _0695_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.545 ps=5.09 w=1 l=0.15
X4031 VGND _0323_ _0695_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.35425 ps=3.69 w=0.65 l=0.15
X4032 VGND _0695_/a_80_21# _0327_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X4033 _0695_/a_300_47# _0312_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X4034 _0695_/a_217_297# _0250_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4035 _0695_/a_80_21# _0250_ _0695_/a_300_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4036 _0695_/a_472_297# _0323_ _0695_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4037 _0695_/a_80_21# _0326_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4038 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4039 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4040 net103 clknet_1_1__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4041 VGND clknet_1_1__leaf__0461_ net103 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4042 net103 clknet_1_1__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4043 VPWR clknet_1_1__leaf__0461_ net103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4044 comp0.B\[0\] _1032_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4045 _1032_/a_891_413# _1032_/a_193_47# _1032_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4046 _1032_/a_561_413# _1032_/a_27_47# _1032_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4047 VPWR net118 _1032_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4048 comp0.B\[0\] _1032_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4049 _1032_/a_381_47# net202 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4050 VGND _1032_/a_634_159# _1032_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4051 VPWR _1032_/a_891_413# _1032_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4052 _1032_/a_466_413# _1032_/a_193_47# _1032_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4053 VPWR _1032_/a_634_159# _1032_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4054 _1032_/a_634_159# _1032_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4055 _1032_/a_634_159# _1032_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4056 _1032_/a_975_413# _1032_/a_193_47# _1032_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4057 VGND _1032_/a_1059_315# _1032_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4058 _1032_/a_193_47# _1032_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4059 _1032_/a_891_413# _1032_/a_27_47# _1032_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4060 _1032_/a_592_47# _1032_/a_193_47# _1032_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4061 VPWR _1032_/a_1059_315# _1032_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4062 _1032_/a_1017_47# _1032_/a_27_47# _1032_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4063 _1032_/a_193_47# _1032_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4064 _1032_/a_466_413# _1032_/a_27_47# _1032_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4065 VGND _1032_/a_891_413# _1032_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4066 _1032_/a_381_47# net202 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4067 VGND net118 _1032_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4068 VGND _0218_ _0816_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4069 _0816_/a_68_297# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4070 _0426_ _0816_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4071 VPWR _0218_ _0816_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4072 _0426_ _0816_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4073 _0816_/a_150_297# net67 _0816_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4074 VGND _0369_ _0747_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X4075 _0747_/a_510_47# _0371_ _0747_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X4076 _0747_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X4077 VPWR _0371_ _0747_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4078 _0747_/a_79_21# net216 _0747_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X4079 _0747_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4080 _0747_/a_79_21# _0352_ _0747_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X4081 VPWR _0747_/a_79_21# _0104_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4082 VGND _0747_/a_79_21# _0104_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4083 _0747_/a_215_47# net216 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4084 VGND _0308_ _0678_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4085 _0678_/a_68_297# _0309_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4086 _0310_ _0678_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4087 VPWR _0308_ _0678_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4088 _0310_ _0678_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4089 _0678_/a_150_297# _0309_ _0678_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4090 VGND acc0.A\[23\] _0601_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4091 _0601_/a_68_297# net51 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4092 _0233_ _0601_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4093 VPWR acc0.A\[23\] _0601_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4094 _0233_ _0601_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4095 _0601_/a_150_297# net51 _0601_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4096 _0532_/a_81_21# _0198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4097 _0532_/a_299_297# _0198_ _0532_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4098 VPWR _0532_/a_81_21# _0146_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4099 VPWR net218 _0532_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4100 VGND _0532_/a_81_21# _0146_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4101 VGND _0195_ _0532_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4102 _0532_/a_299_297# _0195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4103 _0532_/a_384_47# net218 _0532_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4104 comp0.B\[15\] _1015_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4105 _1015_/a_891_413# _1015_/a_193_47# _1015_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4106 _1015_/a_561_413# _1015_/a_27_47# _1015_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4107 VPWR net101 _1015_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4108 comp0.B\[15\] _1015_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4109 _1015_/a_381_47# _0113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4110 VGND _1015_/a_634_159# _1015_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4111 VPWR _1015_/a_891_413# _1015_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4112 _1015_/a_466_413# _1015_/a_193_47# _1015_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4113 VPWR _1015_/a_634_159# _1015_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4114 _1015_/a_634_159# _1015_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4115 _1015_/a_634_159# _1015_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4116 _1015_/a_975_413# _1015_/a_193_47# _1015_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4117 VGND _1015_/a_1059_315# _1015_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4118 _1015_/a_193_47# _1015_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4119 _1015_/a_891_413# _1015_/a_27_47# _1015_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4120 _1015_/a_592_47# _1015_/a_193_47# _1015_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4121 VPWR _1015_/a_1059_315# _1015_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4122 _1015_/a_1017_47# _1015_/a_27_47# _1015_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4123 _1015_/a_193_47# _1015_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4124 _1015_/a_466_413# _1015_/a_27_47# _1015_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4125 VGND _1015_/a_891_413# _1015_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4126 _1015_/a_381_47# _0113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4127 VGND net101 _1015_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4128 net84 clknet_1_0__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4129 VGND clknet_1_0__leaf__0459_ net84 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4130 net84 clknet_1_0__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4131 VPWR clknet_1_0__leaf__0459_ net84 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4132 VPWR clknet_0__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X4133 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X4134 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4135 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4136 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4137 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4138 clkbuf_1_1__f__0461_/a_110_47# clknet_0__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4139 clkbuf_1_1__f__0461_/a_110_47# clknet_0__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X4140 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X4141 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4142 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4143 clkbuf_1_1__f__0461_/a_110_47# clknet_0__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4144 VGND clknet_0__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4145 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4146 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4147 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4148 VGND clknet_0__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4149 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4150 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4151 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4152 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4153 clkbuf_1_1__f__0461_/a_110_47# clknet_0__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4154 VPWR clknet_0__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4155 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4156 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4157 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4158 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4159 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4160 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4161 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4162 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4163 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4164 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4165 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4166 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4167 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4168 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4169 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4170 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4171 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4176 _0515_/a_81_21# _0189_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4177 _0515_/a_299_297# _0189_ _0515_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4178 VPWR _0515_/a_81_21# _0154_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4179 VPWR net181 _0515_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4180 VGND _0515_/a_81_21# _0154_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4181 VGND _0179_ _0515_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4182 _0515_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4183 _0515_/a_384_47# net181 _0515_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4186 net40 _0995_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4187 _0995_/a_891_413# _0995_/a_193_47# _0995_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4188 _0995_/a_561_413# _0995_/a_27_47# _0995_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4189 VPWR net81 _0995_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4190 net40 _0995_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4191 _0995_/a_381_47# _0093_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4192 VGND _0995_/a_634_159# _0995_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4193 VPWR _0995_/a_891_413# _0995_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4194 _0995_/a_466_413# _0995_/a_193_47# _0995_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4195 VPWR _0995_/a_634_159# _0995_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4196 _0995_/a_634_159# _0995_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4197 _0995_/a_634_159# _0995_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4198 _0995_/a_975_413# _0995_/a_193_47# _0995_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4199 VGND _0995_/a_1059_315# _0995_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4200 _0995_/a_193_47# _0995_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4201 _0995_/a_891_413# _0995_/a_27_47# _0995_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4202 _0995_/a_592_47# _0995_/a_193_47# _0995_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4203 VPWR _0995_/a_1059_315# _0995_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4204 _0995_/a_1017_47# _0995_/a_27_47# _0995_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4205 _0995_/a_193_47# _0995_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4206 _0995_/a_466_413# _0995_/a_27_47# _0995_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4207 VGND _0995_/a_891_413# _0995_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4208 _0995_/a_381_47# _0093_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4209 VGND net81 _0995_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4210 VPWR _0463_ clkbuf_0__0463_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X4211 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X4212 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4213 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4214 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4215 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4216 clkbuf_0__0463_/a_110_47# _0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4217 clkbuf_0__0463_/a_110_47# _0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X4218 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X4219 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4220 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4221 clkbuf_0__0463_/a_110_47# _0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4222 VGND _0463_ clkbuf_0__0463_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4223 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4224 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4225 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4226 VGND _0463_ clkbuf_0__0463_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4227 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4228 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4229 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4230 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4231 clkbuf_0__0463_/a_110_47# _0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4232 VPWR _0463_ clkbuf_0__0463_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4233 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4234 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4235 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4236 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4237 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4238 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4239 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4240 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4241 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4242 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4243 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4244 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4245 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4246 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4247 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4248 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4249 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4250 _0397_ _0780_/a_35_297# _0780_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X4251 _0397_ _0308_ _0780_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X4252 _0780_/a_35_297# _0308_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X4253 _0780_/a_117_297# _0308_ _0780_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X4254 VPWR _0308_ _0780_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4255 VGND _0387_ _0780_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4256 VGND _0780_/a_35_297# _0397_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4257 _0780_/a_285_297# _0387_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4258 VPWR _0387_ _0780_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4259 _0780_/a_285_47# _0387_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4262 VPWR input5/a_75_212# net5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4263 input5/a_75_212# A[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4264 input5/a_75_212# A[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4265 VGND input5/a_75_212# net5 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4266 VPWR _0466_ _0978_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X4267 _0978_/a_27_297# _0481_ _0978_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X4268 VGND _0466_ _0978_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X4269 _0168_ _0978_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4270 _0978_/a_27_297# _0481_ _0978_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X4271 _0978_/a_109_297# net226 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4272 _0978_/a_373_47# net226 _0978_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4273 _0168_ _0978_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4274 _0978_/a_109_297# _0488_ _0978_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4275 _0978_/a_109_47# _0488_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4276 VPWR _0248_ _0384_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.53 ps=5.06 w=1 l=0.15
X4277 _0384_ _0236_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4278 _0763_/a_193_47# _0248_ _0763_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1755 ps=1.84 w=0.65 l=0.15
X4279 _0384_ _0236_ _0763_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4280 _0384_ _0372_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4281 _0763_/a_109_47# _0372_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4282 VPWR _0350_ _0439_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4283 _0439_ _0350_ _0832_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4284 _0832_/a_113_47# _0438_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4285 _0439_ _0438_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4286 VPWR _0324_ _0326_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4287 _0326_ _0324_ _0694_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4288 _0694_/a_113_47# _0325_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4289 _0326_ _0325_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4296 acc0.A\[31\] _1031_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4297 _1031_/a_891_413# _1031_/a_193_47# _1031_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4298 _1031_/a_561_413# _1031_/a_27_47# _1031_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4299 VPWR net117 _1031_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4300 acc0.A\[31\] _1031_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4301 _1031_/a_381_47# net163 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4302 VGND _1031_/a_634_159# _1031_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4303 VPWR _1031_/a_891_413# _1031_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4304 _1031_/a_466_413# _1031_/a_193_47# _1031_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4305 VPWR _1031_/a_634_159# _1031_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4306 _1031_/a_634_159# _1031_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4307 _1031_/a_634_159# _1031_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4308 _1031_/a_975_413# _1031_/a_193_47# _1031_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4309 VGND _1031_/a_1059_315# _1031_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4310 _1031_/a_193_47# _1031_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4311 _1031_/a_891_413# _1031_/a_27_47# _1031_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4312 _1031_/a_592_47# _1031_/a_193_47# _1031_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4313 VPWR _1031_/a_1059_315# _1031_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4314 _1031_/a_1017_47# _1031_/a_27_47# _1031_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4315 _1031_/a_193_47# _1031_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4316 _1031_/a_466_413# _1031_/a_27_47# _1031_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4317 VGND _1031_/a_891_413# _1031_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4318 _1031_/a_381_47# net163 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4319 VGND net117 _1031_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4320 VPWR input30/a_75_212# net30 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4321 input30/a_75_212# B[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4322 input30/a_75_212# B[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4323 VGND input30/a_75_212# net30 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4326 _0746_/a_81_21# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4327 _0746_/a_299_297# _0346_ _0746_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4328 VPWR _0746_/a_81_21# _0371_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4329 VPWR _0359_ _0746_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4330 VGND _0746_/a_81_21# _0371_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4331 VGND _0370_ _0746_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4332 _0746_/a_299_297# _0370_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4333 _0746_/a_384_47# _0359_ _0746_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4334 _0815_/a_199_47# _0290_ _0425_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X4335 _0815_/a_113_297# _0401_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X4336 _0425_ _0423_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4337 VPWR _0290_ _0815_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4338 _0815_/a_113_297# _0423_ _0425_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X4339 VGND _0401_ _0815_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4340 _0677_/a_377_297# acc0.A\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X4341 _0677_/a_47_47# net44 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4342 _0677_/a_129_47# net44 _0677_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X4343 _0677_/a_285_47# net44 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X4344 _0309_ _0677_/a_47_47# _0677_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X4345 VGND acc0.A\[17\] _0677_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4346 VPWR acc0.A\[17\] _0677_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4347 VPWR _0677_/a_47_47# _0309_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X4348 _0309_ net44 _0677_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4349 _0677_/a_285_47# acc0.A\[17\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4350 _0600_/a_103_199# _0231_ _0600_/a_253_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.39 ps=3.8 w=0.65 l=0.15
X4351 VPWR _0600_/a_103_199# _0232_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.36 ps=2.72 w=1 l=0.15
X4352 _0600_/a_337_297# _0223_ _0600_/a_253_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.27 ps=2.54 w=1 l=0.15
X4353 _0600_/a_103_199# _0230_ _0600_/a_337_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.425 pd=2.85 as=0 ps=0 w=1 l=0.15
X4354 _0600_/a_253_297# _0225_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4355 VPWR _0231_ _0600_/a_103_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4356 VGND _0600_/a_103_199# _0232_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.234 ps=2.02 w=0.65 l=0.15
X4357 _0600_/a_253_47# _0225_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4358 _0600_/a_253_47# _0230_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4359 VGND _0223_ _0600_/a_253_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4360 VPWR net9 _0531_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X4361 _0531_/a_27_297# _0182_ _0531_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X4362 VGND net9 _0531_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X4363 _0198_ _0531_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4364 _0531_/a_27_297# _0182_ _0531_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X4365 _0531_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4366 _0531_/a_373_47# _0180_ _0531_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4367 _0198_ _0531_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4368 _0531_/a_109_297# net175 _0531_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4369 _0531_/a_109_47# net175 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4372 acc0.A\[0\] _1014_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4373 _1014_/a_891_413# _1014_/a_193_47# _1014_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4374 _1014_/a_561_413# _1014_/a_27_47# _1014_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4375 VPWR net100 _1014_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4376 acc0.A\[0\] _1014_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4377 _1014_/a_381_47# _0112_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4378 VGND _1014_/a_634_159# _1014_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4379 VPWR _1014_/a_891_413# _1014_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4380 _1014_/a_466_413# _1014_/a_193_47# _1014_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4381 VPWR _1014_/a_634_159# _1014_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4382 _1014_/a_634_159# _1014_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4383 _1014_/a_634_159# _1014_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4384 _1014_/a_975_413# _1014_/a_193_47# _1014_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4385 VGND _1014_/a_1059_315# _1014_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4386 _1014_/a_193_47# _1014_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4387 _1014_/a_891_413# _1014_/a_27_47# _1014_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4388 _1014_/a_592_47# _1014_/a_193_47# _1014_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4389 VPWR _1014_/a_1059_315# _1014_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4390 _1014_/a_1017_47# _1014_/a_27_47# _1014_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4391 _1014_/a_193_47# _1014_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4392 _1014_/a_466_413# _1014_/a_27_47# _1014_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4393 VGND _1014_/a_891_413# _1014_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4394 _1014_/a_381_47# _0112_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4395 VGND net100 _1014_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4396 VGND _0350_ _0729_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4397 _0729_/a_68_297# net242 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4398 _0358_ _0729_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4399 VPWR _0350_ _0729_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4400 _0358_ _0729_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4401 _0729_/a_150_297# net242 _0729_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4402 net141 clknet_1_1__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4403 VGND clknet_1_1__leaf__0465_ net141 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4404 net141 clknet_1_1__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4405 VPWR clknet_1_1__leaf__0465_ net141 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4406 VPWR clknet_0__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X4407 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X4408 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4409 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4410 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4411 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4412 clkbuf_1_1__f__0460_/a_110_47# clknet_0__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4413 clkbuf_1_1__f__0460_/a_110_47# clknet_0__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X4414 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X4415 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4416 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4417 clkbuf_1_1__f__0460_/a_110_47# clknet_0__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4418 VGND clknet_0__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4419 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4420 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4421 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4422 VGND clknet_0__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4423 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4424 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4425 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4426 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4427 clkbuf_1_1__f__0460_/a_110_47# clknet_0__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4428 VPWR clknet_0__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4429 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4430 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4431 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4432 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4433 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4434 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4435 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4436 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4437 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4438 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4439 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4440 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4441 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4442 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4443 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4444 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4445 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4446 net71 clknet_1_0__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4447 VGND clknet_1_0__leaf__0458_ net71 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4448 net71 clknet_1_0__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4449 VPWR clknet_1_0__leaf__0458_ net71 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4454 net88 clknet_1_0__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4455 VGND clknet_1_0__leaf__0460_ net88 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4456 net88 clknet_1_0__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4457 VPWR clknet_1_0__leaf__0460_ net88 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4460 VPWR net2 _0514_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X4461 _0514_/a_27_297# _0186_ _0514_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X4462 VGND net2 _0514_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X4463 _0189_ _0514_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4464 _0514_/a_27_297# _0186_ _0514_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X4465 _0514_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4466 _0514_/a_373_47# _0181_ _0514_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4467 _0189_ _0514_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4468 _0514_/a_109_297# acc0.A\[10\] _0514_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4469 _0514_/a_109_47# acc0.A\[10\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4476 net122 clknet_1_1__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4477 VGND clknet_1_1__leaf__0463_ net122 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4478 net122 clknet_1_1__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4479 VPWR clknet_1_1__leaf__0463_ net122 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4480 net136 clknet_1_0__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4481 VGND clknet_1_0__leaf__0464_ net136 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4482 net136 clknet_1_0__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4483 VPWR clknet_1_0__leaf__0464_ net136 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4484 net39 _0994_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4485 _0994_/a_891_413# _0994_/a_193_47# _0994_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4486 _0994_/a_561_413# _0994_/a_27_47# _0994_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4487 VPWR net80 _0994_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4488 net39 _0994_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4489 _0994_/a_381_47# _0092_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4490 VGND _0994_/a_634_159# _0994_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4491 VPWR _0994_/a_891_413# _0994_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4492 _0994_/a_466_413# _0994_/a_193_47# _0994_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4493 VPWR _0994_/a_634_159# _0994_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4494 _0994_/a_634_159# _0994_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4495 _0994_/a_634_159# _0994_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4496 _0994_/a_975_413# _0994_/a_193_47# _0994_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4497 VGND _0994_/a_1059_315# _0994_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4498 _0994_/a_193_47# _0994_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4499 _0994_/a_891_413# _0994_/a_27_47# _0994_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4500 _0994_/a_592_47# _0994_/a_193_47# _0994_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4501 VPWR _0994_/a_1059_315# _0994_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4502 _0994_/a_1017_47# _0994_/a_27_47# _0994_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4503 _0994_/a_193_47# _0994_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4504 _0994_/a_466_413# _0994_/a_27_47# _0994_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4505 VGND _0994_/a_891_413# _0994_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4506 _0994_/a_381_47# _0092_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4507 VGND net80 _0994_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4508 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4509 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4510 VPWR _0462_ clkbuf_0__0462_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X4511 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X4512 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4513 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4514 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4515 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4516 clkbuf_0__0462_/a_110_47# _0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4517 clkbuf_0__0462_/a_110_47# _0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X4518 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X4519 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4520 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4521 clkbuf_0__0462_/a_110_47# _0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4522 VGND _0462_ clkbuf_0__0462_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4523 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4524 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4525 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4526 VGND _0462_ clkbuf_0__0462_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4527 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4528 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4529 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4530 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4531 clkbuf_0__0462_/a_110_47# _0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4532 VPWR _0462_ clkbuf_0__0462_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4533 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4534 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4535 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4536 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4537 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4538 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4539 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4540 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4541 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4542 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4543 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4544 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4545 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4546 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4547 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4548 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4549 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4552 VPWR input6/a_75_212# net6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4553 input6/a_75_212# A[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4554 input6/a_75_212# A[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4555 VGND input6/a_75_212# net6 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4556 VPWR _0977_/a_75_212# _0167_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4557 _0977_/a_75_212# _0489_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4558 _0977_/a_75_212# _0489_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4559 VGND _0977_/a_75_212# _0167_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4562 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4565 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4566 _0438_ _0831_/a_35_297# _0831_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X4567 _0438_ _0434_ _0831_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X4568 _0831_/a_35_297# _0434_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X4569 _0831_/a_117_297# _0434_ _0831_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X4570 VPWR _0434_ _0831_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4571 VGND _0253_ _0831_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4572 VGND _0831_/a_35_297# _0438_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4573 _0831_/a_285_297# _0253_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4574 VPWR _0253_ _0831_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4575 _0831_/a_285_47# _0253_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4576 VGND _0369_ _0762_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X4577 _0762_/a_510_47# _0383_ _0762_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X4578 _0762_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X4579 VPWR _0383_ _0762_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4580 _0762_/a_79_21# net213 _0762_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X4581 _0762_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4582 _0762_/a_79_21# _0352_ _0762_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X4583 VPWR _0762_/a_79_21# _0101_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4584 VGND _0762_/a_79_21# _0101_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4585 _0762_/a_215_47# net213 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4586 VGND acc0.A\[24\] _0693_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4587 _0693_/a_68_297# net52 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4588 _0325_ _0693_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4589 VPWR acc0.A\[24\] _0693_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4590 _0325_ _0693_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4591 _0693_/a_150_297# net52 _0693_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4596 acc0.A\[30\] _1030_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4597 _1030_/a_891_413# _1030_/a_193_47# _1030_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4598 _1030_/a_561_413# _1030_/a_27_47# _1030_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4599 VPWR net116 _1030_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4600 acc0.A\[30\] _1030_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4601 _1030_/a_381_47# net209 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4602 VGND _1030_/a_634_159# _1030_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4603 VPWR _1030_/a_891_413# _1030_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4604 _1030_/a_466_413# _1030_/a_193_47# _1030_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4605 VPWR _1030_/a_634_159# _1030_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4606 _1030_/a_634_159# _1030_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4607 _1030_/a_634_159# _1030_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4608 _1030_/a_975_413# _1030_/a_193_47# _1030_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4609 VGND _1030_/a_1059_315# _1030_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4610 _1030_/a_193_47# _1030_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4611 _1030_/a_891_413# _1030_/a_27_47# _1030_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4612 _1030_/a_592_47# _1030_/a_193_47# _1030_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4613 VPWR _1030_/a_1059_315# _1030_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4614 _1030_/a_1017_47# _1030_/a_27_47# _1030_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4615 _1030_/a_193_47# _1030_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4616 _1030_/a_466_413# _1030_/a_27_47# _1030_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4617 VGND _1030_/a_891_413# _1030_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4618 _1030_/a_381_47# net209 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4619 VGND net116 _1030_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4620 VPWR input20/a_75_212# net20 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4621 input20/a_75_212# B[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4622 input20/a_75_212# B[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4623 VGND input20/a_75_212# net20 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4624 VPWR input31/a_75_212# net31 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4625 input31/a_75_212# B[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4626 input31/a_75_212# B[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4627 VGND input31/a_75_212# net31 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4628 VPWR _0423_ _0814_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2415 ps=2.83 w=0.42 l=0.15
X4629 VPWR _0401_ _0814_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4630 _0814_/a_181_47# _0290_ _0814_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0882 pd=1.26 as=0.0882 ps=1.26 w=0.42 l=0.15
X4631 VGND _0401_ _0814_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4632 _0814_/a_27_47# _0290_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4633 _0424_ _0814_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4634 _0424_ _0814_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4635 _0814_/a_109_47# _0423_ _0814_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4636 VPWR _0250_ _0370_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.53 ps=5.06 w=1 l=0.15
X4637 _0370_ _0326_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4638 _0745_/a_193_47# _0250_ _0745_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1755 ps=1.84 w=0.65 l=0.15
X4639 _0370_ _0326_ _0745_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4640 _0370_ _0312_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4641 _0745_/a_109_47# _0312_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4642 VPWR _0306_ _0308_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4643 _0308_ _0306_ _0676_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4644 _0676_/a_113_47# _0307_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4645 _0308_ _0307_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4648 _0530_/a_81_21# _0197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4649 _0530_/a_299_297# _0197_ _0530_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4650 VPWR _0530_/a_81_21# _0147_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4651 VPWR net175 _0530_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4652 VGND _0530_/a_81_21# _0147_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4653 VGND _0195_ _0530_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4654 _0530_/a_299_297# _0195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4655 _0530_/a_384_47# net175 _0530_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4656 net60 _1013_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4657 _1013_/a_891_413# _1013_/a_193_47# _1013_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4658 _1013_/a_561_413# _1013_/a_27_47# _1013_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4659 VPWR net99 _1013_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4660 net60 _1013_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4661 _1013_/a_381_47# _0111_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4662 VGND _1013_/a_634_159# _1013_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4663 VPWR _1013_/a_891_413# _1013_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4664 _1013_/a_466_413# _1013_/a_193_47# _1013_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4665 VPWR _1013_/a_634_159# _1013_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4666 _1013_/a_634_159# _1013_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4667 _1013_/a_634_159# _1013_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4668 _1013_/a_975_413# _1013_/a_193_47# _1013_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4669 VGND _1013_/a_1059_315# _1013_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4670 _1013_/a_193_47# _1013_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4671 _1013_/a_891_413# _1013_/a_27_47# _1013_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4672 _1013_/a_592_47# _1013_/a_193_47# _1013_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4673 VPWR _1013_/a_1059_315# _1013_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4674 _1013_/a_1017_47# _1013_/a_27_47# _1013_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4675 _1013_/a_193_47# _1013_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4676 _1013_/a_466_413# _1013_/a_27_47# _1013_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4677 VGND _1013_/a_891_413# _1013_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4678 _1013_/a_381_47# _0111_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4679 VGND net99 _1013_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4680 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4681 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4682 VPWR _0356_ _0728_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4683 _0357_ _0728_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X4684 VGND _0356_ _0728_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4685 _0728_/a_59_75# _0333_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4686 _0357_ _0728_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X4687 _0728_/a_145_75# _0333_ _0728_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X4688 VGND acc0.A\[8\] _0659_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4689 _0659_/a_68_297# net66 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4690 _0291_ _0659_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4691 VPWR acc0.A\[8\] _0659_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4692 _0291_ _0659_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4693 _0659_/a_150_297# net66 _0659_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4694 _0513_/a_81_21# _0188_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4695 _0513_/a_299_297# _0188_ _0513_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4696 VPWR _0513_/a_81_21# _0155_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4697 VPWR net188 _0513_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4698 VGND _0513_/a_81_21# _0155_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4699 VGND _0179_ _0513_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4700 _0513_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4701 _0513_/a_384_47# net188 _0513_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4703 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4708 net38 _0993_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4709 _0993_/a_891_413# _0993_/a_193_47# _0993_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4710 _0993_/a_561_413# _0993_/a_27_47# _0993_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4711 VPWR net79 _0993_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4712 net38 _0993_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4713 _0993_/a_381_47# _0091_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4714 VGND _0993_/a_634_159# _0993_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4715 VPWR _0993_/a_891_413# _0993_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4716 _0993_/a_466_413# _0993_/a_193_47# _0993_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4717 VPWR _0993_/a_634_159# _0993_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4718 _0993_/a_634_159# _0993_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4719 _0993_/a_634_159# _0993_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4720 _0993_/a_975_413# _0993_/a_193_47# _0993_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4721 VGND _0993_/a_1059_315# _0993_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4722 _0993_/a_193_47# _0993_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4723 _0993_/a_891_413# _0993_/a_27_47# _0993_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4724 _0993_/a_592_47# _0993_/a_193_47# _0993_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4725 VPWR _0993_/a_1059_315# _0993_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4726 _0993_/a_1017_47# _0993_/a_27_47# _0993_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4727 _0993_/a_193_47# _0993_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4728 _0993_/a_466_413# _0993_/a_27_47# _0993_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4729 VGND _0993_/a_891_413# _0993_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4730 _0993_/a_381_47# _0091_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4731 VGND net79 _0993_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4732 VPWR _0461_ clkbuf_0__0461_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X4733 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X4734 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4735 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4736 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4737 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4738 clkbuf_0__0461_/a_110_47# _0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4739 clkbuf_0__0461_/a_110_47# _0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X4740 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X4741 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4742 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4743 clkbuf_0__0461_/a_110_47# _0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4744 VGND _0461_ clkbuf_0__0461_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4745 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4746 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4747 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4748 VGND _0461_ clkbuf_0__0461_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4749 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4750 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4751 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4752 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4753 clkbuf_0__0461_/a_110_47# _0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4754 VPWR _0461_ clkbuf_0__0461_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4755 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4756 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4757 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4758 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4759 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4760 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4761 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4762 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4763 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4764 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4765 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4766 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4767 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4768 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4769 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4770 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4771 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4774 VPWR input7/a_75_212# net7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4775 input7/a_75_212# A[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4776 input7/a_75_212# A[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4777 VGND input7/a_75_212# net7 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4778 VPWR _0976_/a_505_21# _0976_/a_535_374# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4779 _0976_/a_505_21# control0.count\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4780 _0976_/a_218_374# control0.count\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4781 VGND _0976_/a_505_21# _0976_/a_439_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4782 _0976_/a_76_199# _0488_ _0976_/a_218_374# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4783 _0976_/a_505_21# control0.count\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X4784 _0976_/a_439_47# _0488_ _0976_/a_76_199# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4785 _0976_/a_535_374# _0466_ _0976_/a_76_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X4786 _0976_/a_76_199# _0466_ _0976_/a_218_47# VGND sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4787 _0976_/a_218_47# control0.count\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4788 VPWR _0976_/a_76_199# _0489_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X4789 VGND _0976_/a_76_199# _0489_ VGND sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4792 VGND _0369_ _0830_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X4793 _0830_/a_510_47# _0437_ _0830_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X4794 _0830_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X4795 VPWR _0437_ _0830_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4796 _0830_/a_79_21# net212 _0830_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X4797 _0830_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4798 _0830_/a_79_21# _0399_ _0830_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X4799 VPWR _0830_/a_79_21# _0087_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4800 VGND _0830_/a_79_21# _0087_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4801 _0830_/a_215_47# net212 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4802 VPWR _0219_ _0383_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4803 _0383_ _0219_ _0761_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4804 _0761_/a_113_47# _0382_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4805 _0383_ _0382_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4806 VPWR acc0.A\[24\] _0324_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4807 _0324_ acc0.A\[24\] _0692_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4808 _0692_/a_113_47# net52 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4809 _0324_ net52 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4812 VPWR _0959_/a_80_21# _0160_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X4813 _0959_/a_80_21# _0477_ _0959_/a_472_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.31 ps=2.62 w=1 l=0.15
X4814 VPWR _0467_ _0959_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.545 ps=5.09 w=1 l=0.15
X4815 VGND _0470_ _0959_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.35425 ps=3.69 w=0.65 l=0.15
X4816 VGND _0959_/a_80_21# _0160_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X4817 _0959_/a_300_47# _0467_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X4818 _0959_/a_217_297# net33 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4819 _0959_/a_80_21# net33 _0959_/a_300_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4820 _0959_/a_472_297# _0470_ _0959_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4821 _0959_/a_80_21# _0477_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4824 net95 clknet_1_1__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4825 VGND clknet_1_1__leaf__0460_ net95 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4826 net95 clknet_1_1__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4827 VPWR clknet_1_1__leaf__0460_ net95 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4828 VPWR input10/a_75_212# net10 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4829 input10/a_75_212# A[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4830 input10/a_75_212# A[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4831 VGND input10/a_75_212# net10 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4832 VPWR input21/a_75_212# net21 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4833 input21/a_75_212# B[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4834 input21/a_75_212# B[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4835 VGND input21/a_75_212# net21 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4836 VPWR input32/a_75_212# net32 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4837 input32/a_75_212# B[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4838 input32/a_75_212# B[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4839 VGND input32/a_75_212# net32 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4840 VPWR _0288_ _0813_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X4841 VGND _0288_ _0423_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4842 _0813_/a_109_297# _0289_ _0423_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4843 _0423_ _0289_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4844 VPWR _0350_ _0744_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X4845 VGND _0744_/a_27_47# _0369_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X4846 VGND _0744_/a_27_47# _0369_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4847 _0369_ _0744_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X4848 _0369_ _0744_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4849 VGND _0350_ _0744_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X4850 VPWR _0744_/a_27_47# _0369_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4851 _0369_ _0744_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4852 _0369_ _0744_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4853 VPWR _0744_/a_27_47# _0369_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4854 VGND acc0.A\[16\] _0675_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4855 _0675_/a_68_297# net43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4856 _0307_ _0675_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4857 VPWR acc0.A\[16\] _0675_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4858 _0307_ _0675_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4859 _0675_/a_150_297# net43 _0675_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4860 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4861 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4862 net59 _1012_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4863 _1012_/a_891_413# _1012_/a_193_47# _1012_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4864 _1012_/a_561_413# _1012_/a_27_47# _1012_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4865 VPWR net98 _1012_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4866 net59 _1012_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4867 _1012_/a_381_47# _0110_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4868 VGND _1012_/a_634_159# _1012_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4869 VPWR _1012_/a_891_413# _1012_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4870 _1012_/a_466_413# _1012_/a_193_47# _1012_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4871 VPWR _1012_/a_634_159# _1012_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4872 _1012_/a_634_159# _1012_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4873 _1012_/a_634_159# _1012_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4874 _1012_/a_975_413# _1012_/a_193_47# _1012_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4875 VGND _1012_/a_1059_315# _1012_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4876 _1012_/a_193_47# _1012_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4877 _1012_/a_891_413# _1012_/a_27_47# _1012_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4878 _1012_/a_592_47# _1012_/a_193_47# _1012_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4879 VPWR _1012_/a_1059_315# _1012_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4880 _1012_/a_1017_47# _1012_/a_27_47# _1012_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4881 _1012_/a_193_47# _1012_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4882 _1012_/a_466_413# _1012_/a_27_47# _1012_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4883 VGND _1012_/a_891_413# _1012_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4884 _1012_/a_381_47# _0110_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4885 VGND net98 _1012_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4886 _0356_ _0327_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4887 VPWR _0332_ _0356_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X4888 VPWR _0329_ _0356_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4889 _0727_/a_193_47# _0329_ _0727_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4890 _0356_ _0332_ _0727_/a_277_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X4891 _0727_/a_277_47# _0327_ _0727_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4892 _0356_ _0330_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4893 _0727_/a_109_47# _0330_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4894 VPWR acc0.A\[8\] _0290_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4895 _0290_ acc0.A\[8\] _0658_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4896 _0658_/a_113_47# net66 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4897 _0290_ net66 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4898 VPWR acc0.A\[28\] _0221_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4899 _0221_ acc0.A\[28\] _0589_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4900 _0589_/a_113_47# net56 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4901 _0221_ net56 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4902 VPWR net3 _0512_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X4903 _0512_/a_27_297# _0186_ _0512_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X4904 VGND net3 _0512_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X4905 _0188_ _0512_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4906 _0512_/a_27_297# _0186_ _0512_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X4907 _0512_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4908 _0512_/a_373_47# _0181_ _0512_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4909 _0188_ _0512_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4910 _0512_/a_109_297# acc0.A\[11\] _0512_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4911 _0512_/a_109_47# acc0.A\[11\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4912 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4915 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4916 net37 _0992_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4917 _0992_/a_891_413# _0992_/a_193_47# _0992_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4918 _0992_/a_561_413# _0992_/a_27_47# _0992_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4919 VPWR net78 _0992_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4920 net37 _0992_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4921 _0992_/a_381_47# _0090_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4922 VGND _0992_/a_634_159# _0992_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4923 VPWR _0992_/a_891_413# _0992_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4924 _0992_/a_466_413# _0992_/a_193_47# _0992_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4925 VPWR _0992_/a_634_159# _0992_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4926 _0992_/a_634_159# _0992_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4927 _0992_/a_634_159# _0992_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4928 _0992_/a_975_413# _0992_/a_193_47# _0992_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4929 VGND _0992_/a_1059_315# _0992_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4930 _0992_/a_193_47# _0992_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4931 _0992_/a_891_413# _0992_/a_27_47# _0992_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4932 _0992_/a_592_47# _0992_/a_193_47# _0992_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4933 VPWR _0992_/a_1059_315# _0992_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4934 _0992_/a_1017_47# _0992_/a_27_47# _0992_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4935 _0992_/a_193_47# _0992_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4936 _0992_/a_466_413# _0992_/a_27_47# _0992_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4937 VGND _0992_/a_891_413# _0992_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4938 _0992_/a_381_47# _0090_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4939 VGND net78 _0992_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4940 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4941 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4942 VPWR _0460_ clkbuf_0__0460_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X4943 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X4944 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4945 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4946 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4947 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4948 clkbuf_0__0460_/a_110_47# _0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4949 clkbuf_0__0460_/a_110_47# _0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X4950 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X4951 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4952 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4953 clkbuf_0__0460_/a_110_47# _0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4954 VGND _0460_ clkbuf_0__0460_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4955 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4956 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4957 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4958 VGND _0460_ clkbuf_0__0460_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4959 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4960 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4961 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4962 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4963 clkbuf_0__0460_/a_110_47# _0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4964 VPWR _0460_ clkbuf_0__0460_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4965 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4966 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4967 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4968 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4969 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4970 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4971 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4972 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4973 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4974 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4975 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4976 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4977 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4978 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4979 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4980 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4981 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4984 net127 clknet_1_0__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4985 VGND clknet_1_0__leaf__0463_ net127 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4986 net127 clknet_1_0__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4987 VPWR clknet_1_0__leaf__0463_ net127 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4988 VPWR input8/a_75_212# net8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4989 input8/a_75_212# A[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4990 input8/a_75_212# A[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4991 VGND input8/a_75_212# net8 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4992 VPWR _0486_ _0975_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4993 _0488_ _0975_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X4994 VGND _0486_ _0975_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4995 _0975_/a_59_75# control0.state\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4996 _0488_ _0975_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X4997 _0975_/a_145_75# control0.state\[2\] _0975_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X4998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4999 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5000 _0760_/a_377_297# _0237_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X5001 _0760_/a_47_47# _0381_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5002 _0760_/a_129_47# _0381_ _0760_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X5003 _0760_/a_285_47# _0381_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X5004 _0382_ _0760_/a_47_47# _0760_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X5005 VGND _0237_ _0760_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5006 VPWR _0237_ _0760_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5007 VPWR _0760_/a_47_47# _0382_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X5008 _0382_ _0381_ _0760_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5009 _0760_/a_285_47# _0237_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5010 VGND _0315_ _0691_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5011 _0691_/a_68_297# _0322_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5012 _0323_ _0691_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5013 VPWR _0315_ _0691_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X5014 _0323_ _0691_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X5015 _0691_/a_150_297# _0322_ _0691_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5017 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5018 _0958_/a_27_47# _0476_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5019 _0958_/a_197_47# _0471_ _0958_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X5020 _0477_ _0958_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X5021 _0958_/a_303_47# _0476_ _0958_/a_197_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X5022 _0958_/a_27_47# control0.state\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5023 VPWR _0468_ _0958_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X5024 VGND _0468_ _0958_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0.19627 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X5025 VPWR _0471_ _0958_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X5026 _0477_ _0958_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.19627 ps=1.33 w=0.65 l=0.15
X5027 _0958_/a_109_47# control0.state\[1\] _0958_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X5028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5032 _0743_/a_240_47# net237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X5033 _0105_ _0743_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X5034 VGND _0219_ _0743_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5035 _0743_/a_51_297# _0368_ _0743_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X5036 _0743_/a_149_47# _0345_ _0743_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X5037 _0743_/a_240_47# _0367_ _0743_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5038 VPWR _0219_ _0743_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5039 _0105_ _0743_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X5040 _0743_/a_149_47# _0368_ _0743_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5041 _0743_/a_245_297# _0367_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5042 VPWR _0345_ _0743_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5043 _0743_/a_512_297# net237 _0743_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5044 VPWR input11/a_75_212# net11 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5045 input11/a_75_212# A[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5046 input11/a_75_212# A[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5047 VGND input11/a_75_212# net11 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5048 VPWR input22/a_75_212# net22 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5049 input22/a_75_212# B[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5050 input22/a_75_212# B[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5051 VGND input22/a_75_212# net22 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5052 VPWR input33/a_75_212# net33 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5053 input33/a_75_212# init VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5054 input33/a_75_212# init VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5055 VGND input33/a_75_212# net33 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5056 VGND _0369_ _0812_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X5057 _0812_/a_510_47# _0422_ _0812_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X5058 _0812_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X5059 VPWR _0422_ _0812_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5060 _0812_/a_79_21# net217 _0812_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X5061 _0812_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5062 _0812_/a_79_21# _0399_ _0812_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X5063 VPWR _0812_/a_79_21# _0090_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5064 VGND _0812_/a_79_21# _0090_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5065 _0812_/a_215_47# net217 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5066 VPWR acc0.A\[16\] _0306_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5067 _0306_ acc0.A\[16\] _0674_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5068 _0674_/a_113_47# net43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5069 _0306_ net43 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5070 VPWR clknet_0_clk clkbuf_1_0__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X5071 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X5072 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5073 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5074 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5075 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5076 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5077 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X5078 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X5079 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5080 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5081 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5082 VGND clknet_0_clk clkbuf_1_0__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5083 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5084 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5085 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5086 VGND clknet_0_clk clkbuf_1_0__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5087 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5088 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5089 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5090 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5091 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5092 VPWR clknet_0_clk clkbuf_1_0__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5093 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5094 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5095 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5096 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5097 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5098 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5099 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5100 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5101 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5102 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5103 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5104 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5105 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5106 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5107 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5108 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5109 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5112 net99 clknet_1_1__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5113 VGND clknet_1_1__leaf__0461_ net99 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5114 net99 clknet_1_1__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5115 VPWR clknet_1_1__leaf__0461_ net99 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5116 net57 _1011_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5117 _1011_/a_891_413# _1011_/a_193_47# _1011_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5118 _1011_/a_561_413# _1011_/a_27_47# _1011_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5119 VPWR net97 _1011_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5120 net57 _1011_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5121 _1011_/a_381_47# _0109_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5122 VGND _1011_/a_634_159# _1011_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5123 VPWR _1011_/a_891_413# _1011_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5124 _1011_/a_466_413# _1011_/a_193_47# _1011_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5125 VPWR _1011_/a_634_159# _1011_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5126 _1011_/a_634_159# _1011_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5127 _1011_/a_634_159# _1011_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5128 _1011_/a_975_413# _1011_/a_193_47# _1011_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5129 VGND _1011_/a_1059_315# _1011_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5130 _1011_/a_193_47# _1011_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5131 _1011_/a_891_413# _1011_/a_27_47# _1011_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5132 _1011_/a_592_47# _1011_/a_193_47# _1011_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5133 VPWR _1011_/a_1059_315# _1011_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5134 _1011_/a_1017_47# _1011_/a_27_47# _1011_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5135 _1011_/a_193_47# _1011_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5136 _1011_/a_466_413# _1011_/a_27_47# _1011_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5137 VGND _1011_/a_891_413# _1011_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5138 _1011_/a_381_47# _0109_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5139 VGND net97 _1011_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5140 _0726_/a_240_47# net227 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X5141 _0109_ _0726_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X5142 VGND _0219_ _0726_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5143 _0726_/a_51_297# _0355_ _0726_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X5144 _0726_/a_149_47# _0345_ _0726_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X5145 _0726_/a_240_47# _0354_ _0726_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5146 VPWR _0219_ _0726_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5147 _0109_ _0726_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X5148 _0726_/a_149_47# _0355_ _0726_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5149 _0726_/a_245_297# _0354_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5150 VPWR _0345_ _0726_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5151 _0726_/a_512_297# net227 _0726_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5152 VPWR acc0.A\[30\] _0220_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5153 _0220_ acc0.A\[30\] _0588_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5154 _0588_/a_113_47# net59 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5155 _0220_ net59 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5158 VPWR acc0.A\[9\] _0657_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5159 VGND acc0.A\[9\] _0289_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5160 _0657_/a_109_297# net67 _0289_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5161 _0289_ net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5162 _0511_/a_81_21# _0187_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X5163 _0511_/a_299_297# _0187_ _0511_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X5164 VPWR _0511_/a_81_21# _0156_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5165 VPWR net192 _0511_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5166 VGND _0511_/a_81_21# _0156_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5167 VGND _0179_ _0511_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X5168 _0511_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5169 _0511_/a_384_47# net192 _0511_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5170 net80 clknet_1_1__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5171 VGND clknet_1_1__leaf__0459_ net80 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5172 net80 clknet_1_1__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5173 VPWR clknet_1_1__leaf__0459_ net80 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5174 VPWR acc0.A\[31\] _0341_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5175 _0341_ acc0.A\[31\] _0709_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5176 _0709_/a_113_47# net60 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5177 _0341_ net60 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5178 net67 _0991_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5179 _0991_/a_891_413# _0991_/a_193_47# _0991_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5180 _0991_/a_561_413# _0991_/a_27_47# _0991_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5181 VPWR net77 _0991_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5182 net67 _0991_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5183 _0991_/a_381_47# _0089_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5184 VGND _0991_/a_634_159# _0991_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5185 VPWR _0991_/a_891_413# _0991_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5186 _0991_/a_466_413# _0991_/a_193_47# _0991_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5187 VPWR _0991_/a_634_159# _0991_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5188 _0991_/a_634_159# _0991_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5189 _0991_/a_634_159# _0991_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5190 _0991_/a_975_413# _0991_/a_193_47# _0991_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5191 VGND _0991_/a_1059_315# _0991_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5192 _0991_/a_193_47# _0991_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5193 _0991_/a_891_413# _0991_/a_27_47# _0991_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5194 _0991_/a_592_47# _0991_/a_193_47# _0991_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5195 VPWR _0991_/a_1059_315# _0991_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5196 _0991_/a_1017_47# _0991_/a_27_47# _0991_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5197 _0991_/a_193_47# _0991_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5198 _0991_/a_466_413# _0991_/a_27_47# _0991_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5199 VGND _0991_/a_891_413# _0991_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5200 _0991_/a_381_47# _0089_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5201 VGND net77 _0991_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5202 net114 clknet_1_1__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5203 VGND clknet_1_1__leaf__0462_ net114 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5204 net114 clknet_1_1__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5205 VPWR clknet_1_1__leaf__0462_ net114 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5206 VPWR A[2] input9/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5207 net9 input9/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5208 net9 input9/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5209 VGND A[2] input9/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5210 _0974_/a_222_93# _0468_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5211 VPWR net159 _0974_/a_544_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5212 VGND _0974_/a_79_199# _0166_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5213 _0974_/a_222_93# _0468_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0 ps=0 w=0.42 l=0.15
X5214 VGND _0486_ _0974_/a_448_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.38675 ps=3.79 w=0.65 l=0.15
X5215 _0974_/a_448_47# _0974_/a_222_93# _0974_/a_79_199# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5216 _0974_/a_79_199# _0974_/a_222_93# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0 ps=0 w=1 l=0.15
X5217 _0974_/a_544_297# _0486_ _0974_/a_79_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5218 _0974_/a_448_47# net159 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5219 VPWR _0974_/a_79_199# _0166_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5226 VGND _0318_ _0690_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5227 _0690_/a_68_297# _0321_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5228 _0322_ _0690_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5229 VPWR _0318_ _0690_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X5230 _0322_ _0690_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X5231 _0690_/a_150_297# _0321_ _0690_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5236 VPWR _0475_ _0957_/a_304_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X5237 _0957_/a_304_297# _0472_ _0957_/a_220_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5238 VGND _0474_ _0957_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X5239 _0957_/a_220_297# _0474_ _0957_/a_114_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X5240 _0957_/a_32_297# _0473_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X5241 _0957_/a_32_297# _0472_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5242 VPWR _0957_/a_32_297# _0476_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5243 _0476_ _0957_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5244 VGND _0475_ _0957_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X5245 VPWR _0957_/a_32_297# _0476_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5246 _0476_ _0957_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X5247 _0476_ _0957_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5248 _0476_ _0957_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X5249 _0957_/a_114_297# _0473_ _0957_/a_32_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X5250 VGND _0957_/a_32_297# _0476_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5251 VGND _0957_/a_32_297# _0476_ VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X5252 net74 clknet_1_1__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5253 VGND clknet_1_1__leaf__0458_ net74 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5254 net74 clknet_1_1__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5255 VPWR clknet_1_1__leaf__0458_ net74 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5258 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5259 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5262 _0673_/a_103_199# _0304_ _0673_/a_253_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.39 ps=3.8 w=0.65 l=0.15
X5263 VPWR _0673_/a_103_199# _0305_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.36 ps=2.72 w=1 l=0.15
X5264 _0673_/a_337_297# _0289_ _0673_/a_253_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.27 ps=2.54 w=1 l=0.15
X5265 _0673_/a_103_199# _0295_ _0673_/a_337_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.425 pd=2.85 as=0 ps=0 w=1 l=0.15
X5266 _0673_/a_253_297# _0287_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5267 VPWR _0304_ _0673_/a_103_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5268 VGND _0673_/a_103_199# _0305_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.234 ps=2.02 w=0.65 l=0.15
X5269 _0673_/a_253_47# _0287_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5270 _0673_/a_253_47# _0295_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5271 VGND _0289_ _0673_/a_253_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5272 VPWR input12/a_75_212# net12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5273 input12/a_75_212# A[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5274 input12/a_75_212# A[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5275 VGND input12/a_75_212# net12 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5276 VPWR rst input34/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5277 net34 input34/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5278 net34 input34/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5279 VGND rst input34/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5282 VPWR input23/a_75_212# net23 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5283 input23/a_75_212# B[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5284 input23/a_75_212# B[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5285 VGND input23/a_75_212# net23 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5286 VPWR clknet_0__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X5287 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X5288 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5289 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5290 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5291 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5292 clkbuf_1_0__f__0465_/a_110_47# clknet_0__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5293 clkbuf_1_0__f__0465_/a_110_47# clknet_0__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X5294 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X5295 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5296 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5297 clkbuf_1_0__f__0465_/a_110_47# clknet_0__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5298 VGND clknet_0__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5299 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5300 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5301 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5302 VGND clknet_0__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5303 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5304 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5305 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5306 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5307 clkbuf_1_0__f__0465_/a_110_47# clknet_0__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5308 VPWR clknet_0__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5309 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5310 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5311 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5312 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5313 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5314 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5315 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5316 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5317 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5318 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5319 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5320 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5321 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5322 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5323 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5324 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5325 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5326 _0742_/a_81_21# _0343_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X5327 _0742_/a_299_297# _0343_ _0742_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X5328 VPWR _0742_/a_81_21# _0368_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5329 VPWR _0315_ _0742_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5330 VGND _0742_/a_81_21# _0368_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5331 VGND _0366_ _0742_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X5332 _0742_/a_299_297# _0366_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5333 _0742_/a_384_47# _0315_ _0742_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5334 _0811_/a_81_21# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X5335 _0811_/a_299_297# _0346_ _0811_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X5336 VPWR _0811_/a_81_21# _0422_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5337 VPWR _0402_ _0811_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5338 VGND _0811_/a_81_21# _0422_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5339 VGND _0421_ _0811_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X5340 _0811_/a_299_297# _0421_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5341 _0811_/a_384_47# _0402_ _0811_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5342 net56 _1010_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5343 _1010_/a_891_413# _1010_/a_193_47# _1010_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5344 _1010_/a_561_413# _1010_/a_27_47# _1010_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5345 VPWR net96 _1010_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5346 net56 _1010_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5347 _1010_/a_381_47# _0108_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5348 VGND _1010_/a_634_159# _1010_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5349 VPWR _1010_/a_891_413# _1010_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5350 _1010_/a_466_413# _1010_/a_193_47# _1010_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5351 VPWR _1010_/a_634_159# _1010_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5352 _1010_/a_634_159# _1010_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5353 _1010_/a_634_159# _1010_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5354 _1010_/a_975_413# _1010_/a_193_47# _1010_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5355 VGND _1010_/a_1059_315# _1010_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5356 _1010_/a_193_47# _1010_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5357 _1010_/a_891_413# _1010_/a_27_47# _1010_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5358 _1010_/a_592_47# _1010_/a_193_47# _1010_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5359 VPWR _1010_/a_1059_315# _1010_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5360 _1010_/a_1017_47# _1010_/a_27_47# _1010_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5361 _1010_/a_193_47# _1010_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5362 _1010_/a_466_413# _1010_/a_27_47# _1010_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5363 VGND _1010_/a_891_413# _1010_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5364 _1010_/a_381_47# _0108_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5365 VGND net96 _1010_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5366 VPWR _0725_/a_80_21# _0355_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X5367 _0725_/a_209_297# _0353_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.65 pd=5.3 as=0 ps=0 w=1 l=0.15
X5368 _0725_/a_303_47# _0333_ _0725_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.208 ps=1.94 w=0.65 l=0.15
X5369 _0725_/a_209_47# _0353_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5370 VGND _0725_/a_80_21# _0355_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X5371 VGND _0343_ _0725_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X5372 _0725_/a_80_21# _0221_ _0725_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5373 VPWR _0333_ _0725_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5374 _0725_/a_80_21# _0343_ _0725_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0 ps=0 w=1 l=0.15
X5375 _0725_/a_209_297# _0221_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5376 VPWR net67 _0656_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5377 _0288_ _0656_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X5378 VGND net67 _0656_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5379 _0656_/a_59_75# acc0.A\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5380 _0288_ _0656_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X5381 _0656_/a_145_75# acc0.A\[9\] _0656_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X5382 VPWR _0218_ _0587_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X5383 VGND _0587_/a_27_47# _0219_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X5384 VGND _0587_/a_27_47# _0219_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5385 _0219_ _0587_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X5386 _0219_ _0587_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5387 VGND _0218_ _0587_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X5388 VPWR _0587_/a_27_47# _0219_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5389 _0219_ _0587_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5390 _0219_ _0587_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5391 VPWR _0587_/a_27_47# _0219_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5394 VPWR net4 _0510_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X5395 _0510_/a_27_297# _0186_ _0510_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X5396 VGND net4 _0510_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X5397 _0187_ _0510_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5398 _0510_/a_27_297# _0186_ _0510_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X5399 _0510_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5400 _0510_/a_373_47# _0181_ _0510_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5401 _0187_ _0510_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5402 _0510_/a_109_297# acc0.A\[12\] _0510_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5403 _0510_/a_109_47# acc0.A\[12\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5404 VPWR acc0.A\[5\] hold1/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5405 VGND hold1/a_285_47# hold1/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5406 net148 hold1/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5407 VGND acc0.A\[5\] hold1/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5408 VPWR hold1/a_285_47# hold1/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5409 hold1/a_285_47# hold1/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X5410 hold1/a_285_47# hold1/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X5411 net148 hold1/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5414 VGND acc0.A\[31\] _0708_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5415 _0708_/a_68_297# net60 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5416 _0340_ _0708_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5417 VPWR acc0.A\[31\] _0708_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X5418 _0340_ _0708_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X5419 _0708_/a_150_297# net60 _0708_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5422 VPWR _0256_ _0639_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5423 VGND _0256_ _0271_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5424 _0639_/a_109_297# _0270_ _0271_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5425 _0271_ _0270_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5426 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5427 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5428 net66 _0990_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5429 _0990_/a_891_413# _0990_/a_193_47# _0990_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5430 _0990_/a_561_413# _0990_/a_27_47# _0990_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5431 VPWR net76 _0990_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5432 net66 _0990_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5433 _0990_/a_381_47# _0088_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5434 VGND _0990_/a_634_159# _0990_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5435 VPWR _0990_/a_891_413# _0990_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5436 _0990_/a_466_413# _0990_/a_193_47# _0990_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5437 VPWR _0990_/a_634_159# _0990_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5438 _0990_/a_634_159# _0990_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5439 _0990_/a_634_159# _0990_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5440 _0990_/a_975_413# _0990_/a_193_47# _0990_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5441 VGND _0990_/a_1059_315# _0990_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5442 _0990_/a_193_47# _0990_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5443 _0990_/a_891_413# _0990_/a_27_47# _0990_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5444 _0990_/a_592_47# _0990_/a_193_47# _0990_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5445 VPWR _0990_/a_1059_315# _0990_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5446 _0990_/a_1017_47# _0990_/a_27_47# _0990_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5447 _0990_/a_193_47# _0990_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5448 _0990_/a_466_413# _0990_/a_27_47# _0990_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5449 VGND _0990_/a_891_413# _0990_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5450 _0990_/a_381_47# _0088_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5451 VGND net76 _0990_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5456 net118 clknet_1_1__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5457 VGND clknet_1_1__leaf__0463_ net118 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5458 net118 clknet_1_1__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5459 VPWR clknet_1_1__leaf__0463_ net118 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5460 VPWR _0161_ _0973_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X5461 _0973_/a_27_297# _0487_ _0973_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X5462 VGND _0161_ _0973_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X5463 _0165_ _0973_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5464 _0973_/a_27_297# _0487_ _0973_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X5465 _0973_/a_109_297# net240 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5466 _0973_/a_373_47# net240 _0973_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5467 _0165_ _0973_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5468 _0973_/a_109_297# _0369_ _0973_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5469 _0973_/a_109_47# _0369_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5472 VPWR comp0.B\[2\] _0956_/a_304_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5473 _0956_/a_304_297# comp0.B\[1\] _0956_/a_220_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5474 VGND comp0.B\[0\] _0956_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.4225 ps=3.9 w=0.65 l=0.15
X5475 _0956_/a_220_297# comp0.B\[0\] _0956_/a_114_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.38 ps=2.76 w=1 l=0.15
X5476 _0956_/a_32_297# comp0.B\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5477 _0956_/a_32_297# comp0.B\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5478 VPWR _0956_/a_32_297# _0475_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.54 ps=5.08 w=1 l=0.15
X5479 _0475_ _0956_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5480 VGND comp0.B\[2\] _0956_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5481 VPWR _0956_/a_32_297# _0475_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5482 _0475_ _0956_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X5483 _0475_ _0956_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5484 _0475_ _0956_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5485 _0956_/a_114_297# comp0.B\[15\] _0956_/a_32_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5486 VGND _0956_/a_32_297# _0475_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5487 VGND _0956_/a_32_297# _0475_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5492 VPWR _0283_ _0421_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5493 _0421_ _0283_ _0810_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5494 _0810_/a_113_47# _0420_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5495 _0421_ _0420_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5496 VPWR input13/a_75_212# net13 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5497 input13/a_75_212# A[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5498 input13/a_75_212# A[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5499 VGND input13/a_75_212# net13 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5500 VPWR input24/a_75_212# net24 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5501 input24/a_75_212# B[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5502 input24/a_75_212# B[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5503 VGND input24/a_75_212# net24 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5504 VPWR clknet_0__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X5505 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X5506 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5507 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5508 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5509 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5510 clkbuf_1_0__f__0464_/a_110_47# clknet_0__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5511 clkbuf_1_0__f__0464_/a_110_47# clknet_0__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X5512 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X5513 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5514 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5515 clkbuf_1_0__f__0464_/a_110_47# clknet_0__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5516 VGND clknet_0__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5517 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5518 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5519 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5520 VGND clknet_0__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5521 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5522 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5523 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5524 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5525 clkbuf_1_0__f__0464_/a_110_47# clknet_0__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5526 VPWR clknet_0__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5527 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5528 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5529 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5530 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5531 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5532 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5533 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5534 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5535 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5536 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5537 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5538 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5539 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5540 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5541 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5542 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5543 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5544 VPWR _0315_ _0741_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5545 VGND _0315_ _0367_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5546 _0741_/a_109_297# _0366_ _0367_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5547 _0367_ _0366_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5548 VGND _0280_ _0672_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X5549 _0672_/a_510_47# _0301_ _0672_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X5550 _0672_/a_79_21# _0303_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X5551 VPWR _0301_ _0672_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5552 _0672_/a_79_21# _0296_ _0672_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X5553 _0672_/a_297_297# _0280_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5554 _0672_/a_79_21# _0303_ _0672_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X5555 VPWR _0672_/a_79_21# _0304_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5556 VGND _0672_/a_79_21# _0304_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5557 _0672_/a_215_47# _0296_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5560 _0655_/a_109_93# _0286_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5561 _0655_/a_215_53# _0283_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.74 as=0 ps=0 w=0.42 l=0.15
X5562 VGND _0655_/a_109_93# _0655_/a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5563 VGND _0280_ _0655_/a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5564 VPWR _0280_ _0655_/a_369_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1365 ps=1.49 w=0.42 l=0.15
X5565 _0655_/a_369_297# _0283_ _0655_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X5566 _0287_ _0655_/a_215_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0 ps=0 w=1 l=0.15
X5567 _0655_/a_297_297# _0655_/a_109_93# _0655_/a_215_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5568 _0655_/a_109_93# _0286_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5569 _0287_ _0655_/a_215_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X5570 VPWR _0586_/a_27_47# _0218_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5571 _0218_ _0586_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5572 VPWR control0.add _0586_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5573 _0218_ _0586_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X5574 VGND _0586_/a_27_47# _0218_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5575 VGND control0.add _0586_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5576 _0724_/a_199_47# _0221_ _0354_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X5577 _0724_/a_113_297# _0333_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X5578 _0354_ _0353_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5579 VPWR _0221_ _0724_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5580 _0724_/a_113_297# _0353_ _0354_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X5581 VGND _0333_ _0724_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5584 control0.count\[0\] _1069_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5585 _1069_/a_891_413# _1069_/a_193_47# _1069_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5586 _1069_/a_561_413# _1069_/a_27_47# _1069_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5587 VPWR clknet_1_0__leaf_clk _1069_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5588 control0.count\[0\] _1069_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5589 _1069_/a_381_47# _0167_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5590 VGND _1069_/a_634_159# _1069_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5591 VPWR _1069_/a_891_413# _1069_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5592 _1069_/a_466_413# _1069_/a_193_47# _1069_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5593 VPWR _1069_/a_634_159# _1069_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5594 _1069_/a_634_159# _1069_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5595 _1069_/a_634_159# _1069_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5596 _1069_/a_975_413# _1069_/a_193_47# _1069_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5597 VGND _1069_/a_1059_315# _1069_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5598 _1069_/a_193_47# _1069_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5599 _1069_/a_891_413# _1069_/a_27_47# _1069_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5600 _1069_/a_592_47# _1069_/a_193_47# _1069_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5601 VPWR _1069_/a_1059_315# _1069_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5602 _1069_/a_1017_47# _1069_/a_27_47# _1069_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5603 _1069_/a_193_47# _1069_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5604 _1069_/a_466_413# _1069_/a_27_47# _1069_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5605 VGND _1069_/a_891_413# _1069_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5606 _1069_/a_381_47# _0167_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5607 VGND clknet_1_0__leaf_clk _1069_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5608 VPWR acc0.A\[0\] hold2/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5609 VGND hold2/a_285_47# hold2/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5610 net149 hold2/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5611 VGND acc0.A\[0\] hold2/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5612 VPWR hold2/a_285_47# hold2/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5613 hold2/a_285_47# hold2/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X5614 hold2/a_285_47# hold2/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X5615 net149 hold2/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5616 _0707_/a_75_199# _0338_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.38025 pd=3.77 as=0 ps=0 w=0.65 l=0.15
X5617 _0707_/a_208_47# _0334_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=2.07 as=0 ps=0 w=0.65 l=0.15
X5618 _0707_/a_315_47# _0333_ _0707_/a_208_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=2.34 as=0 ps=0 w=0.65 l=0.15
X5619 VGND _0335_ _0707_/a_75_199# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5620 _0707_/a_75_199# _0221_ _0707_/a_315_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5621 _0707_/a_75_199# _0338_ _0707_/a_544_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.415 ps=2.83 w=1 l=0.15
X5622 _0707_/a_544_297# _0335_ _0707_/a_201_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.655 ps=5.31 w=1 l=0.15
X5623 VPWR _0707_/a_75_199# _0339_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.285 ps=2.57 w=1 l=0.15
X5624 _0707_/a_201_297# _0334_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5625 VPWR _0333_ _0707_/a_201_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5626 _0707_/a_201_297# _0221_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5627 VGND _0707_/a_75_199# _0339_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5628 VPWR _0216_ _0569_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X5629 _0569_/a_27_297# _0195_ _0569_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X5630 VGND _0216_ _0569_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X5631 _0127_ _0569_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5632 _0569_/a_27_297# _0195_ _0569_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X5633 _0569_/a_109_297# acc0.A\[29\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5634 _0569_/a_373_47# acc0.A\[29\] _0569_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5635 _0127_ _0569_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5636 _0569_/a_109_297# net190 _0569_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5637 _0569_/a_109_47# net190 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5638 VPWR acc0.A\[4\] _0638_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5639 VGND acc0.A\[4\] _0270_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5640 _0638_/a_109_297# net62 _0270_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5641 _0270_ net62 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5644 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5645 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5650 _0972_/a_93_21# control0.state\[1\] _0972_/a_346_47# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X5651 _0972_/a_93_21# _0487_ _0972_/a_250_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X5652 _0972_/a_584_47# _0487_ _0972_/a_93_21# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X5653 VPWR _0972_/a_93_21# _0164_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X5654 VGND net231 _0972_/a_584_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5655 _0972_/a_256_47# _0468_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.16737 ps=1.165 w=0.65 l=0.15
X5656 _0972_/a_250_297# net231 _0972_/a_93_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5657 VGND _0972_/a_93_21# _0164_ VGND sky130_fd_pr__nfet_01v8 ad=0.16737 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X5658 _0972_/a_250_297# _0468_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X5659 VPWR _0471_ _0972_/a_250_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X5660 _0972_/a_250_297# control0.state\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X5661 _0972_/a_346_47# _0471_ _0972_/a_256_47# VGND sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X5662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5666 VPWR comp0.B\[6\] _0955_/a_304_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5667 _0955_/a_304_297# comp0.B\[5\] _0955_/a_220_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5668 VGND comp0.B\[4\] _0955_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.4225 ps=3.9 w=0.65 l=0.15
X5669 _0955_/a_220_297# comp0.B\[4\] _0955_/a_114_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.38 ps=2.76 w=1 l=0.15
X5670 _0955_/a_32_297# comp0.B\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5671 _0955_/a_32_297# comp0.B\[5\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5672 VPWR _0955_/a_32_297# _0474_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.54 ps=5.08 w=1 l=0.15
X5673 _0474_ _0955_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5674 VGND comp0.B\[6\] _0955_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5675 VPWR _0955_/a_32_297# _0474_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5676 _0474_ _0955_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X5677 _0474_ _0955_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5678 _0474_ _0955_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5679 _0955_/a_114_297# comp0.B\[3\] _0955_/a_32_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5680 VGND _0955_/a_32_297# _0474_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5681 VGND _0955_/a_32_297# _0474_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5682 VPWR _0324_ _0366_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5683 _0366_ _0324_ _0740_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5684 _0740_/a_113_47# _0359_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5685 _0366_ _0359_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5686 VPWR input14/a_75_212# net14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5687 input14/a_75_212# A[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5688 input14/a_75_212# A[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5689 VGND input14/a_75_212# net14 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5690 VPWR input25/a_75_212# net25 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5691 input25/a_75_212# B[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5692 input25/a_75_212# B[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5693 VGND input25/a_75_212# net25 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5694 VPWR clknet_0__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X5695 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X5696 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5697 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5698 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5699 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5700 clkbuf_1_0__f__0463_/a_110_47# clknet_0__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5701 clkbuf_1_0__f__0463_/a_110_47# clknet_0__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X5702 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X5703 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5704 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5705 clkbuf_1_0__f__0463_/a_110_47# clknet_0__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5706 VGND clknet_0__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5707 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5708 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5709 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5710 VGND clknet_0__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5711 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5712 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5713 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5714 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5715 clkbuf_1_0__f__0463_/a_110_47# clknet_0__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5716 VPWR clknet_0__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5717 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5718 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5719 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5720 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5721 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5722 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5723 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5724 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5725 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5726 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5727 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5728 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5729 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5730 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5731 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5732 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5733 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5734 _0671_/a_199_47# acc0.A\[15\] _0303_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X5735 _0671_/a_113_297# net42 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X5736 _0303_ _0302_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5737 VPWR acc0.A\[15\] _0671_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5738 _0671_/a_113_297# _0302_ _0303_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X5739 VGND net42 _0671_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5740 VPWR clknet_1_0__leaf__0457_ _0869_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5741 _0459_ _0869_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5742 _0459_ _0869_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5743 VGND clknet_1_0__leaf__0457_ _0869_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5744 net91 clknet_1_0__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5745 VGND clknet_1_0__leaf__0460_ net91 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5746 net91 clknet_1_0__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5747 VPWR clknet_1_0__leaf__0460_ net91 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5748 VPWR _0334_ _0723_/a_207_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1218 ps=1.42 w=0.42 l=0.15
X5749 _0353_ _0723_/a_207_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5750 _0723_/a_297_47# _0723_/a_27_413# _0723_/a_207_413# VGND sky130_fd_pr__nfet_01v8 ad=0.1008 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5751 _0353_ _0723_/a_207_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5752 _0723_/a_207_413# _0723_/a_27_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5753 VPWR _0335_ _0723_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5754 VGND _0334_ _0723_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5755 _0723_/a_27_413# _0335_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5758 VPWR _0285_ _0654_/a_207_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1218 ps=1.42 w=0.42 l=0.15
X5759 _0286_ _0654_/a_207_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5760 _0654_/a_297_47# _0654_/a_27_413# _0654_/a_207_413# VGND sky130_fd_pr__nfet_01v8 ad=0.1008 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5761 _0286_ _0654_/a_207_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5762 _0654_/a_207_413# _0654_/a_27_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5763 VPWR _0284_ _0654_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5764 VGND _0285_ _0654_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5765 _0654_/a_27_413# _0284_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5766 VPWR net1 _0585_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X5767 _0585_/a_27_297# _0216_ _0585_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X5768 VGND net1 _0585_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X5769 _0112_ _0585_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5770 _0585_/a_27_297# _0216_ _0585_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X5771 _0585_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5772 _0585_/a_373_47# _0181_ _0585_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5773 _0112_ _0585_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5774 _0585_/a_109_297# net149 _0585_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5775 _0585_/a_109_47# net149 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5776 net35 _1068_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5777 _1068_/a_891_413# _1068_/a_193_47# _1068_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5778 _1068_/a_561_413# _1068_/a_27_47# _1068_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5779 VPWR clknet_1_0__leaf_clk _1068_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5780 net35 _1068_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5781 _1068_/a_381_47# _0166_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5782 VGND _1068_/a_634_159# _1068_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5783 VPWR _1068_/a_891_413# _1068_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5784 _1068_/a_466_413# _1068_/a_193_47# _1068_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5785 VPWR _1068_/a_634_159# _1068_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5786 _1068_/a_634_159# _1068_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5787 _1068_/a_634_159# _1068_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5788 _1068_/a_975_413# _1068_/a_193_47# _1068_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5789 VGND _1068_/a_1059_315# _1068_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5790 _1068_/a_193_47# _1068_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5791 _1068_/a_891_413# _1068_/a_27_47# _1068_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5792 _1068_/a_592_47# _1068_/a_193_47# _1068_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5793 VPWR _1068_/a_1059_315# _1068_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5794 _1068_/a_1017_47# _1068_/a_27_47# _1068_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5795 _1068_/a_193_47# _1068_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5796 _1068_/a_466_413# _1068_/a_27_47# _1068_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5797 VGND _1068_/a_891_413# _1068_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5798 _1068_/a_381_47# _0166_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5799 VGND clknet_1_0__leaf_clk _1068_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5800 VPWR acc0.A\[21\] hold3/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5801 VGND hold3/a_285_47# hold3/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5802 net150 hold3/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5803 VGND acc0.A\[21\] hold3/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5804 VPWR hold3/a_285_47# hold3/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5805 hold3/a_285_47# hold3/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X5806 hold3/a_285_47# hold3/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X5807 net150 hold3/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5808 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5810 _0338_ _0337_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5811 VGND _0337_ _0338_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5812 _0338_ _0337_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5813 VPWR _0337_ _0338_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5814 _0637_/a_56_297# _0263_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X5815 VPWR _0267_ _0637_/a_56_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5816 _0269_ _0261_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.35425 pd=3.69 as=0 ps=0 w=0.65 l=0.15
X5817 _0637_/a_139_47# _0267_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X5818 _0637_/a_311_297# _0268_ _0637_/a_56_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X5819 _0269_ _0261_ _0637_/a_311_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0 ps=0 w=1 l=0.15
X5820 VGND _0268_ _0269_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5821 _0269_ _0263_ _0637_/a_139_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5822 VPWR _0216_ _0568_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X5823 _0568_/a_27_297# _0195_ _0568_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X5824 VGND _0216_ _0568_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X5825 _0128_ _0568_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5826 _0568_/a_27_297# _0195_ _0568_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X5827 _0568_/a_109_297# net208 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5828 _0568_/a_373_47# net208 _0568_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5829 _0128_ _0568_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5830 _0568_/a_109_297# acc0.A\[29\] _0568_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5831 _0568_/a_109_47# acc0.A\[29\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5832 VPWR control0.sh _0499_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5833 _0178_ _0499_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X5834 VGND control0.sh _0499_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5835 _0499_/a_59_75# _0171_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5836 _0178_ _0499_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X5837 _0499_/a_145_75# _0171_ _0499_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X5838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5839 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5845 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5846 _0971_/a_81_21# _0467_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X5847 _0971_/a_299_297# _0467_ _0971_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X5848 VPWR _0971_/a_81_21# _0163_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5849 VPWR _0181_ _0971_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5850 VGND _0971_/a_81_21# _0163_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5851 VGND _0487_ _0971_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X5852 _0971_/a_299_297# _0487_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5853 _0971_/a_384_47# _0181_ _0971_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5856 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5857 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5858 VPWR comp0.B\[14\] _0954_/a_304_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5859 _0954_/a_304_297# comp0.B\[13\] _0954_/a_220_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5860 VGND comp0.B\[12\] _0954_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.4225 ps=3.9 w=0.65 l=0.15
X5861 _0954_/a_220_297# comp0.B\[12\] _0954_/a_114_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.38 ps=2.76 w=1 l=0.15
X5862 _0954_/a_32_297# comp0.B\[11\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5863 _0954_/a_32_297# comp0.B\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5864 VPWR _0954_/a_32_297# _0473_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.54 ps=5.08 w=1 l=0.15
X5865 _0473_ _0954_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5866 VGND comp0.B\[14\] _0954_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5867 VPWR _0954_/a_32_297# _0473_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5868 _0473_ _0954_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X5869 _0473_ _0954_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5870 _0473_ _0954_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5871 _0954_/a_114_297# comp0.B\[11\] _0954_/a_32_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5872 VGND _0954_/a_32_297# _0473_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5873 VGND _0954_/a_32_297# _0473_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5874 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5875 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5876 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5877 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5878 VPWR input15/a_75_212# net15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5879 input15/a_75_212# A[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5880 input15/a_75_212# A[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5881 VGND input15/a_75_212# net15 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5882 VPWR input26/a_75_212# net26 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5883 input26/a_75_212# B[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5884 input26/a_75_212# B[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5885 VGND input26/a_75_212# net26 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5886 VPWR clknet_0__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X5887 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X5888 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5889 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5890 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5891 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5892 clkbuf_1_0__f__0462_/a_110_47# clknet_0__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5893 clkbuf_1_0__f__0462_/a_110_47# clknet_0__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X5894 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X5895 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5896 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5897 clkbuf_1_0__f__0462_/a_110_47# clknet_0__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5898 VGND clknet_0__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5899 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5900 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5901 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5902 VGND clknet_0__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5903 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5904 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5905 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5906 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5907 clkbuf_1_0__f__0462_/a_110_47# clknet_0__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5908 VPWR clknet_0__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5909 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5910 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5911 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5912 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5913 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5914 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5915 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5916 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5917 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5918 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5919 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5920 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5921 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5922 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5923 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5924 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5925 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5926 VGND acc0.A\[15\] _0670_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X5927 _0670_/a_510_47# net41 _0670_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X5928 _0670_/a_79_21# acc0.A\[14\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X5929 VPWR net41 _0670_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5930 _0670_/a_79_21# net42 _0670_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X5931 _0670_/a_297_297# acc0.A\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5932 _0670_/a_79_21# acc0.A\[14\] _0670_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X5933 VPWR _0670_/a_79_21# _0302_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5934 VGND _0670_/a_79_21# _0302_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5935 _0670_/a_215_47# net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5936 VPWR _0799_/a_80_21# _0413_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X5937 _0799_/a_209_297# _0404_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.65 pd=5.3 as=0 ps=0 w=1 l=0.15
X5938 _0799_/a_303_47# _0298_ _0799_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.208 ps=1.94 w=0.65 l=0.15
X5939 _0799_/a_209_47# _0404_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5940 VGND _0799_/a_80_21# _0413_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X5941 VGND _0343_ _0799_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X5942 _0799_/a_80_21# _0411_ _0799_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5943 VPWR _0298_ _0799_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5944 _0799_/a_80_21# _0343_ _0799_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0 ps=0 w=1 l=0.15
X5945 _0799_/a_209_297# _0411_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5946 VPWR acc0.A\[11\] _0285_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5947 _0285_ acc0.A\[11\] _0653_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5948 _0653_/a_113_47# net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5949 _0285_ net38 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5950 VGND _0347_ _0722_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X5951 _0722_/a_510_47# _0351_ _0722_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X5952 _0722_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X5953 VPWR _0351_ _0722_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5954 _0722_/a_79_21# _0349_ _0722_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X5955 _0722_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5956 _0722_/a_79_21# _0352_ _0722_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X5957 VPWR _0722_/a_79_21# _0110_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5958 VGND _0722_/a_79_21# _0110_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5959 _0722_/a_215_47# _0349_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5960 VPWR net23 _0584_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X5961 _0584_/a_27_297# _0216_ _0584_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X5962 VGND net23 _0584_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X5963 _0113_ _0584_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5964 _0584_/a_27_297# _0216_ _0584_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X5965 _0584_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5966 _0584_/a_373_47# _0181_ _0584_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5967 _0113_ _0584_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5968 _0584_/a_109_297# net157 _0584_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5969 _0584_/a_109_47# net157 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5970 control0.add _1067_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5971 _1067_/a_891_413# _1067_/a_193_47# _1067_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5972 _1067_/a_561_413# _1067_/a_27_47# _1067_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5973 VPWR clknet_1_1__leaf_clk _1067_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5974 control0.add _1067_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5975 _1067_/a_381_47# _0165_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5976 VGND _1067_/a_634_159# _1067_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5977 VPWR _1067_/a_891_413# _1067_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5978 _1067_/a_466_413# _1067_/a_193_47# _1067_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5979 VPWR _1067_/a_634_159# _1067_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5980 _1067_/a_634_159# _1067_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5981 _1067_/a_634_159# _1067_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5982 _1067_/a_975_413# _1067_/a_193_47# _1067_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5983 VGND _1067_/a_1059_315# _1067_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5984 _1067_/a_193_47# _1067_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5985 _1067_/a_891_413# _1067_/a_27_47# _1067_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5986 _1067_/a_592_47# _1067_/a_193_47# _1067_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5987 VPWR _1067_/a_1059_315# _1067_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5988 _1067_/a_1017_47# _1067_/a_27_47# _1067_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5989 _1067_/a_193_47# _1067_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5990 _1067_/a_466_413# _1067_/a_27_47# _1067_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5991 VGND _1067_/a_891_413# _1067_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5992 _1067_/a_381_47# _0165_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5993 VGND clknet_1_1__leaf_clk _1067_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5994 VPWR _0120_ hold4/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5995 VGND hold4/a_285_47# hold4/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5996 net151 hold4/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5997 VGND _0120_ hold4/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5998 VPWR hold4/a_285_47# hold4/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5999 hold4/a_285_47# hold4/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6000 hold4/a_285_47# hold4/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6001 net151 hold4/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6002 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6006 VPWR net61 _0636_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6007 _0268_ _0636_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X6008 VGND net61 _0636_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6009 _0636_/a_59_75# acc0.A\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6010 _0268_ _0636_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6011 _0636_/a_145_75# acc0.A\[3\] _0636_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X6012 VPWR _0336_ _0705_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6013 _0337_ _0705_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X6014 VGND _0336_ _0705_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6015 _0705_/a_59_75# _0220_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6016 _0337_ _0705_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6017 _0705_/a_145_75# _0220_ _0705_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X6018 _0498_/a_240_47# net7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6019 _0159_ _0498_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6020 VGND _0172_ _0498_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6021 _0498_/a_51_297# net247 _0498_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X6022 _0498_/a_149_47# _0177_ _0498_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X6023 _0498_/a_240_47# _0174_ _0498_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6024 VPWR _0172_ _0498_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6025 _0159_ _0498_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X6026 _0498_/a_149_47# net247 _0498_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6027 _0498_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6028 VPWR _0177_ _0498_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6029 _0498_/a_512_297# net7 _0498_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6030 VPWR _0216_ _0567_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X6031 _0567_/a_27_297# _0195_ _0567_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X6032 VGND _0216_ _0567_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X6033 _0129_ _0567_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6034 _0567_/a_27_297# _0195_ _0567_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X6035 _0567_/a_109_297# net162 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6036 _0567_/a_373_47# net162 _0567_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6037 _0129_ _0567_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6038 _0567_/a_109_297# acc0.A\[30\] _0567_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6039 _0567_/a_109_47# acc0.A\[30\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6042 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6044 net129 clknet_1_1__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6045 VGND clknet_1_1__leaf__0464_ net129 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6046 net129 clknet_1_1__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6047 VPWR clknet_1_1__leaf__0464_ net129 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6048 net143 clknet_1_1__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6049 VGND clknet_1_1__leaf__0465_ net143 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6050 net143 clknet_1_1__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6051 VPWR clknet_1_1__leaf__0465_ net143 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6053 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6054 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6055 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6056 VGND acc0.A\[7\] _0619_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6057 _0619_/a_68_297# net65 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6058 _0251_ _0619_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6059 VPWR acc0.A\[7\] _0619_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6060 _0251_ _0619_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6061 _0619_/a_150_297# net65 _0619_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6066 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6068 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6069 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6070 VGND _0484_ _0970_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X6071 VGND _0487_ _0162_ VGND sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X6072 _0162_ _0485_ _0970_/a_114_47# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08937 ps=0.925 w=0.65 l=0.15
X6073 _0970_/a_114_47# _0484_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08937 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X6074 _0970_/a_27_297# _0487_ _0162_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X6075 _0970_/a_27_297# _0485_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6076 _0162_ _0487_ _0970_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6077 VPWR _0484_ _0970_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X6078 _0970_/a_27_297# _0484_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6079 VPWR _0485_ _0970_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X6080 _0970_/a_285_47# _0485_ _0162_ VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X6081 _0162_ _0487_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X6082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6084 net110 clknet_1_0__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6085 VGND clknet_1_0__leaf__0462_ net110 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6086 net110 clknet_1_0__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6087 VPWR clknet_1_0__leaf__0462_ net110 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6088 net124 clknet_1_0__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6089 VGND clknet_1_0__leaf__0463_ net124 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6090 net124 clknet_1_0__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6091 VPWR clknet_1_0__leaf__0463_ net124 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6094 VPWR comp0.B\[10\] _0953_/a_304_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6095 _0953_/a_304_297# comp0.B\[9\] _0953_/a_220_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6096 VGND comp0.B\[8\] _0953_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.4225 ps=3.9 w=0.65 l=0.15
X6097 _0953_/a_220_297# comp0.B\[8\] _0953_/a_114_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.38 ps=2.76 w=1 l=0.15
X6098 _0953_/a_32_297# comp0.B\[7\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6099 _0953_/a_32_297# comp0.B\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6100 VPWR _0953_/a_32_297# _0472_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.54 ps=5.08 w=1 l=0.15
X6101 _0472_ _0953_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6102 VGND comp0.B\[10\] _0953_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6103 VPWR _0953_/a_32_297# _0472_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6104 _0472_ _0953_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6105 _0472_ _0953_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6106 _0472_ _0953_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6107 _0953_/a_114_297# comp0.B\[7\] _0953_/a_32_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6108 VGND _0953_/a_32_297# _0472_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6109 VGND _0953_/a_32_297# _0472_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6112 VPWR input16/a_75_212# net16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6113 input16/a_75_212# A[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6114 input16/a_75_212# A[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6115 VGND input16/a_75_212# net16 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6116 VPWR input27/a_75_212# net27 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6117 input27/a_75_212# B[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6118 input27/a_75_212# B[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6119 VGND input27/a_75_212# net27 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6120 VPWR clknet_0__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X6121 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X6122 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6123 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6124 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6125 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6126 clkbuf_1_0__f__0461_/a_110_47# clknet_0__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6127 clkbuf_1_0__f__0461_/a_110_47# clknet_0__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X6128 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X6129 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6130 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6131 clkbuf_1_0__f__0461_/a_110_47# clknet_0__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6132 VGND clknet_0__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6133 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6134 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6135 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6136 VGND clknet_0__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6137 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6138 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6139 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6140 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6141 clkbuf_1_0__f__0461_/a_110_47# clknet_0__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6142 VPWR clknet_0__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6143 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6144 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6145 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6146 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6147 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6148 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6149 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6150 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6151 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6152 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6153 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6154 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6155 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6156 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6157 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6158 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6159 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6160 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6161 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6162 _0798_/a_199_47# _0298_ _0412_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X6163 _0798_/a_113_297# _0404_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X6164 _0412_ _0411_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6165 VPWR _0298_ _0798_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6166 _0798_/a_113_297# _0411_ _0412_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X6167 VGND _0404_ _0798_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6168 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6172 VPWR _0208_ _0721_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X6173 VGND _0721_/a_27_47# _0352_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X6174 VGND _0721_/a_27_47# _0352_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6175 _0352_ _0721_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X6176 _0352_ _0721_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6177 VGND _0208_ _0721_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X6178 VPWR _0721_/a_27_47# _0352_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6179 _0352_ _0721_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6180 _0352_ _0721_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6181 VPWR _0721_/a_27_47# _0352_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6182 VPWR _0183_ _0583_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X6183 _0583_/a_27_297# _0217_ _0583_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X6184 VGND _0183_ _0583_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X6185 _0114_ _0583_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6186 _0583_/a_27_297# _0217_ _0583_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X6187 _0583_/a_109_297# acc0.A\[16\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6188 _0583_/a_373_47# acc0.A\[16\] _0583_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6189 _0114_ _0583_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6190 _0583_/a_109_297# net165 _0583_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6191 _0583_/a_109_47# net165 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6192 VPWR acc0.A\[11\] _0652_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6193 VGND acc0.A\[11\] _0284_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6194 _0652_/a_109_297# net38 _0284_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6195 _0284_ net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6198 control0.sh _1066_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6199 _1066_/a_891_413# _1066_/a_193_47# _1066_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6200 _1066_/a_561_413# _1066_/a_27_47# _1066_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6201 VPWR clknet_1_1__leaf_clk _1066_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6202 control0.sh _1066_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6203 _1066_/a_381_47# net232 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6204 VGND _1066_/a_634_159# _1066_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6205 VPWR _1066_/a_891_413# _1066_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6206 _1066_/a_466_413# _1066_/a_193_47# _1066_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6207 VPWR _1066_/a_634_159# _1066_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6208 _1066_/a_634_159# _1066_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6209 _1066_/a_634_159# _1066_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6210 _1066_/a_975_413# _1066_/a_193_47# _1066_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6211 VGND _1066_/a_1059_315# _1066_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6212 _1066_/a_193_47# _1066_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6213 _1066_/a_891_413# _1066_/a_27_47# _1066_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6214 _1066_/a_592_47# _1066_/a_193_47# _1066_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6215 VPWR _1066_/a_1059_315# _1066_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6216 _1066_/a_1017_47# _1066_/a_27_47# _1066_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6217 _1066_/a_193_47# _1066_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6218 _1066_/a_466_413# _1066_/a_27_47# _1066_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6219 VGND _1066_/a_891_413# _1066_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6220 _1066_/a_381_47# net232 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6221 VGND clknet_1_1__leaf_clk _1066_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6222 VPWR comp0.B\[10\] hold5/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6223 VGND hold5/a_285_47# hold5/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6224 net152 hold5/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6225 VGND comp0.B\[10\] hold5/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6226 VPWR hold5/a_285_47# hold5/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6227 hold5/a_285_47# hold5/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6228 hold5/a_285_47# hold5/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6229 net152 hold5/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6230 VPWR _0182_ _0566_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X6231 VGND _0566_/a_27_47# _0216_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X6232 VGND _0566_/a_27_47# _0216_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6233 _0216_ _0566_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X6234 _0216_ _0566_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6235 VGND _0182_ _0566_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X6236 VPWR _0566_/a_27_47# _0216_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6237 _0216_ _0566_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6238 _0216_ _0566_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6239 VPWR _0566_/a_27_47# _0216_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6240 _0267_ _0265_ _0635_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X6241 VPWR _0266_ _0267_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X6242 _0635_/a_27_47# _0265_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X6243 _0267_ _0266_ _0635_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6244 _0635_/a_109_297# _0264_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6245 VGND _0264_ _0635_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6246 VGND acc0.A\[30\] _0704_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6247 _0704_/a_68_297# net59 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6248 _0336_ _0704_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6249 VPWR acc0.A\[30\] _0704_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6250 _0336_ _0704_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6251 _0704_/a_150_297# net59 _0704_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6254 VGND acc0.A\[15\] _0497_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6255 _0497_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6256 _0177_ _0497_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6257 VPWR acc0.A\[15\] _0497_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6258 _0177_ _0497_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6259 _0497_/a_150_297# _0176_ _0497_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6260 acc0.A\[3\] _1049_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6261 _1049_/a_891_413# _1049_/a_193_47# _1049_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6262 _1049_/a_561_413# _1049_/a_27_47# _1049_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6263 VPWR net135 _1049_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6264 acc0.A\[3\] _1049_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6265 _1049_/a_381_47# _0147_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6266 VGND _1049_/a_634_159# _1049_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6267 VPWR _1049_/a_891_413# _1049_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6268 _1049_/a_466_413# _1049_/a_193_47# _1049_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6269 VPWR _1049_/a_634_159# _1049_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6270 _1049_/a_634_159# _1049_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6271 _1049_/a_634_159# _1049_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6272 _1049_/a_975_413# _1049_/a_193_47# _1049_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6273 VGND _1049_/a_1059_315# _1049_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6274 _1049_/a_193_47# _1049_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6275 _1049_/a_891_413# _1049_/a_27_47# _1049_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6276 _1049_/a_592_47# _1049_/a_193_47# _1049_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6277 VPWR _1049_/a_1059_315# _1049_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6278 _1049_/a_1017_47# _1049_/a_27_47# _1049_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6279 _1049_/a_193_47# _1049_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6280 _1049_/a_466_413# _1049_/a_27_47# _1049_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6281 VGND _1049_/a_891_413# _1049_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6282 _1049_/a_381_47# _0147_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6283 VGND net135 _1049_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6286 VGND _0222_ _0618_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X6287 _0618_/a_510_47# _0232_ _0618_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X6288 _0618_/a_79_21# _0249_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X6289 VPWR _0232_ _0618_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6290 _0618_/a_79_21# _0223_ _0618_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X6291 _0618_/a_297_297# _0222_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6292 _0618_/a_79_21# _0249_ _0618_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X6293 VPWR _0618_/a_79_21# _0250_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6294 VGND _0618_/a_79_21# _0250_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6295 _0618_/a_215_47# _0223_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6296 VGND net171 _0549_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6297 _0549_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6298 _0207_ _0549_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6299 VPWR net171 _0549_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6300 _0207_ _0549_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6301 _0549_/a_150_297# _0176_ _0549_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6314 _0471_ control0.state\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6315 VGND control0.state\[0\] _0471_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6316 _0471_ control0.state\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6317 VPWR control0.state\[0\] _0471_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6320 net102 clknet_1_1__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6321 VGND clknet_1_1__leaf__0461_ net102 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6322 net102 clknet_1_1__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6323 VPWR clknet_1_1__leaf__0461_ net102 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6324 VPWR input17/a_75_212# net17 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6325 input17/a_75_212# B[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6326 input17/a_75_212# B[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6327 VGND input17/a_75_212# net17 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6328 VPWR input28/a_75_212# net28 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6329 input28/a_75_212# B[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6330 input28/a_75_212# B[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6331 VGND input28/a_75_212# net28 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6332 VPWR clknet_0__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X6333 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X6334 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6335 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6336 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6337 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6338 clkbuf_1_0__f__0460_/a_110_47# clknet_0__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6339 clkbuf_1_0__f__0460_/a_110_47# clknet_0__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X6340 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X6341 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6342 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6343 clkbuf_1_0__f__0460_/a_110_47# clknet_0__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6344 VGND clknet_0__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6345 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6346 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6347 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6348 VGND clknet_0__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6349 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6350 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6351 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6352 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6353 clkbuf_1_0__f__0460_/a_110_47# clknet_0__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6354 VPWR clknet_0__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6355 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6356 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6357 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6358 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6359 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6360 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6361 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6362 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6363 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6364 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6365 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6366 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6367 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6368 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6369 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6370 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6371 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6372 VPWR clknet_1_1__leaf__0457_ _0935_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6373 _0465_ _0935_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6374 _0465_ _0935_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6375 VGND clknet_1_1__leaf__0457_ _0935_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6378 VPWR _0299_ _0797_/a_207_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1218 ps=1.42 w=0.42 l=0.15
X6379 _0411_ _0797_/a_207_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6380 _0797_/a_297_47# _0797_/a_27_413# _0797_/a_207_413# VGND sky130_fd_pr__nfet_01v8 ad=0.1008 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X6381 _0411_ _0797_/a_207_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6382 _0797_/a_207_413# _0797_/a_27_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6383 VPWR _0297_ _0797_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6384 VGND _0299_ _0797_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6385 _0797_/a_27_413# _0297_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6388 VGND _0350_ _0720_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6389 _0720_/a_68_297# net239 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6390 _0351_ _0720_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6391 VPWR _0350_ _0720_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6392 _0351_ _0720_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6393 _0720_/a_150_297# net239 _0720_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6396 VPWR _0281_ _0283_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6397 _0283_ _0281_ _0651_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X6398 _0651_/a_113_47# _0282_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6399 _0283_ _0282_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6400 VPWR _0183_ _0582_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X6401 _0582_/a_27_297# _0217_ _0582_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X6402 VGND _0183_ _0582_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X6403 _0115_ _0582_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6404 _0582_/a_27_297# _0217_ _0582_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X6405 _0582_/a_109_297# net219 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6406 _0582_/a_373_47# net219 _0582_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6407 _0115_ _0582_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6408 _0582_/a_109_297# net221 _0582_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6409 _0582_/a_109_47# net221 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6410 net83 clknet_1_1__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6411 VGND clknet_1_1__leaf__0459_ net83 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6412 net83 clknet_1_1__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6413 VPWR clknet_1_1__leaf__0459_ net83 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6414 control0.reset _1065_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6415 _1065_/a_891_413# _1065_/a_193_47# _1065_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6416 _1065_/a_561_413# _1065_/a_27_47# _1065_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6417 VPWR clknet_1_1__leaf_clk _1065_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6418 control0.reset _1065_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6419 _1065_/a_381_47# _0163_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6420 VGND _1065_/a_634_159# _1065_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6421 VPWR _1065_/a_891_413# _1065_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6422 _1065_/a_466_413# _1065_/a_193_47# _1065_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6423 VPWR _1065_/a_634_159# _1065_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6424 _1065_/a_634_159# _1065_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6425 _1065_/a_634_159# _1065_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6426 _1065_/a_975_413# _1065_/a_193_47# _1065_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6427 VGND _1065_/a_1059_315# _1065_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6428 _1065_/a_193_47# _1065_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6429 _1065_/a_891_413# _1065_/a_27_47# _1065_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6430 _1065_/a_592_47# _1065_/a_193_47# _1065_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6431 VPWR _1065_/a_1059_315# _1065_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6432 _1065_/a_1017_47# _1065_/a_27_47# _1065_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6433 _1065_/a_193_47# _1065_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6434 _1065_/a_466_413# _1065_/a_27_47# _1065_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6435 VGND _1065_/a_891_413# _1065_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6436 _1065_/a_381_47# _0163_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6437 VGND clknet_1_1__leaf_clk _1065_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6438 VGND _0219_ _0849_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X6439 _0849_/a_510_47# _0451_ _0849_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X6440 _0849_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X6441 VPWR _0451_ _0849_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6442 _0849_/a_79_21# net222 _0849_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X6443 _0849_/a_297_297# _0219_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6444 _0849_/a_79_21# _0399_ _0849_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X6445 VPWR _0849_/a_79_21# _0082_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6446 VGND _0849_/a_79_21# _0082_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6447 _0849_/a_215_47# net222 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6448 VPWR _0139_ hold6/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6449 VGND hold6/a_285_47# hold6/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6450 net153 hold6/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6451 VGND _0139_ hold6/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6452 VPWR hold6/a_285_47# hold6/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6453 hold6/a_285_47# hold6/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6454 hold6/a_285_47# hold6/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6455 net153 hold6/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6456 VPWR acc0.A\[29\] _0703_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6457 VGND acc0.A\[29\] _0335_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6458 _0703_/a_109_297# net57 _0335_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6459 _0335_ net57 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6460 VPWR _0175_ _0496_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X6461 VPWR _0496_/a_27_47# _0176_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6462 VGND _0175_ _0496_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X6463 _0176_ _0496_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X6464 _0176_ _0496_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X6465 VGND _0496_/a_27_47# _0176_ VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6466 _0565_/a_240_47# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6467 _0130_ _0565_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6468 VGND _0208_ _0565_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6469 _0565_/a_51_297# net201 _0565_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X6470 _0565_/a_149_47# _0215_ _0565_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X6471 _0565_/a_240_47# _0173_ _0565_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6472 VPWR _0208_ _0565_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6473 _0130_ _0565_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X6474 _0565_/a_149_47# net201 _0565_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6475 _0565_/a_245_297# _0173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6476 VPWR _0215_ _0565_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6477 _0565_/a_512_297# net17 _0565_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6478 VPWR acc0.A\[1\] _0266_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6479 _0266_ acc0.A\[1\] _0634_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X6480 _0634_/a_113_47# net47 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6481 _0266_ net47 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6484 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6492 acc0.A\[2\] _1048_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6493 _1048_/a_891_413# _1048_/a_193_47# _1048_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6494 _1048_/a_561_413# _1048_/a_27_47# _1048_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6495 VPWR net134 _1048_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6496 acc0.A\[2\] _1048_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6497 _1048_/a_381_47# _0146_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6498 VGND _1048_/a_634_159# _1048_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6499 VPWR _1048_/a_891_413# _1048_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6500 _1048_/a_466_413# _1048_/a_193_47# _1048_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6501 VPWR _1048_/a_634_159# _1048_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6502 _1048_/a_634_159# _1048_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6503 _1048_/a_634_159# _1048_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6504 _1048_/a_975_413# _1048_/a_193_47# _1048_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6505 VGND _1048_/a_1059_315# _1048_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6506 _1048_/a_193_47# _1048_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6507 _1048_/a_891_413# _1048_/a_27_47# _1048_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6508 _1048_/a_592_47# _1048_/a_193_47# _1048_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6509 VPWR _1048_/a_1059_315# _1048_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6510 _1048_/a_1017_47# _1048_/a_27_47# _1048_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6511 _1048_/a_193_47# _1048_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6512 _1048_/a_466_413# _1048_/a_27_47# _1048_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6513 VGND _1048_/a_891_413# _1048_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6514 _1048_/a_381_47# _0146_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6515 VGND net134 _1048_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6516 VPWR clknet_0_clk clkbuf_1_1__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X6517 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X6518 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6519 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6520 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6521 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6522 clkbuf_1_1__f_clk/a_110_47# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6523 clkbuf_1_1__f_clk/a_110_47# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X6524 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X6525 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6526 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6527 clkbuf_1_1__f_clk/a_110_47# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6528 VGND clknet_0_clk clkbuf_1_1__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6529 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6530 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6531 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6532 VGND clknet_0_clk clkbuf_1_1__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6533 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6534 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6535 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6536 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6537 clkbuf_1_1__f_clk/a_110_47# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6538 VPWR clknet_0_clk clkbuf_1_1__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6539 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6540 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6541 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6542 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6543 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6544 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6545 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6546 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6547 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6548 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6549 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6550 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6551 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6552 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6553 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6554 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6555 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6556 _0548_/a_240_47# net31 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6557 _0138_ _0548_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6558 VGND _0172_ _0548_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6559 _0548_/a_51_297# net173 _0548_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X6560 _0548_/a_149_47# _0206_ _0548_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X6561 _0548_/a_240_47# _0174_ _0548_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6562 VPWR _0172_ _0548_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6563 _0138_ _0548_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X6564 _0548_/a_149_47# net173 _0548_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6565 _0548_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6566 VPWR _0206_ _0548_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6567 _0548_/a_512_297# net31 _0548_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6568 VGND _0238_ _0617_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6569 _0617_/a_68_297# _0248_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6570 _0249_ _0617_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6571 VPWR _0238_ _0617_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6572 _0249_ _0617_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6573 _0617_/a_150_297# _0248_ _0617_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6578 net69 clknet_1_0__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6579 VGND clknet_1_0__leaf__0458_ net69 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6580 net69 clknet_1_0__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6581 VPWR clknet_1_0__leaf__0458_ net69 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6584 _0951_/a_109_93# control0.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6585 _0470_ _0951_/a_209_311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X6586 _0951_/a_109_93# control0.state\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6587 _0951_/a_296_53# _0951_/a_109_93# _0951_/a_209_311# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.10783 ps=1.36 w=0.42 l=0.15
X6588 VPWR comp0.B\[0\] _0951_/a_209_311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.07438 ps=0.815 w=0.42 l=0.15
X6589 _0951_/a_368_53# _0161_ _0951_/a_296_53# VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6590 _0470_ _0951_/a_209_311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12228 ps=1.08 w=0.65 l=0.15
X6591 _0951_/a_209_311# _0161_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07438 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X6592 VPWR _0951_/a_109_93# _0951_/a_209_311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X6593 VGND comp0.B\[0\] _0951_/a_368_53# VGND sky130_fd_pr__nfet_01v8 ad=0.12228 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X6594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6596 VPWR input18/a_75_212# net18 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6597 input18/a_75_212# B[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6598 input18/a_75_212# B[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6599 VGND input18/a_75_212# net18 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6600 VPWR input29/a_75_212# net29 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6601 input29/a_75_212# B[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6602 input29/a_75_212# B[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6603 VGND input29/a_75_212# net29 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6604 VGND _0369_ _0796_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X6605 _0796_/a_510_47# _0410_ _0796_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X6606 _0796_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X6607 VPWR _0410_ _0796_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6608 _0796_/a_79_21# net238 _0796_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X6609 _0796_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6610 _0796_/a_79_21# _0399_ _0796_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X6611 VPWR _0796_/a_79_21# _0094_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6612 VGND _0796_/a_79_21# _0094_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6613 _0796_/a_215_47# net238 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6616 VPWR _0183_ _0581_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X6617 _0581_/a_27_297# _0217_ _0581_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X6618 VGND _0183_ _0581_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X6619 _0116_ _0581_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6620 _0581_/a_27_297# _0217_ _0581_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X6621 _0581_/a_109_297# net206 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6622 _0581_/a_373_47# net206 _0581_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6623 _0116_ _0581_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6624 _0581_/a_109_297# net219 _0581_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6625 _0581_/a_109_47# net219 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6626 VGND acc0.A\[10\] _0650_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6627 _0650_/a_68_297# net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6628 _0282_ _0650_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6629 VPWR acc0.A\[10\] _0650_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6630 _0282_ _0650_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6631 _0650_/a_150_297# net37 _0650_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6632 control0.state\[2\] _1064_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6633 _1064_/a_891_413# _1064_/a_193_47# _1064_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6634 _1064_/a_561_413# _1064_/a_27_47# _1064_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6635 VPWR clknet_1_0__leaf_clk _1064_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6636 control0.state\[2\] _1064_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6637 _1064_/a_381_47# _0162_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6638 VGND _1064_/a_634_159# _1064_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6639 VPWR _1064_/a_891_413# _1064_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6640 _1064_/a_466_413# _1064_/a_193_47# _1064_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6641 VPWR _1064_/a_634_159# _1064_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6642 _1064_/a_634_159# _1064_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6643 _1064_/a_634_159# _1064_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6644 _1064_/a_975_413# _1064_/a_193_47# _1064_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6645 VGND _1064_/a_1059_315# _1064_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6646 _1064_/a_193_47# _1064_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6647 _1064_/a_891_413# _1064_/a_27_47# _1064_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6648 _1064_/a_592_47# _1064_/a_193_47# _1064_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6649 VPWR _1064_/a_1059_315# _1064_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6650 _1064_/a_1017_47# _1064_/a_27_47# _1064_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6651 _1064_/a_193_47# _1064_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6652 _1064_/a_466_413# _1064_/a_27_47# _1064_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6653 VGND _1064_/a_891_413# _1064_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6654 _1064_/a_381_47# _0162_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6655 VGND clknet_1_0__leaf_clk _1064_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6658 net140 clknet_1_0__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6659 VGND clknet_1_0__leaf__0465_ net140 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6660 net140 clknet_1_0__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6661 VPWR clknet_1_0__leaf__0465_ net140 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6662 _0451_ _0450_ _0848_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X6663 VPWR _0350_ _0451_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X6664 _0848_/a_27_47# _0450_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X6665 _0451_ _0350_ _0848_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6666 _0848_/a_109_297# _0446_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6667 VGND _0446_ _0848_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6668 VGND _0347_ _0779_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X6669 _0779_/a_510_47# _0396_ _0779_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X6670 _0779_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X6671 VPWR _0396_ _0779_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6672 _0779_/a_79_21# _0395_ _0779_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X6673 _0779_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6674 _0779_/a_79_21# _0352_ _0779_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X6675 VPWR _0779_/a_79_21# _0097_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6676 VGND _0779_/a_79_21# _0097_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6677 _0779_/a_215_47# _0395_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6678 VPWR acc0.A\[4\] hold7/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6679 VGND hold7/a_285_47# hold7/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6680 net154 hold7/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6681 VGND acc0.A\[4\] hold7/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6682 VPWR hold7/a_285_47# hold7/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6683 hold7/a_285_47# hold7/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6684 hold7/a_285_47# hold7/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6685 net154 hold7/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6686 VPWR acc0.A\[29\] _0334_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6687 _0334_ acc0.A\[29\] _0702_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X6688 _0702_/a_113_47# net57 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6689 _0334_ net57 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6694 VPWR acc0.A\[1\] _0633_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6695 VGND acc0.A\[1\] _0265_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6696 _0633_/a_109_297# net47 _0265_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6697 _0265_ net47 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6698 VGND control0.reset _0495_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6699 _0495_/a_68_297# control0.sh VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6700 _0175_ _0495_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6701 VPWR control0.reset _0495_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6702 _0175_ _0495_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6703 _0495_/a_150_297# control0.sh _0495_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6704 VGND comp0.B\[0\] _0564_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6705 _0564_/a_68_297# _0175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6706 _0215_ _0564_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6707 VPWR comp0.B\[0\] _0564_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6708 _0215_ _0564_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6709 _0564_/a_150_297# _0175_ _0564_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6710 acc0.A\[1\] _1047_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6711 _1047_/a_891_413# _1047_/a_193_47# _1047_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6712 _1047_/a_561_413# _1047_/a_27_47# _1047_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6713 VPWR net133 _1047_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6714 acc0.A\[1\] _1047_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6715 _1047_/a_381_47# _0145_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6716 VGND _1047_/a_634_159# _1047_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6717 VPWR _1047_/a_891_413# _1047_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6718 _1047_/a_466_413# _1047_/a_193_47# _1047_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6719 VPWR _1047_/a_634_159# _1047_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6720 _1047_/a_634_159# _1047_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6721 _1047_/a_634_159# _1047_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6722 _1047_/a_975_413# _1047_/a_193_47# _1047_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6723 VGND _1047_/a_1059_315# _1047_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6724 _1047_/a_193_47# _1047_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6725 _1047_/a_891_413# _1047_/a_27_47# _1047_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6726 _1047_/a_592_47# _1047_/a_193_47# _1047_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6727 VPWR _1047_/a_1059_315# _1047_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6728 _1047_/a_1017_47# _1047_/a_27_47# _1047_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6729 _1047_/a_193_47# _1047_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6730 _1047_/a_466_413# _1047_/a_27_47# _1047_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6731 VGND _1047_/a_891_413# _1047_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6732 _1047_/a_381_47# _0145_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6733 VGND net133 _1047_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6737 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6738 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6740 net121 clknet_1_1__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6741 VGND clknet_1_1__leaf__0463_ net121 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6742 net121 clknet_1_1__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6743 VPWR clknet_1_1__leaf__0463_ net121 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6744 net135 clknet_1_0__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6745 VGND clknet_1_0__leaf__0464_ net135 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6746 net135 clknet_1_0__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6747 VPWR clknet_1_0__leaf__0464_ net135 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6750 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6751 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6752 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6753 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6754 _0616_/a_78_199# _0247_ _0616_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.5655 ps=5.64 w=0.65 l=0.15
X6755 VPWR _0240_ _0616_/a_493_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6756 _0616_/a_493_297# _0246_ _0616_/a_78_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.47 ps=2.94 w=1 l=0.15
X6757 VPWR _0616_/a_78_199# _0248_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X6758 VGND _0246_ _0616_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6759 _0616_/a_78_199# _0241_ _0616_/a_292_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.235 ps=2.47 w=1 l=0.15
X6760 _0616_/a_215_47# _0240_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6761 _0616_/a_215_47# _0241_ _0616_/a_78_199# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6762 _0616_/a_292_297# _0247_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6763 VGND _0616_/a_78_199# _0248_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6768 VGND comp0.B\[8\] _0547_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6769 _0547_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6770 _0206_ _0547_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6771 VPWR comp0.B\[8\] _0547_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6772 _0206_ _0547_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6773 _0547_/a_150_297# _0176_ _0547_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6778 net116 clknet_1_1__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6779 VGND clknet_1_1__leaf__0462_ net116 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6780 net116 clknet_1_1__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6781 VPWR clknet_1_1__leaf__0462_ net116 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6782 VPWR _0950_/a_75_212# _0161_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6783 _0950_/a_75_212# _0469_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6784 _0950_/a_75_212# _0469_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6785 VGND _0950_/a_75_212# _0161_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6786 VPWR clknet_0__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X6787 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X6788 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6789 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6790 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6791 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6792 clkbuf_1_1__f__0459_/a_110_47# clknet_0__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6793 clkbuf_1_1__f__0459_/a_110_47# clknet_0__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X6794 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X6795 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6796 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6797 clkbuf_1_1__f__0459_/a_110_47# clknet_0__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6798 VGND clknet_0__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6799 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6800 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6801 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6802 VGND clknet_0__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6803 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6804 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6805 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6806 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6807 clkbuf_1_1__f__0459_/a_110_47# clknet_0__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6808 VPWR clknet_0__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6809 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6810 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6811 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6812 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6813 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6814 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6815 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6816 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6817 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6818 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6819 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6820 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6821 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6822 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6823 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6824 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6825 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6828 VPWR input19/a_75_212# net19 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6829 input19/a_75_212# B[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6830 input19/a_75_212# B[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6831 VGND input19/a_75_212# net19 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6834 _0795_/a_81_21# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X6835 _0795_/a_299_297# _0346_ _0795_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X6836 VPWR _0795_/a_81_21# _0410_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6837 VPWR _0405_ _0795_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6838 VGND _0795_/a_81_21# _0410_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6839 VGND _0409_ _0795_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X6840 _0795_/a_299_297# _0409_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6841 _0795_/a_384_47# _0405_ _0795_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6844 VPWR _0183_ _0580_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X6845 _0580_/a_27_297# _0217_ _0580_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X6846 VGND _0183_ _0580_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X6847 _0117_ _0580_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6848 _0580_/a_27_297# _0217_ _0580_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X6849 _0580_/a_109_297# acc0.A\[19\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6850 _0580_/a_373_47# acc0.A\[19\] _0580_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6851 _0117_ _0580_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6852 _0580_/a_109_297# net206 _0580_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6853 _0580_/a_109_47# net206 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6856 control0.state\[1\] _1063_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6857 _1063_/a_891_413# _1063_/a_193_47# _1063_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6858 _1063_/a_561_413# _1063_/a_27_47# _1063_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6859 VPWR clknet_1_1__leaf_clk _1063_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6860 control0.state\[1\] _1063_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6861 _1063_/a_381_47# _0161_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6862 VGND _1063_/a_634_159# _1063_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6863 VPWR _1063_/a_891_413# _1063_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6864 _1063_/a_466_413# _1063_/a_193_47# _1063_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6865 VPWR _1063_/a_634_159# _1063_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6866 _1063_/a_634_159# _1063_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6867 _1063_/a_634_159# _1063_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6868 _1063_/a_975_413# _1063_/a_193_47# _1063_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6869 VGND _1063_/a_1059_315# _1063_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6870 _1063_/a_193_47# _1063_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6871 _1063_/a_891_413# _1063_/a_27_47# _1063_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6872 _1063_/a_592_47# _1063_/a_193_47# _1063_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6873 VPWR _1063_/a_1059_315# _1063_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6874 _1063_/a_1017_47# _1063_/a_27_47# _1063_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6875 _1063_/a_193_47# _1063_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6876 _1063_/a_466_413# _1063_/a_27_47# _1063_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6877 VGND _1063_/a_891_413# _1063_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6878 _1063_/a_381_47# _0161_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6879 VGND clknet_1_1__leaf_clk _1063_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6882 VGND _0218_ _0778_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6883 _0778_/a_68_297# net44 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6884 _0396_ _0778_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6885 VPWR _0218_ _0778_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6886 _0396_ _0778_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6887 _0778_/a_150_297# net44 _0778_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6888 VPWR _0263_ _0847_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6889 VGND _0263_ _0450_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6890 _0847_/a_109_297# _0267_ _0450_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6891 _0450_ _0267_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6894 VPWR acc0.A\[26\] hold8/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6895 VGND hold8/a_285_47# hold8/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6896 net155 hold8/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6897 VGND acc0.A\[26\] hold8/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6898 VPWR hold8/a_285_47# hold8/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6899 hold8/a_285_47# hold8/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6900 hold8/a_285_47# hold8/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6901 net155 hold8/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6904 VPWR _0701_/a_80_21# _0333_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X6905 _0701_/a_209_297# _0330_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.65 pd=5.3 as=0 ps=0 w=1 l=0.15
X6906 _0701_/a_303_47# _0329_ _0701_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.208 ps=1.94 w=0.65 l=0.15
X6907 _0701_/a_209_47# _0330_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6908 VGND _0701_/a_80_21# _0333_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X6909 VGND _0332_ _0701_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X6910 _0701_/a_80_21# _0327_ _0701_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6911 VPWR _0329_ _0701_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6912 _0701_/a_80_21# _0332_ _0701_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0 ps=0 w=1 l=0.15
X6913 _0701_/a_209_297# _0327_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6914 _0563_/a_240_47# net24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6915 _0131_ _0563_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6916 VGND _0208_ _0563_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6917 _0563_/a_51_297# net203 _0563_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X6918 _0563_/a_149_47# _0214_ _0563_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X6919 _0563_/a_240_47# _0173_ _0563_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6920 VPWR _0208_ _0563_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6921 _0131_ _0563_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X6922 _0563_/a_149_47# net203 _0563_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6923 _0563_/a_245_297# _0173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6924 VPWR _0214_ _0563_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6925 _0563_/a_512_297# net24 _0563_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6926 VPWR net149 _0264_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6927 _0264_ net149 _0632_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X6928 _0632_/a_113_47# net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6929 _0264_ net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6932 VPWR _0494_/a_27_47# _0174_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6933 _0174_ _0494_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6934 VPWR _0173_ _0494_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6935 _0174_ _0494_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X6936 VGND _0494_/a_27_47# _0174_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6937 VGND _0173_ _0494_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6938 comp0.B\[14\] _1046_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6939 _1046_/a_891_413# _1046_/a_193_47# _1046_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6940 _1046_/a_561_413# _1046_/a_27_47# _1046_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6941 VPWR net132 _1046_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6942 comp0.B\[14\] _1046_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6943 _1046_/a_381_47# net158 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6944 VGND _1046_/a_634_159# _1046_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6945 VPWR _1046_/a_891_413# _1046_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6946 _1046_/a_466_413# _1046_/a_193_47# _1046_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6947 VPWR _1046_/a_634_159# _1046_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6948 _1046_/a_634_159# _1046_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6949 _1046_/a_634_159# _1046_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6950 _1046_/a_975_413# _1046_/a_193_47# _1046_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6951 VGND _1046_/a_1059_315# _1046_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6952 _1046_/a_193_47# _1046_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6953 _1046_/a_891_413# _1046_/a_27_47# _1046_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6954 _1046_/a_592_47# _1046_/a_193_47# _1046_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6955 VPWR _1046_/a_1059_315# _1046_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6956 _1046_/a_1017_47# _1046_/a_27_47# _1046_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6957 _1046_/a_193_47# _1046_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6958 _1046_/a_466_413# _1046_/a_27_47# _1046_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6959 VGND _1046_/a_891_413# _1046_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6960 _1046_/a_381_47# net158 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6961 VGND net132 _1046_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6968 _0546_/a_240_47# net32 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6969 _0139_ _0546_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6970 VGND _0172_ _0546_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6971 _0546_/a_51_297# net152 _0546_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X6972 _0546_/a_149_47# _0205_ _0546_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X6973 _0546_/a_240_47# _0174_ _0546_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6974 VPWR _0172_ _0546_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6975 _0139_ _0546_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X6976 _0546_/a_149_47# net152 _0546_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6977 _0546_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6978 VPWR _0205_ _0546_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6979 _0546_/a_512_297# net32 _0546_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6980 VPWR _0242_ _0615_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6981 VGND _0242_ _0247_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6982 _0615_/a_109_297# _0244_ _0247_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6983 _0247_ _0244_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6984 acc0.A\[29\] _1029_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6985 _1029_/a_891_413# _1029_/a_193_47# _1029_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6986 _1029_/a_561_413# _1029_/a_27_47# _1029_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6987 VPWR net115 _1029_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6988 acc0.A\[29\] _1029_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6989 _1029_/a_381_47# net191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6990 VGND _1029_/a_634_159# _1029_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6991 VPWR _1029_/a_891_413# _1029_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6992 _1029_/a_466_413# _1029_/a_193_47# _1029_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6993 VPWR _1029_/a_634_159# _1029_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6994 _1029_/a_634_159# _1029_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6995 _1029_/a_634_159# _1029_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6996 _1029_/a_975_413# _1029_/a_193_47# _1029_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6997 VGND _1029_/a_1059_315# _1029_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6998 _1029_/a_193_47# _1029_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6999 _1029_/a_891_413# _1029_/a_27_47# _1029_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7000 _1029_/a_592_47# _1029_/a_193_47# _1029_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7001 VPWR _1029_/a_1059_315# _1029_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7002 _1029_/a_1017_47# _1029_/a_27_47# _1029_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7003 _1029_/a_193_47# _1029_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7004 _1029_/a_466_413# _1029_/a_27_47# _1029_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7005 VGND _1029_/a_891_413# _1029_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7006 _1029_/a_381_47# net191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7007 VGND net115 _1029_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7008 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7009 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7010 VPWR net10 _0529_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X7011 _0529_/a_27_297# _0186_ _0529_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X7012 VGND net10 _0529_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X7013 _0197_ _0529_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7014 _0529_/a_27_297# _0186_ _0529_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X7015 _0529_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7016 _0529_/a_373_47# _0180_ _0529_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7017 _0197_ _0529_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7018 _0529_/a_109_297# net170 _0529_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7019 _0529_/a_109_47# net170 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7020 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7021 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7022 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7023 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7024 VPWR clknet_1_0__leaf__0457_ _0880_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X7025 _0460_ _0880_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X7026 _0460_ _0880_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X7027 VGND clknet_1_0__leaf__0457_ _0880_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X7028 VPWR clknet_0__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X7029 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X7030 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7031 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7032 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7033 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7034 clkbuf_1_1__f__0458_/a_110_47# clknet_0__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7035 clkbuf_1_1__f__0458_/a_110_47# clknet_0__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X7036 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X7037 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7038 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7039 clkbuf_1_1__f__0458_/a_110_47# clknet_0__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7040 VGND clknet_0__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7041 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7042 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7043 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7044 VGND clknet_0__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7045 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7046 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7047 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7048 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7049 clkbuf_1_1__f__0458_/a_110_47# clknet_0__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7050 VPWR clknet_0__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7051 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7052 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7053 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7054 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7055 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7056 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7057 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7058 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7059 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7060 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7061 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7062 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7063 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7064 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7065 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7066 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7067 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7068 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7069 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7070 net94 clknet_1_1__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7071 VGND clknet_1_1__leaf__0460_ net94 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7072 net94 clknet_1_1__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7073 VPWR clknet_1_1__leaf__0460_ net94 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7074 _0794_/a_110_297# _0297_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X7075 VGND _0297_ _0794_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.17225 ps=1.83 w=0.65 l=0.15
X7076 _0409_ _0404_ _0794_/a_110_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X7077 VPWR _0300_ _0409_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X7078 _0794_/a_27_47# _0404_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X7079 _0794_/a_326_47# _0300_ _0794_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.12675 ps=1.04 w=0.65 l=0.15
X7080 _0409_ _0277_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X7081 _0409_ _0277_ _0794_/a_326_47# VGND sky130_fd_pr__nfet_01v8 ad=0.39325 pd=2.51 as=0.06825 ps=0.86 w=0.65 l=0.15
X7082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7088 control0.state\[0\] _1062_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7089 _1062_/a_891_413# _1062_/a_193_47# _1062_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7090 _1062_/a_561_413# _1062_/a_27_47# _1062_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7091 VPWR clknet_1_1__leaf_clk _1062_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7092 control0.state\[0\] _1062_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7093 _1062_/a_381_47# _0160_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7094 VGND _1062_/a_634_159# _1062_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7095 VPWR _1062_/a_891_413# _1062_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7096 _1062_/a_466_413# _1062_/a_193_47# _1062_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7097 VPWR _1062_/a_634_159# _1062_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7098 _1062_/a_634_159# _1062_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7099 _1062_/a_634_159# _1062_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7100 _1062_/a_975_413# _1062_/a_193_47# _1062_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7101 VGND _1062_/a_1059_315# _1062_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7102 _1062_/a_193_47# _1062_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7103 _1062_/a_891_413# _1062_/a_27_47# _1062_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7104 _1062_/a_592_47# _1062_/a_193_47# _1062_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7105 VPWR _1062_/a_1059_315# _1062_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7106 _1062_/a_1017_47# _1062_/a_27_47# _1062_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7107 _1062_/a_193_47# _1062_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7108 _1062_/a_466_413# _1062_/a_27_47# _1062_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7109 VGND _1062_/a_891_413# _1062_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7110 _1062_/a_381_47# _0160_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7111 VGND clknet_1_1__leaf_clk _1062_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7112 _0846_/a_240_47# net233 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X7113 _0083_ _0846_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7114 VGND _0219_ _0846_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7115 _0846_/a_51_297# _0449_ _0846_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X7116 _0846_/a_149_47# _0345_ _0846_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X7117 _0846_/a_240_47# _0448_ _0846_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7118 VPWR _0219_ _0846_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7119 _0083_ _0846_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X7120 _0846_/a_149_47# _0449_ _0846_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7121 _0846_/a_245_297# _0448_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7122 VPWR _0345_ _0846_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7123 _0846_/a_512_297# net233 _0846_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7124 _0777_/a_377_297# _0309_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X7125 _0777_/a_47_47# _0394_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7126 _0777_/a_129_47# _0394_ _0777_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X7127 _0777_/a_285_47# _0394_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X7128 _0395_ _0777_/a_47_47# _0777_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X7129 VGND _0309_ _0777_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7130 VPWR _0309_ _0777_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7131 VPWR _0777_/a_47_47# _0395_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X7132 _0395_ _0394_ _0777_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7133 _0777_/a_285_47# _0309_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7134 VPWR _0125_ hold9/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7135 VGND hold9/a_285_47# hold9/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7136 net156 hold9/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7137 VGND _0125_ hold9/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7138 VPWR hold9/a_285_47# hold9/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7139 hold9/a_285_47# hold9/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7140 hold9/a_285_47# hold9/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7141 net156 hold9/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7142 VPWR _0221_ _0332_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7143 _0332_ _0221_ _0700_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X7144 _0700_/a_113_47# _0331_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7145 _0332_ _0331_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7146 VPWR _0261_ _0631_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7147 VGND _0261_ _0263_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7148 _0631_/a_109_297# _0262_ _0263_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7149 _0263_ _0262_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7150 VGND net201 _0562_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7151 _0562_/a_68_297# _0175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7152 _0214_ _0562_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7153 VPWR net201 _0562_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7154 _0214_ _0562_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7155 _0562_/a_150_297# _0175_ _0562_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7156 VPWR _0171_ _0173_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7157 _0173_ _0171_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7158 VPWR control0.sh _0173_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7159 _0493_/a_27_47# control0.sh VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7160 _0493_/a_27_47# _0171_ _0173_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7161 _0173_ _0171_ _0493_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7162 _0173_ control0.sh VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7163 VGND control0.sh _0493_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7164 comp0.B\[13\] _1045_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7165 _1045_/a_891_413# _1045_/a_193_47# _1045_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7166 _1045_/a_561_413# _1045_/a_27_47# _1045_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7167 VPWR net131 _1045_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7168 comp0.B\[13\] _1045_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7169 _1045_/a_381_47# net184 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7170 VGND _1045_/a_634_159# _1045_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7171 VPWR _1045_/a_891_413# _1045_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7172 _1045_/a_466_413# _1045_/a_193_47# _1045_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7173 VPWR _1045_/a_634_159# _1045_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7174 _1045_/a_634_159# _1045_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7175 _1045_/a_634_159# _1045_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7176 _1045_/a_975_413# _1045_/a_193_47# _1045_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7177 VGND _1045_/a_1059_315# _1045_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7178 _1045_/a_193_47# _1045_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7179 _1045_/a_891_413# _1045_/a_27_47# _1045_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7180 _1045_/a_592_47# _1045_/a_193_47# _1045_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7181 VPWR _1045_/a_1059_315# _1045_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7182 _1045_/a_1017_47# _1045_/a_27_47# _1045_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7183 _1045_/a_193_47# _1045_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7184 _1045_/a_466_413# _1045_/a_27_47# _1045_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7185 VGND _1045_/a_891_413# _1045_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7186 _1045_/a_381_47# net184 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7187 VGND net131 _1045_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7188 _0437_ _0435_ _0829_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X7189 VPWR _0436_ _0437_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X7190 _0829_/a_27_47# _0435_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X7191 _0437_ _0436_ _0829_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7192 _0829_/a_109_297# _0429_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7193 VGND _0429_ _0829_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7194 _0246_ _0614_/a_29_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X7195 _0614_/a_111_297# _0245_ _0614_/a_29_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.26 as=0.1092 ps=1.36 w=0.42 l=0.15
X7196 _0246_ _0614_/a_29_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7197 _0614_/a_183_297# _0244_ _0614_/a_111_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1386 pd=1.5 as=0 ps=0 w=0.42 l=0.15
X7198 VPWR _0243_ _0614_/a_183_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7199 _0614_/a_29_53# _0244_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.74 as=0 ps=0 w=0.42 l=0.15
X7200 VGND _0245_ _0614_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7201 VGND _0243_ _0614_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7206 VGND comp0.B\[9\] _0545_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7207 _0545_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7208 _0205_ _0545_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7209 VPWR comp0.B\[9\] _0545_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7210 _0205_ _0545_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7211 _0545_/a_150_297# _0176_ _0545_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7212 acc0.A\[28\] _1028_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7213 _1028_/a_891_413# _1028_/a_193_47# _1028_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7214 _1028_/a_561_413# _1028_/a_27_47# _1028_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7215 VPWR net114 _1028_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7216 acc0.A\[28\] _1028_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7217 _1028_/a_381_47# _0126_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7218 VGND _1028_/a_634_159# _1028_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7219 VPWR _1028_/a_891_413# _1028_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7220 _1028_/a_466_413# _1028_/a_193_47# _1028_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7221 VPWR _1028_/a_634_159# _1028_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7222 _1028_/a_634_159# _1028_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7223 _1028_/a_634_159# _1028_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7224 _1028_/a_975_413# _1028_/a_193_47# _1028_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7225 VGND _1028_/a_1059_315# _1028_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7226 _1028_/a_193_47# _1028_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7227 _1028_/a_891_413# _1028_/a_27_47# _1028_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7228 _1028_/a_592_47# _1028_/a_193_47# _1028_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7229 VPWR _1028_/a_1059_315# _1028_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7230 _1028_/a_1017_47# _1028_/a_27_47# _1028_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7231 _1028_/a_193_47# _1028_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7232 _1028_/a_466_413# _1028_/a_27_47# _1028_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7233 VGND _1028_/a_891_413# _1028_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7234 _1028_/a_381_47# _0126_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7235 VGND net114 _1028_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X7241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X7242 _0528_/a_81_21# _0196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X7243 _0528_/a_299_297# _0196_ _0528_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X7244 VPWR _0528_/a_81_21# _0148_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7245 VPWR net170 _0528_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7246 VGND _0528_/a_81_21# _0148_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7247 VGND _0195_ _0528_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X7248 _0528_/a_299_297# _0195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7249 _0528_/a_384_47# net170 _0528_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7250 VPWR clknet_0__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X7251 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X7252 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7253 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7254 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7255 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7256 clkbuf_1_1__f__0457_/a_110_47# clknet_0__0457_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7257 clkbuf_1_1__f__0457_/a_110_47# clknet_0__0457_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X7258 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X7259 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7260 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7261 clkbuf_1_1__f__0457_/a_110_47# clknet_0__0457_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7262 VGND clknet_0__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7263 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7264 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7265 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7266 VGND clknet_0__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7267 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7268 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7269 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7270 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7271 clkbuf_1_1__f__0457_/a_110_47# clknet_0__0457_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7272 VPWR clknet_0__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7273 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7274 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7275 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7276 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7277 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7278 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7279 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7280 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7281 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7282 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7283 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7284 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7285 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7286 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7287 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7288 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7289 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7290 net107 clknet_1_0__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7291 VGND clknet_1_0__leaf__0461_ net107 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7292 net107 clknet_1_0__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7293 VPWR clknet_1_0__leaf__0461_ net107 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7294 _0793_/a_240_47# net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X7295 _0095_ _0793_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7296 VGND _0219_ _0793_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7297 _0793_/a_51_297# _0408_ _0793_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X7298 _0793_/a_149_47# _0345_ _0793_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X7299 _0793_/a_240_47# _0407_ _0793_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7300 VPWR _0219_ _0793_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7301 _0095_ _0793_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X7302 _0793_/a_149_47# _0408_ _0793_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7303 _0793_/a_245_297# _0407_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7304 VPWR _0345_ _0793_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7305 _0793_/a_512_297# net42 _0793_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7306 VPWR _0459_ clkbuf_0__0459_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X7307 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X7308 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7309 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7310 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7311 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7312 clkbuf_0__0459_/a_110_47# _0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7313 clkbuf_0__0459_/a_110_47# _0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X7314 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X7315 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7316 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7317 clkbuf_0__0459_/a_110_47# _0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7318 VGND _0459_ clkbuf_0__0459_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7319 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7320 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7321 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7322 VGND _0459_ clkbuf_0__0459_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7323 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7324 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7325 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7326 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7327 clkbuf_0__0459_/a_110_47# _0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7328 VPWR _0459_ clkbuf_0__0459_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7329 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7330 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7331 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7332 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7333 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7334 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7335 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7336 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7337 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7338 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7339 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7340 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7341 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7342 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7343 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7344 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7345 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7346 net98 clknet_1_1__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7347 VGND clknet_1_1__leaf__0461_ net98 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7348 net98 clknet_1_1__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7349 VPWR clknet_1_1__leaf__0461_ net98 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7350 acc0.A\[15\] _1061_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7351 VPWR _1061_/a_1059_315# acc0.A\[15\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7352 _1061_/a_891_413# _1061_/a_193_47# _1061_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7353 _1061_/a_561_413# _1061_/a_27_47# _1061_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7354 VPWR net147 _1061_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7355 acc0.A\[15\] _1061_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7356 _1061_/a_381_47# _0159_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7357 VGND _1061_/a_634_159# _1061_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7358 VGND _1061_/a_1059_315# acc0.A\[15\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7359 VPWR _1061_/a_891_413# _1061_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7360 _1061_/a_466_413# _1061_/a_193_47# _1061_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7361 VPWR _1061_/a_634_159# _1061_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7362 _1061_/a_634_159# _1061_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7363 _1061_/a_634_159# _1061_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X7364 _1061_/a_975_413# _1061_/a_193_47# _1061_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7365 VGND _1061_/a_1059_315# _1061_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7366 _1061_/a_193_47# _1061_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7367 _1061_/a_891_413# _1061_/a_27_47# _1061_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7368 _1061_/a_592_47# _1061_/a_193_47# _1061_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7369 VPWR _1061_/a_1059_315# _1061_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7370 _1061_/a_1017_47# _1061_/a_27_47# _1061_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7371 _1061_/a_193_47# _1061_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7372 _1061_/a_466_413# _1061_/a_27_47# _1061_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7373 VGND _1061_/a_891_413# _1061_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7374 _1061_/a_381_47# _0159_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7375 VGND net147 _1061_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7376 _0449_ _0350_ _0845_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X7377 _0449_ _0447_ _0845_/a_193_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X7378 _0845_/a_193_297# _0446_ _0845_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7379 VGND _0446_ _0845_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7380 VPWR _0350_ _0449_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X7381 _0845_/a_109_47# _0447_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X7382 _0845_/a_109_297# _0261_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7383 _0845_/a_109_47# _0261_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7384 _0394_ _0308_ _0776_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X7385 VPWR _0306_ _0394_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X7386 _0776_/a_27_47# _0308_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X7387 _0394_ _0306_ _0776_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7388 _0776_/a_109_297# _0387_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7389 VGND _0387_ _0776_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7392 net132 clknet_1_1__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7393 VGND clknet_1_1__leaf__0464_ net132 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7394 net132 clknet_1_1__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7395 VPWR clknet_1_1__leaf__0464_ net132 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7396 net146 clknet_1_1__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7397 VGND clknet_1_1__leaf__0465_ net146 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7398 net146 clknet_1_1__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7399 VPWR clknet_1_1__leaf__0465_ net146 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7400 _0561_/a_240_47# net25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X7401 _0132_ _0561_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7402 VGND _0208_ _0561_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7403 _0561_/a_51_297# net185 _0561_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X7404 _0561_/a_149_47# _0213_ _0561_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X7405 _0561_/a_240_47# _0173_ _0561_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7406 VPWR _0208_ _0561_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7407 _0132_ _0561_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X7408 _0561_/a_149_47# net185 _0561_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7409 _0561_/a_245_297# _0173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7410 VPWR _0213_ _0561_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7411 _0561_/a_512_297# net25 _0561_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7412 VPWR _0492_/a_27_47# _0172_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7413 _0172_ _0492_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7414 VPWR _0171_ _0492_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7415 _0172_ _0492_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X7416 VGND _0492_/a_27_47# _0172_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7417 VGND _0171_ _0492_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7418 VPWR acc0.A\[2\] _0630_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7419 VGND acc0.A\[2\] _0262_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7420 _0630_/a_109_297# net58 _0262_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7421 _0262_ net58 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7422 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7423 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7424 comp0.B\[12\] _1044_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7425 _1044_/a_891_413# _1044_/a_193_47# _1044_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7426 _1044_/a_561_413# _1044_/a_27_47# _1044_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7427 VPWR net130 _1044_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7428 comp0.B\[12\] _1044_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7429 _1044_/a_381_47# net194 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7430 VGND _1044_/a_634_159# _1044_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7431 VPWR _1044_/a_891_413# _1044_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7432 _1044_/a_466_413# _1044_/a_193_47# _1044_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7433 VPWR _1044_/a_634_159# _1044_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7434 _1044_/a_634_159# _1044_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7435 _1044_/a_634_159# _1044_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7436 _1044_/a_975_413# _1044_/a_193_47# _1044_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7437 VGND _1044_/a_1059_315# _1044_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7438 _1044_/a_193_47# _1044_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7439 _1044_/a_891_413# _1044_/a_27_47# _1044_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7440 _1044_/a_592_47# _1044_/a_193_47# _1044_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7441 VPWR _1044_/a_1059_315# _1044_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7442 _1044_/a_1017_47# _1044_/a_27_47# _1044_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7443 _1044_/a_193_47# _1044_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7444 _1044_/a_466_413# _1044_/a_27_47# _1044_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7445 VGND _1044_/a_891_413# _1044_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7446 _1044_/a_381_47# net194 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7447 VGND net130 _1044_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7450 net79 clknet_1_1__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7451 VGND clknet_1_1__leaf__0459_ net79 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7452 net79 clknet_1_1__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7453 VPWR clknet_1_1__leaf__0459_ net79 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7454 VPWR _0226_ _0381_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7455 _0381_ _0226_ _0759_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X7456 _0759_/a_113_47# _0373_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7457 _0381_ _0373_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7460 _0828_/a_199_47# _0429_ _0436_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X7461 _0828_/a_113_297# _0435_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X7462 _0436_ _0343_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7463 VPWR _0429_ _0828_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7464 _0828_/a_113_297# _0343_ _0436_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X7465 VGND _0435_ _0828_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7466 net72 clknet_1_1__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7467 VGND clknet_1_1__leaf__0458_ net72 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7468 net72 clknet_1_1__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7469 VPWR clknet_1_1__leaf__0458_ net72 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7476 VPWR acc0.A\[18\] _0613_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7477 VGND acc0.A\[18\] _0245_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7478 _0613_/a_109_297# net45 _0245_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7479 _0245_ net45 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7480 _0544_/a_240_47# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X7481 _0140_ _0544_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7482 VGND _0172_ _0544_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7483 _0544_/a_51_297# net198 _0544_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X7484 _0544_/a_149_47# _0204_ _0544_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X7485 _0544_/a_240_47# _0174_ _0544_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7486 VPWR _0172_ _0544_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7487 _0140_ _0544_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X7488 _0544_/a_149_47# net198 _0544_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7489 _0544_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7490 VPWR _0204_ _0544_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7491 _0544_/a_512_297# net18 _0544_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7492 net113 clknet_1_1__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7493 VGND clknet_1_1__leaf__0462_ net113 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7494 net113 clknet_1_1__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7495 VPWR clknet_1_1__leaf__0462_ net113 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7498 acc0.A\[27\] _1027_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7499 _1027_/a_891_413# _1027_/a_193_47# _1027_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7500 _1027_/a_561_413# _1027_/a_27_47# _1027_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7501 VPWR net113 _1027_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7502 acc0.A\[27\] _1027_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7503 _1027_/a_381_47# net156 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7504 VGND _1027_/a_634_159# _1027_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7505 VPWR _1027_/a_891_413# _1027_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7506 _1027_/a_466_413# _1027_/a_193_47# _1027_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7507 VPWR _1027_/a_634_159# _1027_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7508 _1027_/a_634_159# _1027_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7509 _1027_/a_634_159# _1027_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7510 _1027_/a_975_413# _1027_/a_193_47# _1027_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7511 VGND _1027_/a_1059_315# _1027_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7512 _1027_/a_193_47# _1027_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7513 _1027_/a_891_413# _1027_/a_27_47# _1027_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7514 _1027_/a_592_47# _1027_/a_193_47# _1027_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7515 VPWR _1027_/a_1059_315# _1027_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7516 _1027_/a_1017_47# _1027_/a_27_47# _1027_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7517 _1027_/a_193_47# _1027_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7518 _1027_/a_466_413# _1027_/a_27_47# _1027_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7519 VGND _1027_/a_891_413# _1027_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7520 _1027_/a_381_47# net156 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7521 VGND net113 _1027_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7522 VPWR net53 hold90/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7523 VGND hold90/a_285_47# hold90/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7524 net237 hold90/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7525 VGND net53 hold90/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7526 VPWR hold90/a_285_47# hold90/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7527 hold90/a_285_47# hold90/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7528 hold90/a_285_47# hold90/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7529 net237 hold90/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7530 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7531 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7534 VPWR net11 _0527_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X7535 _0527_/a_27_297# _0186_ _0527_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X7536 VGND net11 _0527_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X7537 _0196_ _0527_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7538 _0527_/a_27_297# _0186_ _0527_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X7539 _0527_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7540 _0527_/a_373_47# _0180_ _0527_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7541 _0196_ _0527_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7542 _0527_/a_109_297# net154 _0527_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7543 _0527_/a_109_47# net154 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7546 VPWR _0792_/a_80_21# _0408_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X7547 _0792_/a_209_297# _0405_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.65 pd=5.3 as=0 ps=0 w=1 l=0.15
X7548 _0792_/a_303_47# _0400_ _0792_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.208 ps=1.94 w=0.65 l=0.15
X7549 _0792_/a_209_47# _0405_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7550 VGND _0792_/a_80_21# _0408_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X7551 VGND _0343_ _0792_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X7552 _0792_/a_80_21# _0406_ _0792_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7553 VPWR _0400_ _0792_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7554 _0792_/a_80_21# _0343_ _0792_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0 ps=0 w=1 l=0.15
X7555 _0792_/a_209_297# _0406_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7557 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7560 VPWR _0458_ clkbuf_0__0458_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X7561 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X7562 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7563 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7564 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7565 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7566 clkbuf_0__0458_/a_110_47# _0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7567 clkbuf_0__0458_/a_110_47# _0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X7568 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X7569 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7570 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7571 clkbuf_0__0458_/a_110_47# _0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7572 VGND _0458_ clkbuf_0__0458_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7573 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7574 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7575 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7576 VGND _0458_ clkbuf_0__0458_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7577 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7578 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7579 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7580 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7581 clkbuf_0__0458_/a_110_47# _0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7582 VPWR _0458_ clkbuf_0__0458_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7583 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7584 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7585 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7586 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7587 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7588 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7589 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7590 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7591 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7592 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7593 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7594 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7595 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7596 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7597 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7598 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7599 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7601 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7604 acc0.A\[14\] _1060_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7605 _1060_/a_891_413# _1060_/a_193_47# _1060_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7606 _1060_/a_561_413# _1060_/a_27_47# _1060_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7607 VPWR net146 _1060_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7608 acc0.A\[14\] _1060_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7609 _1060_/a_381_47# _0158_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7610 VGND _1060_/a_634_159# _1060_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7611 VPWR _1060_/a_891_413# _1060_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7612 _1060_/a_466_413# _1060_/a_193_47# _1060_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7613 VPWR _1060_/a_634_159# _1060_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7614 _1060_/a_634_159# _1060_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7615 _1060_/a_634_159# _1060_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7616 _1060_/a_975_413# _1060_/a_193_47# _1060_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7617 VGND _1060_/a_1059_315# _1060_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7618 _1060_/a_193_47# _1060_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7619 _1060_/a_891_413# _1060_/a_27_47# _1060_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7620 _1060_/a_592_47# _1060_/a_193_47# _1060_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7621 VPWR _1060_/a_1059_315# _1060_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7622 _1060_/a_1017_47# _1060_/a_27_47# _1060_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7623 _1060_/a_193_47# _1060_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7624 _1060_/a_466_413# _1060_/a_27_47# _1060_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7625 VGND _1060_/a_891_413# _1060_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7626 _1060_/a_381_47# _0158_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7627 VGND net146 _1060_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7628 VPWR _0261_ _0844_/a_382_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.305 ps=2.61 w=1 l=0.15
X7629 _0844_/a_297_47# _0447_ _0844_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.3705 pd=3.74 as=0.169 ps=1.82 w=0.65 l=0.15
X7630 _0844_/a_297_47# _0261_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7631 VGND _0446_ _0844_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7632 VPWR _0844_/a_79_21# _0448_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X7633 _0844_/a_79_21# _0447_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.15
X7634 _0844_/a_382_297# _0446_ _0844_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7635 VGND _0844_/a_79_21# _0448_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7636 VPWR clknet_1_1__leaf__0457_ _0913_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X7637 _0463_ _0913_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X7638 _0463_ _0913_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X7639 VGND clknet_1_1__leaf__0457_ _0913_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X7640 VGND _0347_ _0775_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X7641 _0775_/a_510_47# _0393_ _0775_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X7642 _0775_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X7643 VPWR _0393_ _0775_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7644 _0775_/a_79_21# _0392_ _0775_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X7645 _0775_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7646 _0775_/a_79_21# _0352_ _0775_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X7647 VPWR _0775_/a_79_21# _0098_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7648 VGND _0775_/a_79_21# _0098_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7649 _0775_/a_215_47# _0392_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7650 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7652 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7653 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7654 _0171_ control0.reset VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7655 VGND control0.reset _0171_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7656 _0171_ control0.reset VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7657 VPWR control0.reset _0171_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7658 VGND comp0.B\[2\] _0560_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7659 _0560_/a_68_297# _0175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7660 _0213_ _0560_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7661 VPWR comp0.B\[2\] _0560_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7662 _0213_ _0560_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7663 _0560_/a_150_297# _0175_ _0560_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7664 comp0.B\[11\] _1043_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7665 _1043_/a_891_413# _1043_/a_193_47# _1043_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7666 _1043_/a_561_413# _1043_/a_27_47# _1043_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7667 VPWR net129 _1043_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7668 comp0.B\[11\] _1043_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7669 _1043_/a_381_47# net196 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7670 VGND _1043_/a_634_159# _1043_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7671 VPWR _1043_/a_891_413# _1043_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7672 _1043_/a_466_413# _1043_/a_193_47# _1043_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7673 VPWR _1043_/a_634_159# _1043_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7674 _1043_/a_634_159# _1043_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7675 _1043_/a_634_159# _1043_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7676 _1043_/a_975_413# _1043_/a_193_47# _1043_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7677 VGND _1043_/a_1059_315# _1043_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7678 _1043_/a_193_47# _1043_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7679 _1043_/a_891_413# _1043_/a_27_47# _1043_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7680 _1043_/a_592_47# _1043_/a_193_47# _1043_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7681 VPWR _1043_/a_1059_315# _1043_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7682 _1043_/a_1017_47# _1043_/a_27_47# _1043_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7683 _1043_/a_193_47# _1043_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7684 _1043_/a_466_413# _1043_/a_27_47# _1043_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7685 VGND _1043_/a_891_413# _1043_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7686 _1043_/a_381_47# net196 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7687 VGND net129 _1043_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7688 _0435_ _0434_ _0827_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X7689 VPWR _0273_ _0435_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X7690 _0827_/a_27_47# _0434_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X7691 _0435_ _0273_ _0827_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7692 _0827_/a_109_297# _0430_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7693 VGND _0430_ _0827_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7694 VGND _0347_ _0758_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X7695 _0758_/a_510_47# _0380_ _0758_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X7696 _0758_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X7697 VPWR _0380_ _0758_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7698 _0758_/a_79_21# _0379_ _0758_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X7699 _0758_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7700 _0758_/a_79_21# _0352_ _0758_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X7701 VPWR _0758_/a_79_21# _0102_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7702 VGND _0758_/a_79_21# _0102_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7703 _0758_/a_215_47# _0379_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7704 VGND _0319_ _0689_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7705 _0689_/a_68_297# _0320_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7706 _0321_ _0689_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7707 VPWR _0319_ _0689_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7708 _0321_ _0689_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7709 _0689_/a_150_297# _0320_ _0689_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7714 VPWR net45 _0612_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7715 _0244_ _0612_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X7716 VGND net45 _0612_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7717 _0612_/a_59_75# acc0.A\[18\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7718 _0244_ _0612_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7719 _0612_/a_145_75# acc0.A\[18\] _0612_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X7720 VGND net152 _0543_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7721 _0543_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7722 _0204_ _0543_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7723 VPWR net152 _0543_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7724 _0204_ _0543_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7725 _0543_/a_150_297# _0176_ _0543_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7726 acc0.A\[26\] _1026_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7727 _1026_/a_891_413# _1026_/a_193_47# _1026_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7728 _1026_/a_561_413# _1026_/a_27_47# _1026_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7729 VPWR net112 _1026_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7730 acc0.A\[26\] _1026_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7731 _1026_/a_381_47# _0124_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7732 VGND _1026_/a_634_159# _1026_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7733 VPWR _1026_/a_891_413# _1026_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7734 _1026_/a_466_413# _1026_/a_193_47# _1026_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7735 VPWR _1026_/a_634_159# _1026_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7736 _1026_/a_634_159# _1026_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7737 _1026_/a_634_159# _1026_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7738 _1026_/a_975_413# _1026_/a_193_47# _1026_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7739 VGND _1026_/a_1059_315# _1026_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7740 _1026_/a_193_47# _1026_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7741 _1026_/a_891_413# _1026_/a_27_47# _1026_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7742 _1026_/a_592_47# _1026_/a_193_47# _1026_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7743 VPWR _1026_/a_1059_315# _1026_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7744 _1026_/a_1017_47# _1026_/a_27_47# _1026_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7745 _1026_/a_193_47# _1026_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7746 _1026_/a_466_413# _1026_/a_27_47# _1026_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7747 VGND _1026_/a_891_413# _1026_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7748 _1026_/a_381_47# _0124_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7749 VGND net112 _1026_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7750 VPWR net57 hold80/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7751 VGND hold80/a_285_47# hold80/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7752 net227 hold80/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7753 VGND net57 hold80/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7754 VPWR hold80/a_285_47# hold80/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7755 hold80/a_285_47# hold80/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7756 hold80/a_285_47# hold80/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7757 net227 hold80/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7758 VPWR net41 hold91/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7759 VGND hold91/a_285_47# hold91/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7760 net238 hold91/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7761 VGND net41 hold91/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7762 VPWR hold91/a_285_47# hold91/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7763 hold91/a_285_47# hold91/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7764 hold91/a_285_47# hold91/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7765 net238 hold91/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7766 VPWR _0178_ _0526_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X7767 VGND _0526_/a_27_47# _0195_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X7768 VGND _0526_/a_27_47# _0195_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7769 _0195_ _0526_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X7770 _0195_ _0526_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7771 VGND _0178_ _0526_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X7772 VPWR _0526_/a_27_47# _0195_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7773 _0195_ _0526_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7774 _0195_ _0526_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7775 VPWR _0526_/a_27_47# _0195_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7778 net55 _1009_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7779 _1009_/a_891_413# _1009_/a_193_47# _1009_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7780 _1009_/a_561_413# _1009_/a_27_47# _1009_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7781 VPWR net95 _1009_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7782 net55 _1009_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7783 _1009_/a_381_47# _0107_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7784 VGND _1009_/a_634_159# _1009_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7785 VPWR _1009_/a_891_413# _1009_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7786 _1009_/a_466_413# _1009_/a_193_47# _1009_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7787 VPWR _1009_/a_634_159# _1009_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7788 _1009_/a_634_159# _1009_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7789 _1009_/a_634_159# _1009_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7790 _1009_/a_975_413# _1009_/a_193_47# _1009_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7791 VGND _1009_/a_1059_315# _1009_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7792 _1009_/a_193_47# _1009_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7793 _1009_/a_891_413# _1009_/a_27_47# _1009_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7794 _1009_/a_592_47# _1009_/a_193_47# _1009_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7795 VPWR _1009_/a_1059_315# _1009_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7796 _1009_/a_1017_47# _1009_/a_27_47# _1009_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7797 _1009_/a_193_47# _1009_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7798 _1009_/a_466_413# _1009_/a_27_47# _1009_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7799 VGND _1009_/a_891_413# _1009_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7800 _1009_/a_381_47# _0107_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7801 VGND net95 _1009_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7802 net105 clknet_1_0__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7803 VGND clknet_1_0__leaf__0461_ net105 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7804 net105 clknet_1_0__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7805 VPWR clknet_1_0__leaf__0461_ net105 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7808 VPWR _0509_/a_27_47# _0186_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7809 _0186_ _0509_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7810 VPWR _0182_ _0509_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7811 _0186_ _0509_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X7812 VGND _0509_/a_27_47# _0186_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7813 VGND _0182_ _0509_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X7815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X7816 _0791_/a_199_47# _0400_ _0407_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X7817 _0791_/a_113_297# _0405_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X7818 _0407_ _0406_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7819 VPWR _0400_ _0791_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7820 _0791_/a_113_297# _0406_ _0407_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X7821 VGND _0405_ _0791_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7822 net86 clknet_1_0__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7823 VGND clknet_1_0__leaf__0459_ net86 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7824 net86 clknet_1_0__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7825 VPWR clknet_1_0__leaf__0459_ net86 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7826 net65 _0989_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7827 _0989_/a_891_413# _0989_/a_193_47# _0989_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7828 _0989_/a_561_413# _0989_/a_27_47# _0989_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7829 VPWR net75 _0989_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7830 net65 _0989_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7831 _0989_/a_381_47# _0087_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7832 VGND _0989_/a_634_159# _0989_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7833 VPWR _0989_/a_891_413# _0989_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7834 _0989_/a_466_413# _0989_/a_193_47# _0989_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7835 VPWR _0989_/a_634_159# _0989_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7836 _0989_/a_634_159# _0989_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7837 _0989_/a_634_159# _0989_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7838 _0989_/a_975_413# _0989_/a_193_47# _0989_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7839 VGND _0989_/a_1059_315# _0989_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7840 _0989_/a_193_47# _0989_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7841 _0989_/a_891_413# _0989_/a_27_47# _0989_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7842 _0989_/a_592_47# _0989_/a_193_47# _0989_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7843 VPWR _0989_/a_1059_315# _0989_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7844 _0989_/a_1017_47# _0989_/a_27_47# _0989_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7845 _0989_/a_193_47# _0989_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7846 _0989_/a_466_413# _0989_/a_27_47# _0989_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7847 VGND _0989_/a_891_413# _0989_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7848 _0989_/a_381_47# _0087_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7849 VGND net75 _0989_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7850 VPWR _0457_ clkbuf_0__0457_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X7851 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X7852 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7853 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7854 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7855 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7856 clkbuf_0__0457_/a_110_47# _0457_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7857 clkbuf_0__0457_/a_110_47# _0457_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X7858 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X7859 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7860 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7861 clkbuf_0__0457_/a_110_47# _0457_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7862 VGND _0457_ clkbuf_0__0457_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7863 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7864 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7865 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7866 VGND _0457_ clkbuf_0__0457_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7867 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7868 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7869 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7870 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7871 clkbuf_0__0457_/a_110_47# _0457_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7872 VPWR _0457_ clkbuf_0__0457_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7873 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7874 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7875 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7876 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7877 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7878 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7879 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7880 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7881 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7882 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7883 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7884 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7885 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7886 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7887 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7888 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7889 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7894 VGND _0260_ _0843_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7895 _0843_/a_68_297# _0268_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7896 _0447_ _0843_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7897 VPWR _0260_ _0843_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7898 _0447_ _0843_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7899 _0843_/a_150_297# _0268_ _0843_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7900 VGND _0218_ _0774_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7901 _0774_/a_68_297# net45 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7902 _0393_ _0774_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7903 VPWR _0218_ _0774_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7904 _0393_ _0774_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7905 _0774_/a_150_297# net45 _0774_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7908 comp0.B\[10\] _1042_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7909 _1042_/a_891_413# _1042_/a_193_47# _1042_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7910 _1042_/a_561_413# _1042_/a_27_47# _1042_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7911 VPWR net128 _1042_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7912 comp0.B\[10\] _1042_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7913 _1042_/a_381_47# _0140_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7914 VGND _1042_/a_634_159# _1042_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7915 VPWR _1042_/a_891_413# _1042_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7916 _1042_/a_466_413# _1042_/a_193_47# _1042_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7917 VPWR _1042_/a_634_159# _1042_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7918 _1042_/a_634_159# _1042_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7919 _1042_/a_634_159# _1042_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7920 _1042_/a_975_413# _1042_/a_193_47# _1042_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7921 VGND _1042_/a_1059_315# _1042_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7922 _1042_/a_193_47# _1042_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7923 _1042_/a_891_413# _1042_/a_27_47# _1042_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7924 _1042_/a_592_47# _1042_/a_193_47# _1042_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7925 VPWR _1042_/a_1059_315# _1042_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7926 _1042_/a_1017_47# _1042_/a_27_47# _1042_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7927 _1042_/a_193_47# _1042_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7928 _1042_/a_466_413# _1042_/a_27_47# _1042_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7929 VGND _1042_/a_891_413# _1042_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7930 _1042_/a_381_47# _0140_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7931 VGND net128 _1042_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X7933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X7934 _0826_/a_219_297# _0826_/a_27_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X7935 VGND _0433_ _0826_/a_27_53# VGND sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X7936 VPWR _0255_ _0826_/a_301_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X7937 _0434_ _0826_/a_219_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10187 ps=0.99 w=0.65 l=0.15
X7938 _0826_/a_301_297# _0826_/a_27_53# _0826_/a_219_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7939 _0434_ _0826_/a_219_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7940 _0826_/a_27_53# _0433_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7941 VGND _0255_ _0826_/a_219_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7942 VGND _0350_ _0757_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7943 _0757_/a_68_297# net243 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7944 _0380_ _0757_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7945 VPWR _0350_ _0757_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7946 _0380_ _0757_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7947 _0757_/a_150_297# net243 _0757_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7948 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7949 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7950 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7951 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7952 VPWR acc0.A\[26\] _0688_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7953 VGND acc0.A\[26\] _0320_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7954 _0688_/a_109_297# net54 _0320_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7955 _0320_ net54 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7956 net137 clknet_1_1__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7957 VGND clknet_1_1__leaf__0464_ net137 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7958 net137 clknet_1_1__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7959 VPWR clknet_1_1__leaf__0464_ net137 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7961 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7964 _0542_/a_240_47# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X7965 _0141_ _0542_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7966 VGND _0172_ _0542_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7967 _0542_/a_51_297# net195 _0542_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X7968 _0542_/a_149_47# _0203_ _0542_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X7969 _0542_/a_240_47# _0174_ _0542_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7970 VPWR _0172_ _0542_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7971 _0141_ _0542_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X7972 _0542_/a_149_47# net195 _0542_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7973 _0542_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7974 VPWR _0203_ _0542_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7975 _0542_/a_512_297# net19 _0542_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7976 VGND _0241_ _0611_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7977 _0611_/a_68_297# _0242_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7978 _0243_ _0611_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7979 VPWR _0241_ _0611_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7980 _0243_ _0611_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7981 _0611_/a_150_297# _0242_ _0611_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7982 acc0.A\[25\] _1025_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7983 _1025_/a_891_413# _1025_/a_193_47# _1025_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7984 _1025_/a_561_413# _1025_/a_27_47# _1025_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7985 VPWR net111 _1025_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7986 acc0.A\[25\] _1025_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7987 _1025_/a_381_47# net200 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7988 VGND _1025_/a_634_159# _1025_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7989 VPWR _1025_/a_891_413# _1025_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7990 _1025_/a_466_413# _1025_/a_193_47# _1025_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7991 VPWR _1025_/a_634_159# _1025_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7992 _1025_/a_634_159# _1025_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7993 _1025_/a_634_159# _1025_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7994 _1025_/a_975_413# _1025_/a_193_47# _1025_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7995 VGND _1025_/a_1059_315# _1025_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7996 _1025_/a_193_47# _1025_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7997 _1025_/a_891_413# _1025_/a_27_47# _1025_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7998 _1025_/a_592_47# _1025_/a_193_47# _1025_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7999 VPWR _1025_/a_1059_315# _1025_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8000 _1025_/a_1017_47# _1025_/a_27_47# _1025_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8001 _1025_/a_193_47# _1025_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8002 _1025_/a_466_413# _1025_/a_27_47# _1025_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8003 VGND _1025_/a_891_413# _1025_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8004 _1025_/a_381_47# net200 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8005 VGND net111 _1025_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8006 _0809_/a_81_21# _0289_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X8007 _0809_/a_299_297# _0289_ _0809_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X8008 VPWR _0809_/a_81_21# _0420_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8009 VPWR _0295_ _0809_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8010 VGND _0809_/a_81_21# _0420_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8011 VGND _0401_ _0809_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X8012 _0809_/a_299_297# _0401_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8013 _0809_/a_384_47# _0295_ _0809_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8014 VPWR net37 hold70/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8015 VGND hold70/a_285_47# hold70/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8016 net217 hold70/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8017 VGND net37 hold70/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8018 VPWR hold70/a_285_47# hold70/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8019 hold70/a_285_47# hold70/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8020 hold70/a_285_47# hold70/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8021 net217 hold70/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8022 VPWR acc0.A\[12\] hold81/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8023 VGND hold81/a_285_47# hold81/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8024 net228 hold81/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8025 VGND acc0.A\[12\] hold81/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8026 VPWR hold81/a_285_47# hold81/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8027 hold81/a_285_47# hold81/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8028 hold81/a_285_47# hold81/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8029 net228 hold81/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8030 VPWR net59 hold92/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8031 VGND hold92/a_285_47# hold92/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8032 net239 hold92/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8033 VGND net59 hold92/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8034 VPWR hold92/a_285_47# hold92/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8035 hold92/a_285_47# hold92/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8036 hold92/a_285_47# hold92/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8037 net239 hold92/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8038 _0525_/a_81_21# _0194_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X8039 _0525_/a_299_297# _0194_ _0525_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X8040 VPWR _0525_/a_81_21# _0149_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8041 VPWR net154 _0525_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8042 VGND _0525_/a_81_21# _0149_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8043 VGND _0179_ _0525_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X8044 _0525_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8045 _0525_/a_384_47# net154 _0525_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8048 net54 _1008_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8049 _1008_/a_891_413# _1008_/a_193_47# _1008_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8050 _1008_/a_561_413# _1008_/a_27_47# _1008_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8051 VPWR net94 _1008_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8052 net54 _1008_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8053 _1008_/a_381_47# _0106_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8054 VGND _1008_/a_634_159# _1008_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8055 VPWR _1008_/a_891_413# _1008_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8056 _1008_/a_466_413# _1008_/a_193_47# _1008_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8057 VPWR _1008_/a_634_159# _1008_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8058 _1008_/a_634_159# _1008_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8059 _1008_/a_634_159# _1008_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8060 _1008_/a_975_413# _1008_/a_193_47# _1008_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8061 VGND _1008_/a_1059_315# _1008_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8062 _1008_/a_193_47# _1008_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8063 _1008_/a_891_413# _1008_/a_27_47# _1008_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8064 _1008_/a_592_47# _1008_/a_193_47# _1008_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8065 VPWR _1008_/a_1059_315# _1008_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8066 _1008_/a_1017_47# _1008_/a_27_47# _1008_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8067 _1008_/a_193_47# _1008_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8068 _1008_/a_466_413# _1008_/a_27_47# _1008_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8069 VGND _1008_/a_891_413# _1008_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8070 _1008_/a_381_47# _0106_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8071 VGND net94 _1008_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8072 VPWR output60/a_27_47# pp[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8073 pp[31] output60/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8074 VPWR net60 output60/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8075 pp[31] output60/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8076 VGND output60/a_27_47# pp[31] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8077 VGND net60 output60/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8080 _0508_/a_81_21# _0185_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X8081 _0508_/a_299_297# _0185_ _0508_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X8082 VPWR _0508_/a_81_21# _0157_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8083 VPWR net228 _0508_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8084 VGND _0508_/a_81_21# _0157_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8085 VGND _0179_ _0508_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X8086 _0508_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8087 _0508_/a_384_47# net228 _0508_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8088 _0406_ _0790_/a_35_297# _0790_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X8089 _0406_ net42 _0790_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X8090 _0790_/a_35_297# net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8091 _0790_/a_117_297# net42 _0790_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X8092 VPWR net42 _0790_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8093 VGND acc0.A\[15\] _0790_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8094 VGND _0790_/a_35_297# _0406_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8095 _0790_/a_285_297# acc0.A\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8096 VPWR acc0.A\[15\] _0790_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8097 _0790_/a_285_47# acc0.A\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8098 net64 _0988_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8099 _0988_/a_891_413# _0988_/a_193_47# _0988_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8100 _0988_/a_561_413# _0988_/a_27_47# _0988_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8101 VPWR net74 _0988_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8102 net64 _0988_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8103 _0988_/a_381_47# _0086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8104 VGND _0988_/a_634_159# _0988_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8105 VPWR _0988_/a_891_413# _0988_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8106 _0988_/a_466_413# _0988_/a_193_47# _0988_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8107 VPWR _0988_/a_634_159# _0988_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8108 _0988_/a_634_159# _0988_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8109 _0988_/a_634_159# _0988_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8110 _0988_/a_975_413# _0988_/a_193_47# _0988_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8111 VGND _0988_/a_1059_315# _0988_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8112 _0988_/a_193_47# _0988_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8113 _0988_/a_891_413# _0988_/a_27_47# _0988_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8114 _0988_/a_592_47# _0988_/a_193_47# _0988_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8115 VPWR _0988_/a_1059_315# _0988_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8116 _0988_/a_1017_47# _0988_/a_27_47# _0988_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8117 _0988_/a_193_47# _0988_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8118 _0988_/a_466_413# _0988_/a_27_47# _0988_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8119 VGND _0988_/a_891_413# _0988_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8120 _0988_/a_381_47# _0086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8121 VGND net74 _0988_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8122 net90 clknet_1_0__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8123 VGND clknet_1_0__leaf__0460_ net90 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8124 net90 clknet_1_0__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8125 VPWR clknet_1_0__leaf__0460_ net90 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8126 VPWR _0267_ _0842_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8127 _0446_ _0842_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X8128 VGND _0267_ _0842_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8129 _0842_/a_59_75# _0263_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8130 _0446_ _0842_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8131 _0842_/a_145_75# _0263_ _0842_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X8132 _0392_ _0773_/a_35_297# _0773_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X8133 _0392_ _0388_ _0773_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X8134 _0773_/a_35_297# _0388_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8135 _0773_/a_117_297# _0388_ _0773_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X8136 VPWR _0388_ _0773_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8137 VGND _0386_ _0773_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8138 VGND _0773_/a_35_297# _0392_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8139 _0773_/a_285_297# _0386_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8140 VPWR _0386_ _0773_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8141 _0773_/a_285_47# _0386_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8146 comp0.B\[9\] _1041_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8147 _1041_/a_891_413# _1041_/a_193_47# _1041_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8148 _1041_/a_561_413# _1041_/a_27_47# _1041_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8149 VPWR net127 _1041_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8150 comp0.B\[9\] _1041_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8151 _1041_/a_381_47# net153 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8152 VGND _1041_/a_634_159# _1041_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8153 VPWR _1041_/a_891_413# _1041_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8154 _1041_/a_466_413# _1041_/a_193_47# _1041_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8155 VPWR _1041_/a_634_159# _1041_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8156 _1041_/a_634_159# _1041_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8157 _1041_/a_634_159# _1041_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8158 _1041_/a_975_413# _1041_/a_193_47# _1041_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8159 VGND _1041_/a_1059_315# _1041_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8160 _1041_/a_193_47# _1041_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8161 _1041_/a_891_413# _1041_/a_27_47# _1041_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8162 _1041_/a_592_47# _1041_/a_193_47# _1041_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8163 VPWR _1041_/a_1059_315# _1041_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8164 _1041_/a_1017_47# _1041_/a_27_47# _1041_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8165 _1041_/a_193_47# _1041_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8166 _1041_/a_466_413# _1041_/a_27_47# _1041_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8167 VGND _1041_/a_891_413# _1041_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8168 _1041_/a_381_47# net153 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8169 VGND net127 _1041_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8170 VGND _0258_ _0825_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8171 _0825_/a_68_297# _0432_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8172 _0433_ _0825_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8173 VPWR _0258_ _0825_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8174 _0433_ _0825_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8175 _0825_/a_150_297# _0432_ _0825_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8178 VPWR net54 _0687_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8179 _0319_ _0687_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X8180 VGND net54 _0687_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8181 _0687_/a_59_75# acc0.A\[26\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8182 _0319_ _0687_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8183 _0687_/a_145_75# acc0.A\[26\] _0687_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X8184 _0756_/a_377_297# _0225_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X8185 _0756_/a_47_47# _0378_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8186 _0756_/a_129_47# _0378_ _0756_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X8187 _0756_/a_285_47# _0378_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X8188 _0379_ _0756_/a_47_47# _0756_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X8189 VGND _0225_ _0756_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8190 VPWR _0225_ _0756_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8191 VPWR _0756_/a_47_47# _0379_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X8192 _0379_ _0378_ _0756_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8193 _0756_/a_285_47# _0225_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8198 VPWR net46 _0610_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8199 _0242_ _0610_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X8200 VGND net46 _0610_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8201 _0610_/a_59_75# acc0.A\[19\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8202 _0242_ _0610_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8203 _0610_/a_145_75# acc0.A\[19\] _0610_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X8204 VGND comp0.B\[11\] _0541_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8205 _0541_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8206 _0203_ _0541_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8207 VPWR comp0.B\[11\] _0541_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8208 _0203_ _0541_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8209 _0541_/a_150_297# _0176_ _0541_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8210 acc0.A\[24\] _1024_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8211 _1024_/a_891_413# _1024_/a_193_47# _1024_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8212 _1024_/a_561_413# _1024_/a_27_47# _1024_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8213 VPWR net110 _1024_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8214 acc0.A\[24\] _1024_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8215 _1024_/a_381_47# _0122_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8216 VGND _1024_/a_634_159# _1024_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8217 VPWR _1024_/a_891_413# _1024_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8218 _1024_/a_466_413# _1024_/a_193_47# _1024_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8219 VPWR _1024_/a_634_159# _1024_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8220 _1024_/a_634_159# _1024_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8221 _1024_/a_634_159# _1024_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8222 _1024_/a_975_413# _1024_/a_193_47# _1024_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8223 VGND _1024_/a_1059_315# _1024_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8224 _1024_/a_193_47# _1024_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8225 _1024_/a_891_413# _1024_/a_27_47# _1024_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8226 _1024_/a_592_47# _1024_/a_193_47# _1024_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8227 VPWR _1024_/a_1059_315# _1024_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8228 _1024_/a_1017_47# _1024_/a_27_47# _1024_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8229 _1024_/a_193_47# _1024_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8230 _1024_/a_466_413# _1024_/a_27_47# _1024_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8231 VGND _1024_/a_891_413# _1024_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8232 _1024_/a_381_47# _0122_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8233 VGND net110 _1024_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8234 _0808_/a_585_47# _0419_ _0808_/a_266_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.47125 ps=4.05 w=0.65 l=0.15
X8235 VGND _0417_ _0808_/a_266_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8236 VPWR _0808_/a_81_21# _0091_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8237 _0808_/a_81_21# _0345_ _0808_/a_585_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8238 VGND _0808_/a_81_21# _0091_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8239 _0808_/a_266_297# _0346_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0 ps=0 w=1 l=0.15
X8240 _0808_/a_368_297# _0417_ _0808_/a_266_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0 ps=0 w=1 l=0.15
X8241 _0808_/a_266_47# _0418_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8242 _0808_/a_266_47# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8243 _0808_/a_81_21# _0418_ _0808_/a_368_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.535 pd=5.07 as=0 ps=0 w=1 l=0.15
X8244 _0808_/a_81_21# _0345_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8245 VPWR _0419_ _0808_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8246 VGND _0347_ _0739_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X8247 _0739_/a_510_47# _0365_ _0739_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X8248 _0739_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X8249 VPWR _0365_ _0739_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8250 _0739_/a_79_21# _0364_ _0739_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X8251 _0739_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8252 _0739_/a_79_21# _0352_ _0739_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X8253 VPWR _0739_/a_79_21# _0106_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8254 VGND _0739_/a_79_21# _0106_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8255 _0739_/a_215_47# _0364_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8256 VPWR _0117_ hold60/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8257 VGND hold60/a_285_47# hold60/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8258 net207 hold60/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8259 VGND _0117_ hold60/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8260 VPWR hold60/a_285_47# hold60/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8261 hold60/a_285_47# hold60/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8262 hold60/a_285_47# hold60/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8263 net207 hold60/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8264 VPWR acc0.A\[1\] hold71/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8265 VGND hold71/a_285_47# hold71/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8266 net218 hold71/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8267 VGND acc0.A\[1\] hold71/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8268 VPWR hold71/a_285_47# hold71/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8269 hold71/a_285_47# hold71/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8270 hold71/a_285_47# hold71/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8271 net218 hold71/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8272 VPWR acc0.A\[13\] hold82/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8273 VGND hold82/a_285_47# hold82/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8274 net229 hold82/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8275 VGND acc0.A\[13\] hold82/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8276 VPWR hold82/a_285_47# hold82/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8277 hold82/a_285_47# hold82/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8278 hold82/a_285_47# hold82/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8279 net229 hold82/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8280 VPWR control0.state\[1\] hold93/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8281 VGND hold93/a_285_47# hold93/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8282 net240 hold93/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8283 VGND control0.state\[1\] hold93/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8284 VPWR hold93/a_285_47# hold93/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8285 hold93/a_285_47# hold93/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8286 hold93/a_285_47# hold93/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8287 net240 hold93/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8288 VPWR net12 _0524_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X8289 _0524_/a_27_297# _0186_ _0524_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X8290 VGND net12 _0524_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X8291 _0194_ _0524_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8292 _0524_/a_27_297# _0186_ _0524_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X8293 _0524_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8294 _0524_/a_373_47# _0180_ _0524_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8295 _0194_ _0524_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8296 _0524_/a_109_297# net148 _0524_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8297 _0524_/a_109_47# net148 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8298 net53 _1007_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8299 _1007_/a_891_413# _1007_/a_193_47# _1007_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8300 _1007_/a_561_413# _1007_/a_27_47# _1007_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8301 VPWR net93 _1007_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8302 net53 _1007_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8303 _1007_/a_381_47# _0105_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8304 VGND _1007_/a_634_159# _1007_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8305 VPWR _1007_/a_891_413# _1007_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8306 _1007_/a_466_413# _1007_/a_193_47# _1007_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8307 VPWR _1007_/a_634_159# _1007_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8308 _1007_/a_634_159# _1007_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8309 _1007_/a_634_159# _1007_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8310 _1007_/a_975_413# _1007_/a_193_47# _1007_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8311 VGND _1007_/a_1059_315# _1007_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8312 _1007_/a_193_47# _1007_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8313 _1007_/a_891_413# _1007_/a_27_47# _1007_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8314 _1007_/a_592_47# _1007_/a_193_47# _1007_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8315 VPWR _1007_/a_1059_315# _1007_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8316 _1007_/a_1017_47# _1007_/a_27_47# _1007_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8317 _1007_/a_193_47# _1007_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8318 _1007_/a_466_413# _1007_/a_27_47# _1007_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8319 VGND _1007_/a_891_413# _1007_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8320 _1007_/a_381_47# _0105_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8321 VGND net93 _1007_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8323 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8326 VPWR output50/a_27_47# pp[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8327 pp[22] output50/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8328 VPWR net50 output50/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8329 pp[22] output50/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8330 VGND output50/a_27_47# pp[22] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8331 VGND net50 output50/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8332 VPWR net61 output61/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X8333 VGND output61/a_27_47# pp[3] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X8334 VGND output61/a_27_47# pp[3] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8335 pp[3] output61/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X8336 pp[3] output61/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8337 VGND net61 output61/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X8338 VPWR output61/a_27_47# pp[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8339 pp[3] output61/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8340 pp[3] output61/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8341 VPWR output61/a_27_47# pp[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8342 VPWR net5 _0507_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X8343 _0507_/a_27_297# _0183_ _0507_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X8344 VGND net5 _0507_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X8345 _0185_ _0507_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8346 _0507_/a_27_297# _0183_ _0507_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X8347 _0507_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8348 _0507_/a_373_47# _0181_ _0507_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8349 _0185_ _0507_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8350 _0507_/a_109_297# acc0.A\[13\] _0507_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8351 _0507_/a_109_47# acc0.A\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8352 net63 _0987_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8353 _0987_/a_891_413# _0987_/a_193_47# _0987_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8354 _0987_/a_561_413# _0987_/a_27_47# _0987_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8355 VPWR net73 _0987_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8356 net63 _0987_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8357 _0987_/a_381_47# _0085_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8358 VGND _0987_/a_634_159# _0987_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8359 VPWR _0987_/a_891_413# _0987_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8360 _0987_/a_466_413# _0987_/a_193_47# _0987_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8361 VPWR _0987_/a_634_159# _0987_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8362 _0987_/a_634_159# _0987_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8363 _0987_/a_634_159# _0987_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8364 _0987_/a_975_413# _0987_/a_193_47# _0987_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8365 VGND _0987_/a_1059_315# _0987_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8366 _0987_/a_193_47# _0987_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8367 _0987_/a_891_413# _0987_/a_27_47# _0987_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8368 _0987_/a_592_47# _0987_/a_193_47# _0987_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8369 VPWR _0987_/a_1059_315# _0987_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8370 _0987_/a_1017_47# _0987_/a_27_47# _0987_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8371 _0987_/a_193_47# _0987_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8372 _0987_/a_466_413# _0987_/a_27_47# _0987_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8373 VGND _0987_/a_891_413# _0987_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8374 _0987_/a_381_47# _0085_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8375 VGND net73 _0987_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8376 net75 clknet_1_1__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8377 VGND clknet_1_1__leaf__0458_ net75 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8378 net75 clknet_1_1__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8379 VPWR clknet_1_1__leaf__0458_ net75 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8380 net77 clknet_1_0__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8381 VGND clknet_1_0__leaf__0458_ net77 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8382 net77 clknet_1_0__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8383 VPWR clknet_1_0__leaf__0458_ net77 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8388 VGND _0369_ _0772_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X8389 _0772_/a_510_47# _0391_ _0772_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X8390 _0772_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X8391 VPWR _0391_ _0772_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8392 _0772_/a_79_21# net223 _0772_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X8393 _0772_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8394 _0772_/a_79_21# _0352_ _0772_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X8395 VPWR _0772_/a_79_21# _0099_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8396 VGND _0772_/a_79_21# _0099_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8397 _0772_/a_215_47# net223 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8398 VGND _0347_ _0841_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X8399 _0841_/a_510_47# _0445_ _0841_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X8400 _0841_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X8401 VPWR _0445_ _0841_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8402 _0841_/a_79_21# _0444_ _0841_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X8403 _0841_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8404 _0841_/a_79_21# _0399_ _0841_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X8405 VPWR _0841_/a_79_21# _0084_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8406 VGND _0841_/a_79_21# _0084_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8407 _0841_/a_215_47# _0444_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X8411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X8412 comp0.B\[8\] _1040_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8413 _1040_/a_891_413# _1040_/a_193_47# _1040_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8414 _1040_/a_561_413# _1040_/a_27_47# _1040_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8415 VPWR net126 _1040_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8416 comp0.B\[8\] _1040_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8417 _1040_/a_381_47# net174 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8418 VGND _1040_/a_634_159# _1040_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8419 VPWR _1040_/a_891_413# _1040_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8420 _1040_/a_466_413# _1040_/a_193_47# _1040_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8421 VPWR _1040_/a_634_159# _1040_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8422 _1040_/a_634_159# _1040_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8423 _1040_/a_634_159# _1040_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8424 _1040_/a_975_413# _1040_/a_193_47# _1040_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8425 VGND _1040_/a_1059_315# _1040_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8426 _1040_/a_193_47# _1040_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8427 _1040_/a_891_413# _1040_/a_27_47# _1040_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8428 _1040_/a_592_47# _1040_/a_193_47# _1040_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8429 VPWR _1040_/a_1059_315# _1040_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8430 _1040_/a_1017_47# _1040_/a_27_47# _1040_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8431 _1040_/a_193_47# _1040_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8432 _1040_/a_466_413# _1040_/a_27_47# _1040_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8433 VGND _1040_/a_891_413# _1040_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8434 _1040_/a_381_47# net174 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8435 VGND net126 _1040_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8440 VPWR _0271_ _0824_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8441 _0432_ _0824_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X8442 VGND _0271_ _0824_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8443 _0824_/a_59_75# _0431_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8444 _0432_ _0824_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8445 _0824_/a_145_75# _0431_ _0824_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X8446 VPWR _0227_ _0755_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X8447 VGND _0227_ _0378_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8448 _0755_/a_109_297# _0374_ _0378_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8449 _0378_ _0374_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8450 _0686_/a_219_297# _0686_/a_27_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0 ps=0 w=0.42 l=0.15
X8451 VGND _0317_ _0686_/a_27_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8452 VPWR _0316_ _0686_/a_301_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8453 _0318_ _0686_/a_219_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8454 _0686_/a_301_297# _0686_/a_27_53# _0686_/a_219_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8455 _0318_ _0686_/a_219_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8456 _0686_/a_27_53# _0317_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0 ps=0 w=0.42 l=0.15
X8457 VGND _0316_ _0686_/a_219_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8458 net128 clknet_1_1__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8459 VGND clknet_1_1__leaf__0464_ net128 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8460 net128 clknet_1_1__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8461 VPWR clknet_1_1__leaf__0464_ net128 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8462 net142 clknet_1_1__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8463 VGND clknet_1_1__leaf__0465_ net142 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8464 net142 clknet_1_1__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8465 VPWR clknet_1_1__leaf__0465_ net142 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8466 _0540_/a_240_47# net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X8467 _0142_ _0540_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8468 VGND _0172_ _0540_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8469 _0540_/a_51_297# net193 _0540_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X8470 _0540_/a_149_47# _0202_ _0540_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X8471 _0540_/a_240_47# _0174_ _0540_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8472 VPWR _0172_ _0540_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X8473 _0142_ _0540_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X8474 _0540_/a_149_47# net193 _0540_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8475 _0540_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8476 VPWR _0202_ _0540_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8477 _0540_/a_512_297# net20 _0540_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8478 acc0.A\[23\] _1023_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8479 _1023_/a_891_413# _1023_/a_193_47# _1023_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8480 _1023_/a_561_413# _1023_/a_27_47# _1023_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8481 VPWR net109 _1023_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8482 acc0.A\[23\] _1023_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8483 _1023_/a_381_47# net177 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8484 VGND _1023_/a_634_159# _1023_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8485 VPWR _1023_/a_891_413# _1023_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8486 _1023_/a_466_413# _1023_/a_193_47# _1023_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8487 VPWR _1023_/a_634_159# _1023_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8488 _1023_/a_634_159# _1023_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8489 _1023_/a_634_159# _1023_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8490 _1023_/a_975_413# _1023_/a_193_47# _1023_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8491 VGND _1023_/a_1059_315# _1023_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8492 _1023_/a_193_47# _1023_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8493 _1023_/a_891_413# _1023_/a_27_47# _1023_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8494 _1023_/a_592_47# _1023_/a_193_47# _1023_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8495 VPWR _1023_/a_1059_315# _1023_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8496 _1023_/a_1017_47# _1023_/a_27_47# _1023_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8497 _1023_/a_193_47# _1023_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8498 _1023_/a_466_413# _1023_/a_27_47# _1023_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8499 VGND _1023_/a_891_413# _1023_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8500 _1023_/a_381_47# net177 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8501 VGND net109 _1023_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8502 VGND _0218_ _0807_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8503 _0807_/a_68_297# net246 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8504 _0419_ _0807_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8505 VPWR _0218_ _0807_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8506 _0419_ _0807_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8507 _0807_/a_150_297# net246 _0807_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8508 VGND _0350_ _0738_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8509 _0738_/a_68_297# net244 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8510 _0365_ _0738_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8511 VPWR _0350_ _0738_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8512 _0365_ _0738_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8513 _0738_/a_150_297# net244 _0738_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8514 _0301_ _0669_/a_29_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X8515 _0669_/a_111_297# _0300_ _0669_/a_29_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.26 as=0.1092 ps=1.36 w=0.42 l=0.15
X8516 _0301_ _0669_/a_29_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8517 _0669_/a_183_297# _0277_ _0669_/a_111_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1386 pd=1.5 as=0 ps=0 w=0.42 l=0.15
X8518 VPWR _0276_ _0669_/a_183_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8519 _0669_/a_29_53# _0277_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.74 as=0 ps=0 w=0.42 l=0.15
X8520 VGND _0300_ _0669_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8521 VGND _0276_ _0669_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8526 VPWR acc0.A\[27\] hold50/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8527 VGND hold50/a_285_47# hold50/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8528 net197 hold50/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8529 VGND acc0.A\[27\] hold50/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8530 VPWR hold50/a_285_47# hold50/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8531 hold50/a_285_47# hold50/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8532 hold50/a_285_47# hold50/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8533 net197 hold50/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8534 VPWR acc0.A\[30\] hold61/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8535 VGND hold61/a_285_47# hold61/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8536 net208 hold61/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8537 VGND acc0.A\[30\] hold61/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8538 VPWR hold61/a_285_47# hold61/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8539 hold61/a_285_47# hold61/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8540 hold61/a_285_47# hold61/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8541 net208 hold61/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8542 VPWR acc0.A\[17\] hold72/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8543 VGND hold72/a_285_47# hold72/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8544 net219 hold72/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8545 VGND acc0.A\[17\] hold72/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8546 VPWR hold72/a_285_47# hold72/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8547 hold72/a_285_47# hold72/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8548 hold72/a_285_47# hold72/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8549 net219 hold72/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8550 VPWR acc0.A\[6\] hold83/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8551 VGND hold83/a_285_47# hold83/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8552 net230 hold83/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8553 VGND acc0.A\[6\] hold83/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8554 VPWR hold83/a_285_47# hold83/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8555 hold83/a_285_47# hold83/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8556 hold83/a_285_47# hold83/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8557 net230 hold83/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8558 VPWR net51 hold94/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8559 VGND hold94/a_285_47# hold94/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8560 net241 hold94/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8561 VGND net51 hold94/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8562 VPWR hold94/a_285_47# hold94/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8563 hold94/a_285_47# hold94/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8564 hold94/a_285_47# hold94/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8565 net241 hold94/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8568 net109 clknet_1_0__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8569 VGND clknet_1_0__leaf__0462_ net109 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8570 net109 clknet_1_0__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8571 VPWR clknet_1_0__leaf__0462_ net109 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8572 _0523_/a_81_21# _0193_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X8573 _0523_/a_299_297# _0193_ _0523_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X8574 VPWR _0523_/a_81_21# _0150_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8575 VPWR net148 _0523_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8576 VGND _0523_/a_81_21# _0150_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8577 VGND _0179_ _0523_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X8578 _0523_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8579 _0523_/a_384_47# net148 _0523_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8580 net52 _1006_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8581 _1006_/a_891_413# _1006_/a_193_47# _1006_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8582 _1006_/a_561_413# _1006_/a_27_47# _1006_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8583 VPWR net92 _1006_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8584 net52 _1006_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8585 _1006_/a_381_47# _0104_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8586 VGND _1006_/a_634_159# _1006_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8587 VPWR _1006_/a_891_413# _1006_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8588 _1006_/a_466_413# _1006_/a_193_47# _1006_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8589 VPWR _1006_/a_634_159# _1006_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8590 _1006_/a_634_159# _1006_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8591 _1006_/a_634_159# _1006_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8592 _1006_/a_975_413# _1006_/a_193_47# _1006_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8593 VGND _1006_/a_1059_315# _1006_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8594 _1006_/a_193_47# _1006_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8595 _1006_/a_891_413# _1006_/a_27_47# _1006_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8596 _1006_/a_592_47# _1006_/a_193_47# _1006_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8597 VPWR _1006_/a_1059_315# _1006_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8598 _1006_/a_1017_47# _1006_/a_27_47# _1006_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8599 _1006_/a_193_47# _1006_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8600 _1006_/a_466_413# _1006_/a_27_47# _1006_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8601 VGND _1006_/a_891_413# _1006_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8602 _1006_/a_381_47# _0104_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8603 VGND net92 _1006_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X8607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X8608 VPWR output51/a_27_47# pp[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8609 pp[23] output51/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8610 VPWR net51 output51/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8611 pp[23] output51/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8612 VGND output51/a_27_47# pp[23] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8613 VGND net51 output51/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8614 VPWR output40/a_27_47# pp[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8615 pp[13] output40/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8616 VPWR net40 output40/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8617 pp[13] output40/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8618 VGND output40/a_27_47# pp[13] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8619 VGND net40 output40/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8620 VPWR net62 output62/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X8621 VGND output62/a_27_47# pp[4] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X8622 VGND output62/a_27_47# pp[4] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8623 pp[4] output62/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X8624 pp[4] output62/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8625 VGND net62 output62/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X8626 VPWR output62/a_27_47# pp[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8627 pp[4] output62/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8628 pp[4] output62/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8629 VPWR output62/a_27_47# pp[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8632 _0506_/a_81_21# _0184_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X8633 _0506_/a_299_297# _0184_ _0506_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X8634 VPWR _0506_/a_81_21# _0158_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8635 VPWR net229 _0506_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8636 VGND _0506_/a_81_21# _0158_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8637 VGND _0179_ _0506_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X8638 _0506_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8639 _0506_/a_384_47# net229 _0506_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X8643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X8644 net62 _0986_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8645 _0986_/a_891_413# _0986_/a_193_47# _0986_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8646 _0986_/a_561_413# _0986_/a_27_47# _0986_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8647 VPWR net72 _0986_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8648 net62 _0986_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8649 _0986_/a_381_47# _0084_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8650 VGND _0986_/a_634_159# _0986_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8651 VPWR _0986_/a_891_413# _0986_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8652 _0986_/a_466_413# _0986_/a_193_47# _0986_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8653 VPWR _0986_/a_634_159# _0986_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8654 _0986_/a_634_159# _0986_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8655 _0986_/a_634_159# _0986_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8656 _0986_/a_975_413# _0986_/a_193_47# _0986_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8657 VGND _0986_/a_1059_315# _0986_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8658 _0986_/a_193_47# _0986_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8659 _0986_/a_891_413# _0986_/a_27_47# _0986_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8660 _0986_/a_592_47# _0986_/a_193_47# _0986_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8661 VPWR _0986_/a_1059_315# _0986_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8662 _0986_/a_1017_47# _0986_/a_27_47# _0986_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8663 _0986_/a_193_47# _0986_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8664 _0986_/a_466_413# _0986_/a_27_47# _0986_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8665 VGND _0986_/a_891_413# _0986_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8666 _0986_/a_381_47# _0084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8667 VGND net72 _0986_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8668 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8669 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8670 _0771_/a_298_297# _0771_/a_27_413# _0771_/a_215_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.535 pd=5.07 as=0.265 ps=2.53 w=1 l=0.15
X8671 _0771_/a_215_297# _0771_/a_27_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8672 _0771_/a_298_297# _0389_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8673 _0391_ _0771_/a_215_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8674 VPWR _0390_ _0771_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8675 _0391_ _0771_/a_215_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8676 _0771_/a_382_47# _0243_ _0771_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8677 VGND _0390_ _0771_/a_27_413# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X8678 VPWR _0243_ _0771_/a_298_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8679 VGND _0389_ _0771_/a_382_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8680 VGND _0218_ _0840_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8681 _0840_/a_68_297# net62 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8682 _0445_ _0840_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8683 VPWR _0218_ _0840_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8684 _0445_ _0840_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8685 _0840_/a_150_297# net62 _0840_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8686 VPWR _0468_ _0969_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X8687 VGND _0468_ _0487_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8688 _0969_/a_109_297# _0486_ _0487_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8689 _0487_ _0486_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8692 _0754_/a_240_47# net241 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X8693 _0103_ _0754_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8694 VGND _0219_ _0754_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8695 _0754_/a_51_297# _0377_ _0754_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X8696 _0754_/a_149_47# _0345_ _0754_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X8697 _0754_/a_240_47# _0376_ _0754_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8698 VPWR _0219_ _0754_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X8699 _0103_ _0754_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X8700 _0754_/a_149_47# _0377_ _0754_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8701 _0754_/a_245_297# _0376_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8702 VPWR _0345_ _0754_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8703 _0754_/a_512_297# net241 _0754_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8704 VPWR _0260_ _0823_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X8705 VGND _0260_ _0431_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8706 _0823_/a_109_297# _0269_ _0431_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8707 _0431_ _0269_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8708 VGND acc0.A\[27\] _0685_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8709 _0685_/a_68_297# net55 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8710 _0317_ _0685_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8711 VPWR acc0.A\[27\] _0685_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8712 _0317_ _0685_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8713 _0685_/a_150_297# net55 _0685_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X8715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X8716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8718 acc0.A\[22\] _1022_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8719 _1022_/a_891_413# _1022_/a_193_47# _1022_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8720 _1022_/a_561_413# _1022_/a_27_47# _1022_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8721 VPWR net108 _1022_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8722 acc0.A\[22\] _1022_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8723 _1022_/a_381_47# net151 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8724 VGND _1022_/a_634_159# _1022_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8725 VPWR _1022_/a_891_413# _1022_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8726 _1022_/a_466_413# _1022_/a_193_47# _1022_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8727 VPWR _1022_/a_634_159# _1022_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8728 _1022_/a_634_159# _1022_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8729 _1022_/a_634_159# _1022_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8730 _1022_/a_975_413# _1022_/a_193_47# _1022_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8731 VGND _1022_/a_1059_315# _1022_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8732 _1022_/a_193_47# _1022_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8733 _1022_/a_891_413# _1022_/a_27_47# _1022_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8734 _1022_/a_592_47# _1022_/a_193_47# _1022_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8735 VPWR _1022_/a_1059_315# _1022_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8736 _1022_/a_1017_47# _1022_/a_27_47# _1022_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8737 _1022_/a_193_47# _1022_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8738 _1022_/a_466_413# _1022_/a_27_47# _1022_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8739 VGND _1022_/a_891_413# _1022_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8740 _1022_/a_381_47# net151 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8741 VGND net108 _1022_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X8743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X8744 VPWR _0297_ _0668_/a_382_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.305 ps=2.61 w=1 l=0.15
X8745 _0668_/a_297_47# _0299_ _0668_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.3705 pd=3.74 as=0.169 ps=1.82 w=0.65 l=0.15
X8746 _0668_/a_297_47# _0297_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8747 VGND _0298_ _0668_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8748 VPWR _0668_/a_79_21# _0300_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X8749 _0668_/a_79_21# _0299_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.15
X8750 _0668_/a_382_297# _0298_ _0668_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8751 VGND _0668_/a_79_21# _0300_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8752 _0364_ _0737_/a_35_297# _0737_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X8753 _0364_ _0360_ _0737_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X8754 _0737_/a_35_297# _0360_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8755 _0737_/a_117_297# _0360_ _0737_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X8756 VPWR _0360_ _0737_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8757 VGND _0321_ _0737_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8758 VGND _0737_/a_35_297# _0364_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8759 _0737_/a_285_297# _0321_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8760 VPWR _0321_ _0737_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8761 _0737_/a_285_47# _0321_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8762 _0806_/a_199_47# _0281_ _0418_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X8763 _0806_/a_113_297# _0402_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X8764 _0418_ _0286_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8765 VPWR _0281_ _0806_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8766 _0806_/a_113_297# _0286_ _0418_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X8767 VGND _0402_ _0806_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8768 VPWR acc0.A\[23\] _0231_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8769 _0231_ acc0.A\[23\] _0599_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X8770 _0599_/a_113_47# net51 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8771 _0231_ net51 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8774 VPWR acc0.A\[20\] hold40/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8775 VGND hold40/a_285_47# hold40/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8776 net187 hold40/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8777 VGND acc0.A\[20\] hold40/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8778 VPWR hold40/a_285_47# hold40/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8779 hold40/a_285_47# hold40/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8780 hold40/a_285_47# hold40/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8781 net187 hold40/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8782 VPWR comp0.B\[11\] hold51/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8783 VGND hold51/a_285_47# hold51/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8784 net198 hold51/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8785 VGND comp0.B\[11\] hold51/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8786 VPWR hold51/a_285_47# hold51/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8787 hold51/a_285_47# hold51/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8788 hold51/a_285_47# hold51/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8789 net198 hold51/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8790 VPWR _0128_ hold62/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8791 VGND hold62/a_285_47# hold62/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8792 net209 hold62/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8793 VGND _0128_ hold62/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8794 VPWR hold62/a_285_47# hold62/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8795 hold62/a_285_47# hold62/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8796 hold62/a_285_47# hold62/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8797 net209 hold62/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8798 VPWR net48 hold73/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8799 VGND hold73/a_285_47# hold73/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8800 net220 hold73/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8801 VGND net48 hold73/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8802 VPWR hold73/a_285_47# hold73/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8803 hold73/a_285_47# hold73/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8804 hold73/a_285_47# hold73/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8805 net220 hold73/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8806 VPWR control0.sh hold84/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8807 VGND hold84/a_285_47# hold84/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8808 net231 hold84/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8809 VGND control0.sh hold84/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8810 VPWR hold84/a_285_47# hold84/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8811 hold84/a_285_47# hold84/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8812 hold84/a_285_47# hold84/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8813 net231 hold84/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8814 VPWR net56 hold95/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8815 VGND hold95/a_285_47# hold95/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8816 net242 hold95/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8817 VGND net56 hold95/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8818 VPWR hold95/a_285_47# hold95/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8819 hold95/a_285_47# hold95/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8820 hold95/a_285_47# hold95/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8821 net242 hold95/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8822 VPWR net13 _0522_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X8823 _0522_/a_27_297# _0186_ _0522_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X8824 VGND net13 _0522_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X8825 _0193_ _0522_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8826 _0522_/a_27_297# _0186_ _0522_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X8827 _0522_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8828 _0522_/a_373_47# _0180_ _0522_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8829 _0193_ _0522_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8830 _0522_/a_109_297# acc0.A\[6\] _0522_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8831 _0522_/a_109_47# acc0.A\[6\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8834 net51 _1005_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8835 _1005_/a_891_413# _1005_/a_193_47# _1005_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8836 _1005_/a_561_413# _1005_/a_27_47# _1005_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8837 VPWR net91 _1005_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8838 net51 _1005_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8839 _1005_/a_381_47# _0103_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8840 VGND _1005_/a_634_159# _1005_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8841 VPWR _1005_/a_891_413# _1005_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8842 _1005_/a_466_413# _1005_/a_193_47# _1005_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8843 VPWR _1005_/a_634_159# _1005_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8844 _1005_/a_634_159# _1005_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8845 _1005_/a_634_159# _1005_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8846 _1005_/a_975_413# _1005_/a_193_47# _1005_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8847 VGND _1005_/a_1059_315# _1005_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8848 _1005_/a_193_47# _1005_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8849 _1005_/a_891_413# _1005_/a_27_47# _1005_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8850 _1005_/a_592_47# _1005_/a_193_47# _1005_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8851 VPWR _1005_/a_1059_315# _1005_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8852 _1005_/a_1017_47# _1005_/a_27_47# _1005_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8853 _1005_/a_193_47# _1005_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8854 _1005_/a_466_413# _1005_/a_27_47# _1005_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8855 VGND _1005_/a_891_413# _1005_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8856 _1005_/a_381_47# _0103_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8857 VGND net91 _1005_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8858 VPWR output52/a_27_47# pp[24] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8859 pp[24] output52/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8860 VPWR net52 output52/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8861 pp[24] output52/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8862 VGND output52/a_27_47# pp[24] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8863 VGND net52 output52/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8864 VPWR output41/a_27_47# pp[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8865 pp[14] output41/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8866 VPWR net41 output41/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8867 pp[14] output41/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8868 VGND output41/a_27_47# pp[14] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8869 VGND net41 output41/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8870 VPWR net63 output63/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X8871 VGND output63/a_27_47# pp[5] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X8872 VGND output63/a_27_47# pp[5] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8873 pp[5] output63/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X8874 pp[5] output63/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8875 VGND net63 output63/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X8876 VPWR output63/a_27_47# pp[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8877 pp[5] output63/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8878 pp[5] output63/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8879 VPWR output63/a_27_47# pp[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X8883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X8884 VPWR net6 _0505_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X8885 _0505_/a_27_297# _0183_ _0505_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X8886 VGND net6 _0505_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X8887 _0184_ _0505_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8888 _0505_/a_27_297# _0183_ _0505_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X8889 _0505_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8890 _0505_/a_373_47# _0181_ _0505_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8891 _0184_ _0505_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8892 _0505_/a_109_297# acc0.A\[14\] _0505_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8893 _0505_/a_109_47# acc0.A\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
C0 _0199_ control0.sh 0
C1 _0118_ _0208_ 0.00135f
C2 VPWR _1005_/a_891_413# 0.19141f
C3 clknet_1_1__leaf__0459_ hold91/a_49_47# 0
C4 _0790_/a_285_297# _0406_ 0.07186f
C5 _0731_/a_384_47# VPWR 0.00171f
C6 clkbuf_0__0463_/a_110_47# _0494_/a_27_47# 0.00886f
C7 net21 _0473_ 0.01525f
C8 net103 _0219_ 0.00486f
C9 _0985_/a_1059_315# _0844_/a_79_21# 0
C10 _0157_ _0289_ 0
C11 clkbuf_1_1__f__0462_/a_110_47# _1010_/a_466_413# 0
C12 hold33/a_391_47# net22 0
C13 _0463_ _0913_/a_27_47# 0.11004f
C14 hold30/a_49_47# _1023_/a_891_413# 0
C15 hold30/a_391_47# _1023_/a_466_413# 0
C16 output39/a_27_47# _0994_/a_1059_315# 0
C17 _1001_/a_27_47# _1001_/a_193_47# 0.96327f
C18 _0390_ _0386_ 0
C19 _0243_ _0388_ 0.01017f
C20 pp[28] _1030_/a_634_159# 0
C21 net88 net1 0
C22 _0627_/a_109_93# _0274_ 0
C23 net23 clknet_1_0__leaf__0457_ 0.01769f
C24 net189 _0514_/a_109_297# 0
C25 _1057_/a_381_47# net2 0
C26 _1038_/a_891_413# net8 0
C27 _0176_ _1043_/a_1017_47# 0
C28 _0553_/a_51_297# _0957_/a_32_297# 0
C29 _0399_ _0268_ 0
C30 _0217_ hold40/a_49_47# 0.03884f
C31 VPWR _0765_/a_297_297# 0.00799f
C32 _0717_/a_80_21# _0333_ 0.08355f
C33 _1039_/a_975_413# _0473_ 0
C34 _1039_/a_381_47# _0472_ 0.00513f
C35 hold9/a_49_47# _1008_/a_891_413# 0
C36 hold9/a_285_47# _1008_/a_1059_315# 0
C37 net21 clkbuf_1_1__f__0464_/a_110_47# 0.09737f
C38 acc0.A\[29\] acc0.A\[28\] 0.00288f
C39 hold7/a_285_47# _0186_ 0
C40 _0958_/a_303_47# _0471_ 0
C41 net233 _0219_ 0.16267f
C42 _0235_ _0764_/a_81_21# 0
C43 _0339_ _0333_ 0.03397f
C44 _0811_/a_299_297# net228 0.00166f
C45 _0399_ _0090_ 0
C46 _0532_/a_299_297# net175 0
C47 _0198_ _0531_/a_109_47# 0.00201f
C48 _1049_/a_27_47# _1048_/a_466_413# 0
C49 _1049_/a_466_413# _1048_/a_27_47# 0
C50 _1049_/a_634_159# _1048_/a_193_47# 0
C51 acc0.A\[29\] net209 0
C52 _0462_ _0237_ 0
C53 _0225_ _0222_ 0.55444f
C54 hold33/a_391_47# clknet_1_0__leaf__0463_ 0.00491f
C55 hold44/a_285_47# net191 0.00983f
C56 _0461_ net149 0.00163f
C57 clknet_1_1__leaf__0460_ _0310_ 0
C58 hold8/a_49_47# hold8/a_285_47# 0.22264f
C59 VPWR _1011_/a_975_413# 0.00464f
C60 _0375_ _0369_ 0
C61 _0234_ _0383_ 0.00747f
C62 _0429_ _0253_ 0
C63 hold54/a_49_47# _0113_ 0.09107f
C64 _0485_ hold84/a_49_47# 0
C65 VPWR _1006_/a_466_413# 0.26928f
C66 _0678_/a_68_297# net43 0
C67 net36 _0347_ 0
C68 _1055_/a_466_413# A[10] 0
C69 net194 _0538_/a_51_297# 0
C70 _0699_/a_68_297# acc0.A\[28\] 0.18009f
C71 _0736_/a_139_47# _0350_ 0.00195f
C72 acc0.A\[5\] _0835_/a_78_199# 0
C73 _0195_ _1030_/a_891_413# 0.0206f
C74 _0216_ _1030_/a_466_413# 0
C75 net48 _1005_/a_891_413# 0.0213f
C76 VPWR _0986_/a_466_413# 0.265f
C77 acc0.A\[18\] _0773_/a_35_297# 0
C78 _1046_/a_27_47# _1061_/a_27_47# 0
C79 A[10] net181 0.25482f
C80 _0287_ net67 0.02876f
C81 _1019_/a_975_413# _0345_ 0.00255f
C82 _0714_/a_149_47# _0345_ 0.00154f
C83 _0985_/a_1059_315# _0846_/a_240_47# 0
C84 _0550_/a_512_297# _0176_ 0
C85 pp[9] _1058_/a_193_47# 0
C86 net118 _1067_/a_1059_315# 0
C87 _0742_/a_299_297# _0742_/a_384_47# 0
C88 _0951_/a_109_93# _0951_/a_296_53# 0
C89 net64 net182 0
C90 _0199_ net157 0.01586f
C91 _1013_/a_193_47# _0567_/a_27_297# 0
C92 _1013_/a_27_47# _0567_/a_109_297# 0
C93 _0769_/a_299_297# _0462_ 0
C94 _0701_/a_80_21# _0332_ 0.14907f
C95 _1012_/a_592_47# _0110_ 0
C96 _1004_/a_27_47# _0216_ 0.03401f
C97 _0161_ hold93/a_49_47# 0
C98 _0175_ _0560_/a_68_297# 0.12736f
C99 net34 input34/a_27_47# 0.10943f
C100 _0224_ _0103_ 0
C101 _0093_ pp[14] 0.0013f
C102 control0.state\[0\] _0972_/a_584_47# 0.0025f
C103 control0.state\[1\] _0972_/a_346_47# 0.0067f
C104 net46 _0592_/a_68_297# 0
C105 _0216_ _0126_ 0.00158f
C106 _0276_ VPWR 0.42181f
C107 net48 _0765_/a_297_297# 0.00847f
C108 net23 _1062_/a_466_413# 0
C109 _1072_/a_193_47# _1068_/a_27_47# 0
C110 _1072_/a_27_47# _1068_/a_193_47# 0
C111 _0180_ _0522_/a_109_297# 0.02121f
C112 _0532_/a_384_47# _0147_ 0
C113 clkbuf_1_0__f__0461_/a_110_47# _0612_/a_59_75# 0.01201f
C114 _0571_/a_109_47# VPWR 0
C115 comp0.B\[13\] _0538_/a_245_297# 0
C116 _0957_/a_32_297# _0561_/a_149_47# 0
C117 net95 _1009_/a_891_413# 0
C118 clkbuf_0__0464_/a_110_47# comp0.B\[10\] 0
C119 net55 _0322_ 0.20259f
C120 _0183_ clknet_1_1__leaf__0457_ 0
C121 _0289_ acc0.A\[9\] 0.05394f
C122 _0960_/a_27_47# _0169_ 0
C123 _1003_/a_891_413# acc0.A\[21\] 0.00257f
C124 _1003_/a_1059_315# _0227_ 0
C125 _0478_ _1072_/a_27_47# 0
C126 net55 _0327_ 0.36394f
C127 hold75/a_391_47# _0350_ 0.00112f
C128 _1035_/a_634_159# _0208_ 0
C129 _1035_/a_27_47# _0132_ 0.00283f
C130 _1035_/a_891_413# _0173_ 0
C131 net121 _0561_/a_51_297# 0
C132 _0236_ _0345_ 0.644f
C133 _1047_/a_27_47# _1047_/a_466_413# 0.27314f
C134 _1047_/a_193_47# _1047_/a_634_159# 0.11564f
C135 _0255_ _0269_ 0
C136 comp0.B\[8\] _1040_/a_891_413# 0.03417f
C137 _0206_ _1040_/a_1059_315# 0.01602f
C138 acc0.A\[16\] net84 0
C139 hold97/a_285_47# _0317_ 0.00358f
C140 _0957_/a_114_297# _0473_ 0
C141 net216 net52 0.25543f
C142 net53 _0367_ 0
C143 _0248_ _0372_ 0.43613f
C144 _0342_ VPWR 0.55477f
C145 _0172_ _0463_ 0
C146 clknet_1_0__leaf__0460_ hold3/a_49_47# 0.00174f
C147 control0.add hold40/a_285_47# 0
C148 clknet_1_0__leaf__0462_ net177 0.02309f
C149 _1041_/a_634_159# _0174_ 0.0035f
C150 _0312_ _0352_ 0
C151 _0664_/a_79_21# _0664_/a_297_47# 0.03259f
C152 _0346_ _0112_ 0
C153 _0582_/a_373_47# net221 0
C154 _0328_ hold90/a_391_47# 0
C155 _1041_/a_1059_315# comp0.B\[10\] 0.00928f
C156 net234 _1014_/a_27_47# 0
C157 _0855_/a_299_297# _1014_/a_1059_315# 0
C158 _1001_/a_634_159# clknet_1_0__leaf__0461_ 0
C159 _1007_/a_193_47# _1007_/a_975_413# 0
C160 _1007_/a_466_413# _1007_/a_381_47# 0.03733f
C161 _1052_/a_634_159# _1052_/a_592_47# 0
C162 _1007_/a_1059_315# _1007_/a_891_413# 0.31086f
C163 net121 _0133_ 0.01071f
C164 _0177_ _0935_/a_27_47# 0.00322f
C165 hold96/a_285_47# _1004_/a_193_47# 0.00198f
C166 VPWR _0854_/a_79_21# 0.44645f
C167 _0177_ _1061_/a_193_47# 0.00207f
C168 _0837_/a_81_21# _0837_/a_585_47# 0.00695f
C169 _0837_/a_266_297# _0837_/a_266_47# 0
C170 _0443_ _0835_/a_78_199# 0.00127f
C171 _1058_/a_381_47# _1058_/a_561_413# 0.00123f
C172 _1058_/a_27_47# net144 0.21888f
C173 _1058_/a_891_413# _1058_/a_975_413# 0.00851f
C174 _0172_ _1044_/a_1059_315# 0.05641f
C175 _1020_/a_193_47# _0352_ 0.04092f
C176 hold69/a_49_47# _1006_/a_193_47# 0
C177 hold69/a_285_47# _1006_/a_27_47# 0
C178 _0179_ _1052_/a_1059_315# 0.00594f
C179 _0230_ net52 0
C180 VPWR _0334_ 0.67554f
C181 net45 _0240_ 0.0019f
C182 input15/a_75_212# pp[5] 0
C183 _0149_ _0172_ 0.10195f
C184 _0429_ net74 0
C185 net45 _0369_ 0.03416f
C186 net44 _0351_ 0
C187 _0550_/a_51_297# clkbuf_1_0__f__0463_/a_110_47# 0.00167f
C188 clknet_1_1__leaf__0463_ clknet_0_clk 0
C189 net149 _0465_ 0.04747f
C190 _1050_/a_193_47# net11 0.03157f
C191 _1003_/a_27_47# _0487_ 0.01358f
C192 _0261_ _0186_ 0.05003f
C193 _0971_/a_81_21# _0971_/a_299_297# 0.08213f
C194 input22/a_75_212# B[14] 0.1979f
C195 _0462_ _0392_ 0
C196 _1011_/a_1017_47# _0355_ 0
C197 _1011_/a_592_47# net227 0
C198 _1011_/a_381_47# _0109_ 0.13419f
C199 net119 _1065_/a_891_413# 0
C200 _1033_/a_193_47# control0.reset 0.01691f
C201 _1002_/a_561_413# VPWR 0.00317f
C202 _0637_/a_311_297# _0219_ 0
C203 clknet_1_1__leaf__0457_ acc0.A\[15\] 0.13024f
C204 hold74/a_391_47# _0183_ 0
C205 comp0.B\[11\] hold6/a_49_47# 0
C206 clkbuf_0_clk/a_110_47# _1063_/a_27_47# 0.00381f
C207 net61 _0989_/a_27_47# 0.00206f
C208 _0389_ _0616_/a_78_199# 0.00434f
C209 net117 net208 0
C210 _0983_/a_381_47# _0854_/a_79_21# 0
C211 _0617_/a_68_297# _1006_/a_27_47# 0.00771f
C212 _0429_ output61/a_27_47# 0.00932f
C213 _0253_ clknet_1_1__leaf__0458_ 0.00932f
C214 _1059_/a_27_47# _0277_ 0
C215 _1063_/a_27_47# _1063_/a_634_159# 0.13601f
C216 _0422_ _0345_ 0.0058f
C217 _0770_/a_79_21# clkbuf_1_0__f__0457_/a_110_47# 0
C218 _1058_/a_1059_315# _0186_ 0.02109f
C219 _0645_/a_47_47# net42 0.01759f
C220 _0176_ net29 0.09615f
C221 clkbuf_0_clk/a_110_47# _0974_/a_448_47# 0.0032f
C222 _0345_ hold62/a_391_47# 0.0049f
C223 _1027_/a_1059_315# hold50/a_285_47# 0
C224 _0252_ pp[3] 0
C225 _0090_ _0295_ 0
C226 _0346_ _0099_ 0.0265f
C227 net221 clknet_1_0__leaf__0461_ 0
C228 acc0.A\[20\] _0772_/a_79_21# 0
C229 hold80/a_285_47# hold80/a_391_47# 0.41909f
C230 _0195_ net135 0
C231 _0592_/a_150_297# VPWR 0.00228f
C232 _0218_ _0778_/a_68_297# 0.16918f
C233 _0974_/a_222_93# net159 0
C234 hold34/a_285_47# acc0.A\[10\] 0
C235 _1039_/a_193_47# _0177_ 0
C236 _0536_/a_149_47# clkbuf_0__0464_/a_110_47# 0
C237 net158 _1049_/a_27_47# 0
C238 _0984_/a_561_413# VPWR 0.00344f
C239 net63 _0989_/a_634_159# 0
C240 _0336_ hold92/a_285_47# 0
C241 net63 hold1/a_391_47# 0
C242 clkbuf_0__0462_/a_110_47# acc0.A\[25\] 0
C243 _0346_ _0359_ 0.09817f
C244 _0994_/a_592_47# _0218_ 0
C245 _0538_/a_245_297# comp0.B\[9\] 0
C246 clknet_0__0459_ _0670_/a_79_21# 0
C247 output44/a_27_47# acc0.A\[30\] 0.1005f
C248 control0.state\[1\] _0183_ 0
C249 _0981_/a_27_297# _0482_ 0
C250 _0509_/a_27_47# _0186_ 0.16484f
C251 _1011_/a_634_159# acc0.A\[29\] 0.004f
C252 _1004_/a_634_159# net90 0
C253 _0718_/a_47_47# _0333_ 0
C254 _1004_/a_193_47# _1024_/a_27_47# 0
C255 hold41/a_391_47# acc0.A\[10\] 0.00474f
C256 _0369_ _0990_/a_1059_315# 0.00238f
C257 _0183_ _0583_/a_109_47# 0
C258 clkbuf_1_0__f__0462_/a_110_47# _1007_/a_891_413# 0.0129f
C259 _1002_/a_561_413# net48 0
C260 _0308_ _0347_ 0.02458f
C261 _1060_/a_27_47# _1060_/a_634_159# 0.14145f
C262 hold97/a_391_47# clknet_1_1__leaf__0460_ 0.03783f
C263 hold43/a_285_47# _1028_/a_193_47# 0
C264 hold43/a_391_47# _1028_/a_27_47# 0
C265 net15 net65 0
C266 net40 _0797_/a_27_413# 0.02102f
C267 _0195_ net234 0.00845f
C268 _0399_ clkbuf_1_0__f__0461_/a_110_47# 0
C269 pp[26] _0195_ 0.21462f
C270 net54 _0216_ 0.05797f
C271 net196 _1042_/a_1059_315# 0.0039f
C272 _1012_/a_27_47# _0396_ 0
C273 _1030_/a_975_413# acc0.A\[30\] 0.002f
C274 _0273_ _0252_ 0.20052f
C275 _0273_ _0989_/a_381_47# 0
C276 clknet_1_1__leaf__0463_ _0955_/a_220_297# 0
C277 hold56/a_391_47# _1065_/a_193_47# 0
C278 _0179_ clknet_1_1__leaf__0457_ 0.06403f
C279 hold16/a_285_47# hold62/a_285_47# 0
C280 hold16/a_391_47# hold62/a_49_47# 0
C281 _0988_/a_466_413# _0988_/a_592_47# 0.00553f
C282 _0988_/a_634_159# _0988_/a_1017_47# 0
C283 _0856_/a_79_21# _0456_ 0.07732f
C284 _0787_/a_80_21# _0402_ 0.13549f
C285 _0601_/a_68_297# _0350_ 0.00995f
C286 _0553_/a_51_297# _0553_/a_240_47# 0.03076f
C287 output57/a_27_47# net227 0.00549f
C288 _1039_/a_891_413# _0136_ 0.0012f
C289 net120 clkbuf_1_1__f__0463_/a_110_47# 0.00702f
C290 net187 net87 0.10509f
C291 _0485_ _0471_ 0.00157f
C292 net46 net92 0
C293 _1053_/a_466_413# acc0.A\[7\] 0
C294 hold100/a_391_47# _0465_ 0.00397f
C295 clk _1062_/a_193_47# 0
C296 clkbuf_0_clk/a_110_47# _1062_/a_1059_315# 0
C297 _0305_ _0675_/a_150_297# 0
C298 _0782_/a_27_47# clknet_1_0__leaf__0461_ 0.03f
C299 clknet_1_1__leaf__0460_ net96 0.21333f
C300 _1041_/a_27_47# comp0.B\[8\] 0.00294f
C301 _0982_/a_466_413# _0465_ 0.00183f
C302 net10 net196 0
C303 _0953_/a_114_297# comp0.B\[10\] 0.00596f
C304 _0606_/a_215_297# hold94/a_285_47# 0
C305 _0606_/a_109_53# hold94/a_49_47# 0.00137f
C306 VPWR _1014_/a_193_47# 0.31819f
C307 net58 hold100/a_285_47# 0.08214f
C308 acc0.A\[2\] hold100/a_391_47# 0
C309 _0309_ _0780_/a_35_297# 0.00148f
C310 _0542_/a_149_47# net195 0.01274f
C311 _0430_ _0399_ 0.015f
C312 _0542_/a_512_297# net19 0
C313 _0111_ _1031_/a_466_413# 0
C314 hold101/a_391_47# VPWR 0.18193f
C315 _1056_/a_1059_315# _0369_ 0
C316 hold96/a_285_47# net199 0.0125f
C317 net47 _0186_ 0.01984f
C318 _0644_/a_47_47# _0399_ 0
C319 clknet_1_0__leaf__0465_ _0826_/a_219_297# 0
C320 _0982_/a_466_413# acc0.A\[2\] 0
C321 control0.count\[3\] net91 0
C322 _1001_/a_975_413# clknet_1_0__leaf__0457_ 0.00107f
C323 _0461_ _0393_ 0.11178f
C324 net82 _1060_/a_27_47# 0
C325 _0460_ _1062_/a_891_413# 0
C326 _0684_/a_145_75# _0318_ 0
C327 _0316_ _0686_/a_301_297# 0.00141f
C328 _0784_/a_113_47# _0399_ 0
C329 hold14/a_49_47# net121 0.00467f
C330 _0216_ _0584_/a_27_297# 0.12341f
C331 acc0.A\[3\] _0449_ 0
C332 _0399_ _0401_ 0
C333 _1035_/a_975_413# net27 0.00101f
C334 _0399_ acc0.A\[5\] 0.00365f
C335 _1021_/a_891_413# clknet_1_0__leaf__0457_ 0.00832f
C336 _1021_/a_466_413# _0460_ 0.004f
C337 _0701_/a_80_21# _0701_/a_209_47# 0.01013f
C338 clknet_1_1__leaf__0458_ net74 0.30084f
C339 net133 _1047_/a_466_413# 0
C340 B[15] B[4] 0.02168f
C341 _0626_/a_150_297# _0271_ 0
C342 hold67/a_285_47# _0179_ 0
C343 _0583_/a_109_47# acc0.A\[15\] 0
C344 _0580_/a_109_47# acc0.A\[19\] 0.00214f
C345 net194 net11 0
C346 _0278_ _0994_/a_381_47# 0
C347 _1059_/a_1059_315# _0673_/a_253_47# 0
C348 hold79/a_49_47# clknet_1_0__leaf_clk 0.05758f
C349 _1008_/a_891_413# _0739_/a_79_21# 0
C350 clknet_1_1__leaf__0460_ _0315_ 0.18411f
C351 _0536_/a_512_297# net147 0
C352 _0347_ _1008_/a_381_47# 0.00928f
C353 output59/a_27_47# VPWR 0.3031f
C354 _0399_ net222 0.22806f
C355 _0378_ _0374_ 0.11567f
C356 hold45/a_285_47# A[11] 0
C357 _0996_/a_193_47# hold91/a_391_47# 0
C358 _0997_/a_1017_47# _0218_ 0
C359 hold25/a_49_47# _1038_/a_27_47# 0.00248f
C360 _0644_/a_377_297# _0277_ 0.00354f
C361 _0276_ _0794_/a_110_297# 0
C362 pp[30] _1030_/a_1017_47# 0
C363 _0675_/a_68_297# net43 0.1005f
C364 _0538_/a_51_297# _1045_/a_27_47# 0
C365 clkload4/Y _1017_/a_27_47# 0
C366 hold13/a_391_47# _0957_/a_32_297# 0
C367 _0557_/a_240_47# control0.sh 0.00287f
C368 clknet_1_1__leaf__0459_ _0779_/a_79_21# 0
C369 _0467_ hold38/a_49_47# 0
C370 output42/a_27_47# _0405_ 0
C371 _0305_ _0181_ 0.89721f
C372 _0151_ acc0.A\[7\] 0
C373 _0664_/a_382_297# _0402_ 0.00165f
C374 _0267_ net72 0
C375 _0642_/a_298_297# _0988_/a_27_47# 0
C376 hold9/a_285_47# clknet_1_1__leaf__0462_ 0.02229f
C377 _0999_/a_1059_315# net42 0
C378 acc0.A\[29\] _0702_/a_113_47# 0
C379 _0947_/a_109_297# _0467_ 0.01129f
C380 net125 _0173_ 0
C381 _0346_ net228 0.11311f
C382 net234 _0081_ 0
C383 _1001_/a_193_47# _0772_/a_79_21# 0
C384 VPWR _0724_/a_113_297# 0.23916f
C385 hold30/a_391_47# net177 0.1316f
C386 _1001_/a_634_159# _1001_/a_1017_47# 0
C387 _1001_/a_466_413# _1001_/a_592_47# 0.00553f
C388 _0537_/a_68_297# clknet_1_1__leaf__0464_ 0.05327f
C389 _0336_ hold80/a_285_47# 0
C390 _0991_/a_193_47# _0345_ 0.00163f
C391 _1035_/a_27_47# net25 0.00136f
C392 _0399_ _0182_ 0
C393 _1062_/a_193_47# _1062_/a_592_47# 0
C394 _1062_/a_466_413# _1062_/a_561_413# 0.00772f
C395 _1062_/a_634_159# _1062_/a_975_413# 0
C396 _0487_ hold93/a_285_47# 0
C397 _1020_/a_27_47# _1032_/a_381_47# 0
C398 _1020_/a_381_47# _1032_/a_27_47# 0
C399 _1029_/a_193_47# clknet_1_1__leaf__0462_ 0
C400 _1011_/a_27_47# _0353_ 0.00365f
C401 clkbuf_0__0458_/a_110_47# _0840_/a_68_297# 0
C402 _0992_/a_466_413# net228 0
C403 hold38/a_49_47# comp0.B\[0\] 0.00192f
C404 _1021_/a_193_47# _1021_/a_891_413# 0.19685f
C405 _1021_/a_27_47# _1021_/a_381_47# 0.06222f
C406 _1021_/a_634_159# _1021_/a_1059_315# 0
C407 _1003_/a_381_47# net49 0
C408 net61 _0257_ 0.40789f
C409 _0518_/a_109_297# clknet_1_1__leaf__0458_ 0.0077f
C410 net199 _1024_/a_27_47# 0
C411 _0854_/a_79_21# _0453_ 0
C412 _0481_ _0489_ 0
C413 _0419_ net246 0.00751f
C414 _0147_ _1048_/a_27_47# 0
C415 _1049_/a_193_47# net134 0.03751f
C416 _0607_/a_27_297# _0399_ 0
C417 clknet_1_1__leaf__0461_ _0790_/a_35_297# 0
C418 net155 VPWR 0.50585f
C419 _0645_/a_47_47# _0645_/a_377_297# 0.00899f
C420 _0996_/a_1059_315# _0670_/a_79_21# 0
C421 _1037_/a_891_413# net27 0
C422 _0476_ hold84/a_391_47# 0.0022f
C423 _0329_ net114 0
C424 clkbuf_1_0__f__0463_/a_110_47# _0913_/a_27_47# 0
C425 hold64/a_49_47# net45 0
C426 _0791_/a_199_47# net41 0
C427 _0205_ _0545_/a_150_297# 0
C428 _0536_/a_240_47# _0953_/a_32_297# 0
C429 net117 _1031_/a_193_47# 0.01325f
C430 _0963_/a_285_47# control0.count\[0\] 0.00129f
C431 net179 A[10] 0.00173f
C432 _0443_ _0399_ 0.08246f
C433 VPWR _0548_/a_512_297# 0.00846f
C434 _0330_ _0332_ 0.27162f
C435 clkbuf_1_0__f__0465_/a_110_47# _0989_/a_193_47# 0
C436 clknet_1_1__leaf__0464_ _1043_/a_381_47# 0.01784f
C437 net57 _0568_/a_27_297# 0
C438 _0752_/a_300_297# _0378_ 0
C439 _0216_ _1015_/a_634_159# 0.00147f
C440 _0433_ _0825_/a_150_297# 0.00114f
C441 net157 _0498_/a_149_47# 0
C442 _0137_ _0176_ 0.03446f
C443 hold88/a_285_47# _0252_ 0
C444 _0763_/a_193_47# _0462_ 0
C445 _0585_/a_373_47# clknet_1_0__leaf__0461_ 0
C446 _0092_ _0994_/a_891_413# 0
C447 _1034_/a_466_413# clkbuf_1_1__f__0463_/a_110_47# 0.00707f
C448 _1034_/a_27_47# clknet_0__0463_ 0.00542f
C449 _1020_/a_891_413# _0721_/a_27_47# 0
C450 hold26/a_285_47# _0205_ 0
C451 _0258_ net63 0.00253f
C452 hold38/a_285_47# _1034_/a_193_47# 0
C453 _0225_ _1022_/a_466_413# 0
C454 _0714_/a_240_47# _0344_ 0.04114f
C455 hold34/a_391_47# _0181_ 0
C456 _0554_/a_68_297# _0209_ 0
C457 pp[10] _0186_ 0
C458 _0439_ _0369_ 0.27612f
C459 _0561_/a_149_47# _0213_ 0.00154f
C460 VPWR _0240_ 2.3886f
C461 net23 _0160_ 0.05426f
C462 hold29/a_285_47# _1022_/a_27_47# 0
C463 hold100/a_49_47# _0261_ 0.02205f
C464 hold90/a_49_47# _0105_ 0
C465 VPWR _0369_ 6.64798f
C466 _0251_ net235 0
C467 clknet_0__0457_ VPWR 3.32669f
C468 net181 _0514_/a_373_47# 0
C469 _0515_/a_81_21# net2 0.0029f
C470 _0259_ _0218_ 0
C471 _0982_/a_193_47# _0261_ 0
C472 net44 _0338_ 0
C473 net188 _0179_ 0.17965f
C474 _0760_/a_129_47# clknet_1_0__leaf__0460_ 0
C475 _1020_/a_193_47# net106 0.00468f
C476 net11 _0987_/a_193_47# 0.0132f
C477 _0618_/a_79_21# _0618_/a_215_47# 0.04584f
C478 _0473_ _0173_ 0.02885f
C479 _0252_ _0086_ 0
C480 hold39/a_49_47# _0175_ 0
C481 _1036_/a_561_413# clknet_1_1__leaf__0463_ 0
C482 _1036_/a_891_413# net122 0
C483 _0346_ _0792_/a_80_21# 0
C484 _1050_/a_1059_315# clknet_0__0464_ 0
C485 _0348_ _1030_/a_27_47# 0
C486 _0510_/a_27_297# _0181_ 0.11208f
C487 _0233_ _0315_ 0
C488 _0231_ _0366_ 0
C489 _0999_/a_193_47# _0307_ 0
C490 _0461_ _1019_/a_891_413# 0.00603f
C491 hold68/a_391_47# _0222_ 0
C492 _0538_/a_51_297# net132 0
C493 hold96/a_285_47# VPWR 0.28289f
C494 _0555_/a_51_297# _1037_/a_27_47# 0
C495 _0423_ _0345_ 0.01874f
C496 _0683_/a_113_47# _0345_ 0
C497 _0423_ _0814_/a_27_47# 0.22351f
C498 VPWR _0852_/a_117_297# 0.00604f
C499 clknet_1_0__leaf__0459_ _1014_/a_193_47# 0
C500 _1001_/a_634_159# _0218_ 0
C501 net121 _0208_ 0
C502 _1041_/a_634_159# comp0.B\[9\] 0
C503 _1041_/a_891_413# net153 0
C504 _1041_/a_381_47# net127 0.001f
C505 hold34/a_285_47# _0188_ 0
C506 _0329_ _0365_ 0
C507 _1047_/a_27_47# _0145_ 0.10676f
C508 _1047_/a_1059_315# _1047_/a_1017_47# 0
C509 _0723_/a_27_413# hold61/a_285_47# 0
C510 _1030_/a_1017_47# _0339_ 0
C511 clknet_1_1__leaf__0460_ _0742_/a_81_21# 0.00101f
C512 _1037_/a_891_413# _0136_ 0
C513 hold12/a_49_47# _0381_ 0
C514 net83 _0407_ 0
C515 _0401_ _0295_ 0.44341f
C516 _0111_ hold16/a_285_47# 0
C517 _0241_ net47 0
C518 hold25/a_391_47# VPWR 0.19135f
C519 clknet_1_0__leaf_clk _0970_/a_114_47# 0
C520 clknet_0__0465_ _0826_/a_27_53# 0.02113f
C521 _0256_ _0465_ 0.00401f
C522 _0961_/a_199_47# _0480_ 0
C523 net185 _0561_/a_240_47# 0.04111f
C524 control0.state\[0\] _0467_ 0.00574f
C525 _0973_/a_27_297# clknet_1_0__leaf__0461_ 0
C526 _0849_/a_297_297# _0219_ 0.00697f
C527 _0230_ hold94/a_391_47# 0
C528 output53/a_27_47# pp[25] 0.15955f
C529 pp[28] _0355_ 0
C530 net58 net235 0.00178f
C531 comp0.B\[6\] _0176_ 0.54545f
C532 _0461_ net206 0
C533 net188 _0513_/a_81_21# 0.10837f
C534 hold41/a_391_47# _0188_ 0.06451f
C535 _0183_ _1018_/a_1059_315# 0
C536 _0953_/a_32_297# _1046_/a_27_47# 0
C537 hold85/a_285_47# _0959_/a_80_21# 0
C538 _1004_/a_193_47# _0756_/a_47_47# 0
C539 net197 _0689_/a_68_297# 0
C540 _1007_/a_381_47# _0105_ 0.13242f
C541 hold22/a_391_47# _0152_ 0
C542 _0243_ _0216_ 0.06697f
C543 _0180_ _0150_ 0.0693f
C544 _0464_ net170 0
C545 _0536_/a_512_297# _0473_ 0
C546 _0536_/a_51_297# _0472_ 0
C547 net243 _1004_/a_381_47# 0
C548 hold88/a_49_47# net141 0.00152f
C549 _0446_ _0263_ 0.24854f
C550 _0450_ _0261_ 0.0048f
C551 _0502_/a_27_47# net8 0
C552 net197 _1027_/a_1017_47# 0
C553 _0126_ _1027_/a_891_413# 0
C554 _0217_ _0575_/a_27_297# 0.16541f
C555 net48 _0369_ 0.46345f
C556 _0387_ _0776_/a_109_297# 0
C557 clknet_0__0457_ net48 0
C558 clknet_1_1__leaf__0460_ _0309_ 0
C559 hold7/a_391_47# _0987_/a_193_47# 0.00186f
C560 hold7/a_49_47# _0987_/a_466_413# 0.00261f
C561 net58 _0858_/a_27_47# 0
C562 _0629_/a_145_75# _0458_ 0
C563 _1057_/a_634_159# net37 0
C564 _0370_ net52 0.00803f
C565 _0269_ _0843_/a_68_297# 0.01021f
C566 _0220_ _0336_ 0.48593f
C567 _0172_ clkbuf_1_0__f__0463_/a_110_47# 0
C568 _0429_ net61 0.05305f
C569 _0715_/a_27_47# _0347_ 0
C570 control0.state\[0\] comp0.B\[0\] 0
C571 _0301_ net41 0
C572 net57 _0109_ 0.00211f
C573 _0216_ net227 0.00292f
C574 _0960_/a_27_47# _0960_/a_109_47# 0.00517f
C575 _0218_ net221 0
C576 hold24/a_285_47# VPWR 0.29072f
C577 hold42/a_285_47# net67 0.00661f
C578 _1057_/a_1059_315# net67 0.00164f
C579 _0819_/a_299_297# net66 0
C580 _0982_/a_27_47# clknet_1_0__leaf__0461_ 0.00779f
C581 _0757_/a_150_297# acc0.A\[23\] 0
C582 hold25/a_285_47# _0550_/a_51_297# 0.00218f
C583 _1038_/a_193_47# net28 0
C584 _0130_ control0.reset 0
C585 clknet_0__0458_ _0433_ 0.02146f
C586 net220 _0462_ 0
C587 clknet_1_0__leaf__0458_ acc0.A\[18\] 0
C588 _0330_ _0738_/a_68_297# 0
C589 _0983_/a_592_47# _0455_ 0
C590 VPWR input7/a_75_212# 0.26163f
C591 net120 _0163_ 0
C592 _0390_ _0369_ 0
C593 _0326_ acc0.A\[23\] 0
C594 acc0.A\[12\] net38 0
C595 _1046_/a_891_413# net174 0
C596 _1063_/a_891_413# _1063_/a_975_413# 0.00851f
C597 _1063_/a_381_47# _1063_/a_561_413# 0.00123f
C598 A[6] net12 0
C599 _0836_/a_68_297# acc0.A\[8\] 0
C600 VPWR _0844_/a_79_21# 0.2402f
C601 net243 _0225_ 0
C602 clkbuf_1_1__f__0458_/a_110_47# _0434_ 0.03798f
C603 _0712_/a_79_21# _1013_/a_27_47# 0
C604 _0179_ _0155_ 0.11023f
C605 net45 pp[31] 0.0909f
C606 acc0.A\[20\] _1019_/a_27_47# 0
C607 _0399_ _0089_ 0
C608 acc0.A\[8\] net212 0
C609 _0305_ _0507_/a_373_47# 0
C610 hold100/a_49_47# net47 0
C611 hold19/a_391_47# _0115_ 0.00131f
C612 _1037_/a_1017_47# _0208_ 0
C613 VPWR _1024_/a_27_47# 0.68927f
C614 _0161_ clknet_1_0__leaf__0457_ 0
C615 _0585_/a_27_297# _0585_/a_373_47# 0.01338f
C616 _0462_ _1006_/a_592_47# 0
C617 _1071_/a_27_47# _0976_/a_505_21# 0
C618 _0982_/a_193_47# net47 0
C619 hold76/a_285_47# _0352_ 0
C620 net233 net58 0.19475f
C621 clknet_1_0__leaf__0464_ _1050_/a_466_413# 0.0013f
C622 _0748_/a_81_21# _0294_ 0.11014f
C623 _0305_ hold82/a_391_47# 0.02594f
C624 _0677_/a_47_47# net43 0.00123f
C625 net17 clknet_1_0__leaf__0461_ 0.13796f
C626 _0349_ _1012_/a_193_47# 0
C627 VPWR _1048_/a_634_159# 0.1828f
C628 net59 _0567_/a_27_297# 0
C629 net18 _0542_/a_51_297# 0.01959f
C630 _0544_/a_51_297# net19 0
C631 _0343_ net42 0.19747f
C632 _0855_/a_81_21# _0580_/a_27_297# 0
C633 _1028_/a_381_47# clknet_1_1__leaf__0462_ 0.00756f
C634 _1055_/a_27_47# acc0.A\[8\] 0
C635 hold57/a_285_47# _0175_ 0
C636 _0891_/a_27_47# _0721_/a_27_47# 0.00328f
C637 hold46/a_391_47# _0473_ 0
C638 _0131_ net24 0.03905f
C639 net214 _0291_ 0
C640 _0642_/a_27_413# _0253_ 0
C641 _0255_ clkbuf_0__0458_/a_110_47# 0
C642 _0260_ acc0.A\[3\] 0.16271f
C643 _0428_ clkbuf_0__0465_/a_110_47# 0.00603f
C644 _0312_ _0392_ 0
C645 _0170_ _0482_ 0
C646 _0195_ _0569_/a_373_47# 0
C647 net97 acc0.A\[29\] 0
C648 _0216_ _0569_/a_109_297# 0.00824f
C649 net197 net112 0
C650 _0570_/a_109_47# acc0.A\[26\] 0
C651 _0716_/a_27_47# _0403_ 0
C652 VPWR _1010_/a_381_47# 0.0765f
C653 _1000_/a_193_47# _1000_/a_891_413# 0.19329f
C654 _1000_/a_27_47# _1000_/a_381_47# 0.06222f
C655 _1000_/a_634_159# _1000_/a_1059_315# 0
C656 _0140_ net20 0
C657 _1060_/a_891_413# _1060_/a_975_413# 0.00851f
C658 _1060_/a_27_47# net146 0.26322f
C659 _1060_/a_381_47# _1060_/a_561_413# 0.00123f
C660 _1051_/a_193_47# net154 0.02015f
C661 _0513_/a_81_21# _0155_ 0.13864f
C662 hold57/a_391_47# control0.sh 0.04748f
C663 _0168_ _0979_/a_27_297# 0
C664 VPWR _0979_/a_109_47# 0
C665 net230 _0520_/a_373_47# 0
C666 _0151_ _0520_/a_109_297# 0.05529f
C667 _1072_/a_27_47# VPWR 0.43427f
C668 _0238_ _0346_ 0.0245f
C669 _0143_ _1050_/a_1017_47# 0
C670 clknet_1_1__leaf__0458_ _0987_/a_193_47# 0.00141f
C671 VPWR _0846_/a_240_47# 0.00134f
C672 _0233_ _0742_/a_81_21# 0
C673 _0609_/a_109_297# _0241_ 0.01509f
C674 _0320_ _0739_/a_79_21# 0
C675 net208 _0704_/a_68_297# 0
C676 _0553_/a_512_297# _0136_ 0
C677 _0805_/a_181_47# VPWR 0
C678 _0399_ _0986_/a_891_413# 0.00587f
C679 clknet_1_0__leaf__0459_ _0240_ 0
C680 _0973_/a_109_297# _1063_/a_1059_315# 0
C681 net62 net47 1.19133f
C682 net105 hold60/a_49_47# 0
C683 acc0.A\[27\] _0462_ 0
C684 pp[27] net208 0.00341f
C685 VPWR _1009_/a_561_413# 0.00316f
C686 acc0.A\[12\] hold81/a_285_47# 0.02061f
C687 _0698_/a_113_297# _0317_ 0.05024f
C688 hold36/a_391_47# clknet_1_1__leaf__0464_ 0
C689 clknet_1_0__leaf__0459_ _0369_ 0.23205f
C690 hold14/a_391_47# _0173_ 0
C691 _0450_ net47 0
C692 clknet_0__0457_ clknet_1_0__leaf__0459_ 0.16003f
C693 _0457_ _1033_/a_193_47# 0
C694 _0963_/a_35_297# _0963_/a_285_297# 0.02504f
C695 clknet_1_0__leaf__0458_ hold59/a_49_47# 0
C696 hold27/a_285_47# _1039_/a_193_47# 0
C697 _0080_ _0465_ 0.00584f
C698 hold27/a_391_47# _1039_/a_27_47# 0
C699 _0343_ _0379_ 0
C700 _0231_ _0378_ 0
C701 _0161_ _1062_/a_466_413# 0
C702 _0376_ acc0.A\[22\] 0
C703 _0236_ hold94/a_391_47# 0
C704 _0583_/a_109_297# net165 0.0015f
C705 clknet_1_0__leaf__0462_ hold4/a_49_47# 0.01353f
C706 _1071_/a_592_47# VPWR 0
C707 net19 _0141_ 0.00738f
C708 _1056_/a_634_159# net178 0
C709 _0998_/a_1059_315# _0097_ 0
C710 _0343_ _0372_ 0.04387f
C711 _0330_ _0701_/a_209_47# 0.00166f
C712 _0216_ _0567_/a_109_47# 0.00484f
C713 _0985_/a_891_413# _0179_ 0.02746f
C714 clknet_1_0__leaf__0457_ _0391_ 0.03534f
C715 acc0.A\[21\] clknet_1_0__leaf__0461_ 0
C716 clknet_1_1__leaf__0462_ _0739_/a_297_297# 0
C717 _0152_ _0255_ 0
C718 _0369_ _0283_ 0.00234f
C719 _0179_ _1049_/a_634_159# 0.04732f
C720 _0305_ clknet_1_1__leaf__0461_ 0.22802f
C721 _1018_/a_27_47# _0181_ 0
C722 clknet_1_1__leaf__0463_ _1065_/a_27_47# 0.00255f
C723 _0372_ net95 0
C724 net113 _0347_ 0
C725 _0497_/a_68_297# _0173_ 0
C726 _1059_/a_1059_315# _0219_ 0.001f
C727 _0119_ _0460_ 0.00495f
C728 _0684_/a_59_75# _0328_ 0
C729 net36 _0180_ 0.03068f
C730 _0701_/a_303_47# _0333_ 0
C731 _0621_/a_35_297# _0437_ 0
C732 net133 _0145_ 0.00182f
C733 _0573_/a_27_47# _1015_/a_1059_315# 0
C734 net36 net218 0.00321f
C735 _0311_ _0250_ 0.00114f
C736 _0858_/a_27_47# _0262_ 0
C737 _0997_/a_634_159# net41 0.01583f
C738 _0997_/a_27_47# pp[14] 0
C739 _0346_ _0268_ 0
C740 clknet_0__0464_ _1046_/a_891_413# 0.00385f
C741 hold11/a_285_47# net157 0.04296f
C742 net61 clknet_1_1__leaf__0458_ 0.04067f
C743 _1071_/a_634_159# clknet_0_clk 0
C744 hold79/a_285_47# clk 0.00133f
C745 net54 _1027_/a_891_413# 0.00168f
C746 net226 control0.count\[0\] 0
C747 _1008_/a_381_47# _0106_ 0.13113f
C748 _0959_/a_80_21# _0132_ 0
C749 _0346_ _0721_/a_27_47# 0
C750 pp[11] net38 0.01194f
C751 hold13/a_285_47# _0173_ 0
C752 hold13/a_391_47# _0213_ 0
C753 _0397_ _0676_/a_113_47# 0
C754 net185 B[4] 0
C755 hold64/a_49_47# VPWR 0.2669f
C756 net64 _1055_/a_27_47# 0
C757 _0257_ _0431_ 0.02022f
C758 net175 _1048_/a_1017_47# 0
C759 net9 _1048_/a_561_413# 0
C760 comp0.B\[11\] _1043_/a_891_413# 0.00679f
C761 _1055_/a_193_47# _0621_/a_35_297# 0
C762 _0346_ _0090_ 0
C763 _0328_ _0687_/a_145_75# 0
C764 control0.state\[2\] _1066_/a_27_47# 0
C765 _0153_ acc0.A\[10\] 0
C766 _1020_/a_466_413# _0578_/a_109_297# 0
C767 _1020_/a_1059_315# _0578_/a_27_297# 0
C768 _1000_/a_27_47# _1018_/a_466_413# 0
C769 _0119_ _0457_ 0
C770 control0.state\[2\] _1068_/a_27_47# 0
C771 net44 _0396_ 0.21454f
C772 net21 _1045_/a_193_47# 0.02873f
C773 net183 _1045_/a_634_159# 0
C774 _0201_ _1045_/a_1059_315# 0.00435f
C775 net22 _0204_ 0
C776 net149 _1047_/a_975_413# 0.00119f
C777 _0531_/a_109_297# clkbuf_1_1__f__0457_/a_110_47# 0
C778 VPWR _1022_/a_975_413# 0.00481f
C779 clk net17 0
C780 hold10/a_49_47# _0533_/a_27_297# 0.00654f
C781 clknet_1_0__leaf__0463_ _0552_/a_68_297# 0
C782 _0245_ clknet_1_0__leaf__0461_ 0
C783 _0650_/a_68_297# hold81/a_285_47# 0
C784 _0637_/a_139_47# _0465_ 0
C785 _0610_/a_59_75# acc0.A\[19\] 0.12219f
C786 _0852_/a_117_297# _0453_ 0.00595f
C787 _0852_/a_285_47# _0266_ 0
C788 net22 hold6/a_391_47# 0
C789 _0999_/a_1059_315# _0999_/a_891_413# 0.31086f
C790 _0999_/a_193_47# _0999_/a_975_413# 0
C791 _0999_/a_466_413# _0999_/a_381_47# 0.03733f
C792 net17 _1063_/a_891_413# 0.04385f
C793 net214 _0290_ 0.18018f
C794 _0992_/a_466_413# _0090_ 0
C795 _0992_/a_891_413# _0422_ 0
C796 _1001_/a_27_47# _1019_/a_193_47# 0.00217f
C797 _1001_/a_193_47# _1019_/a_27_47# 0.00314f
C798 _1017_/a_466_413# _0115_ 0.00312f
C799 _0772_/a_79_21# _0772_/a_297_297# 0.01735f
C800 _0972_/a_346_47# clknet_1_1__leaf_clk 0
C801 VPWR _0993_/a_27_47# 0.72354f
C802 _0833_/a_297_297# _0186_ 0.00409f
C803 _1001_/a_891_413# net223 0.02535f
C804 _1001_/a_1059_315# _0391_ 0
C805 _1001_/a_634_159# _0099_ 0.00197f
C806 _0340_ _1031_/a_891_413# 0.01063f
C807 net58 _0637_/a_311_297# 0
C808 _1004_/a_1059_315# _0217_ 0.01136f
C809 _0565_/a_51_297# comp0.B\[0\] 0.0061f
C810 clknet_1_0__leaf__0462_ _1007_/a_27_47# 0.04412f
C811 _1041_/a_193_47# hold5/a_391_47# 0
C812 net26 _0176_ 0.00575f
C813 _0290_ _0813_/a_109_297# 0.00289f
C814 acc0.A\[12\] _0282_ 0.05399f
C815 net61 _0263_ 0
C816 _1020_/a_466_413# net202 0
C817 net132 net11 0
C818 net57 _0725_/a_80_21# 0.00515f
C819 _0232_ _0754_/a_149_47# 0
C820 _0600_/a_337_297# _0219_ 0
C821 _0642_/a_27_413# output61/a_27_47# 0.00146f
C822 B[9] _0544_/a_512_297# 0
C823 _0231_ acc0.A\[24\] 0
C824 clknet_1_0__leaf__0465_ _1061_/a_891_413# 0
C825 acc0.A\[14\] _0635_/a_27_47# 0
C826 net56 _0334_ 0
C827 _1021_/a_466_413# _0119_ 0.04444f
C828 _0181_ _0507_/a_373_47# 0.00123f
C829 hold32/a_49_47# _0517_/a_299_297# 0
C830 hold32/a_285_47# _0517_/a_81_21# 0
C831 net31 _0545_/a_68_297# 0
C832 _1017_/a_1017_47# _0459_ 0
C833 clknet_1_0__leaf__0460_ _0969_/a_109_297# 0
C834 _0576_/a_109_47# _0380_ 0
C835 _0174_ _0536_/a_240_47# 0.01466f
C836 net125 _0144_ 0
C837 _0732_/a_209_297# _0368_ 0.00184f
C838 output66/a_27_47# _0512_/a_27_297# 0
C839 _0359_ hold90/a_49_47# 0.0437f
C840 _0510_/a_27_297# _0187_ 0.11063f
C841 _0996_/a_891_413# _0302_ 0
C842 clknet_1_1__leaf__0460_ _0698_/a_199_47# 0
C843 _1017_/a_27_47# _0218_ 0
C844 _1017_/a_193_47# _0294_ 0
C845 _1056_/a_381_47# acc0.A\[12\] 0
C846 hold23/a_285_47# acc0.A\[2\] 0
C847 net39 _0303_ 0
C848 _0461_ comp0.B\[15\] 0
C849 _1049_/a_891_413# clknet_1_1__leaf__0457_ 0
C850 _0690_/a_68_297# clknet_0__0462_ 0.00566f
C851 acc0.A\[20\] hold3/a_391_47# 0
C852 net62 _0988_/a_592_47# 0
C853 VPWR _0138_ 0.30255f
C854 _0211_ VPWR 0.30589f
C855 _0649_/a_113_47# net67 0
C856 hold12/a_49_47# _0468_ 0
C857 _0800_/a_51_297# net81 0.02049f
C858 _0751_/a_29_53# net241 0.08339f
C859 net57 _0128_ 0
C860 _0216_ net208 0.23029f
C861 _0467_ _1068_/a_193_47# 0
C862 _1050_/a_27_47# _0638_/a_109_297# 0
C863 acc0.A\[22\] _0224_ 0.01541f
C864 _0782_/a_27_47# _0112_ 0.01398f
C865 _0461_ _0773_/a_35_297# 0.00277f
C866 _0985_/a_27_47# _0985_/a_634_159# 0.14145f
C867 _0673_/a_337_297# _0288_ 0
C868 control0.count\[1\] _0978_/a_109_47# 0
C869 VPWR _0409_ 0.73938f
C870 _0986_/a_466_413# _0345_ 0
C871 hold19/a_285_47# _1017_/a_381_47# 0
C872 hold85/a_285_47# net232 0.01932f
C873 _0833_/a_215_47# _0253_ 0.00164f
C874 _0243_ hold64/a_285_47# 0
C875 control0.count\[2\] _1071_/a_891_413# 0.04689f
C876 _0535_/a_68_297# _1046_/a_27_47# 0
C877 _0642_/a_215_297# _0642_/a_298_297# 0.07178f
C878 _0173_ _0132_ 0.05368f
C879 hold47/a_285_47# _1050_/a_1059_315# 0.00813f
C880 hold47/a_49_47# _1050_/a_891_413# 0.002f
C881 _0348_ net44 0
C882 VPWR _1067_/a_1017_47# 0
C883 net82 _0094_ 0.01828f
C884 _0279_ _0284_ 0
C885 net176 _1022_/a_891_413# 0
C886 _0264_ _0219_ 0
C887 _1010_/a_27_47# acc0.A\[29\] 0
C888 _0313_ net237 0
C889 _0216_ _0612_/a_145_75# 0.00123f
C890 _0282_ _0650_/a_68_297# 0.12525f
C891 _0582_/a_109_47# net219 0
C892 _0582_/a_27_297# net206 0
C893 _0276_ _0345_ 0.09472f
C894 _1019_/a_193_47# _0459_ 0
C895 _0753_/a_79_21# _0753_/a_561_47# 0
C896 _0753_/a_297_297# _0753_/a_465_47# 0
C897 hold55/a_285_47# clknet_1_0__leaf__0461_ 0.004f
C898 clknet_1_1__leaf__0460_ _0691_/a_150_297# 0
C899 _0530_/a_81_21# _0530_/a_299_297# 0.08213f
C900 VPWR _0756_/a_47_47# 0.34182f
C901 _0187_ _0181_ 0.12375f
C902 _0172_ _0548_/a_245_297# 0
C903 _0734_/a_47_47# _0359_ 0
C904 hold27/a_285_47# clkbuf_0__0464_/a_110_47# 0
C905 VPWR _1027_/a_1059_315# 0.44437f
C906 _0218_ _0772_/a_215_47# 0
C907 _0586_/a_27_47# net223 0
C908 _1000_/a_1059_315# _0242_ 0
C909 _1003_/a_891_413# _0381_ 0
C910 _1003_/a_1059_315# _0237_ 0.00384f
C911 _0997_/a_27_47# _0408_ 0
C912 _0805_/a_181_47# _0283_ 0
C913 _0805_/a_109_47# _0286_ 0
C914 clknet_1_1__leaf__0462_ hold95/a_391_47# 0.00639f
C915 _1031_/a_193_47# _0704_/a_68_297# 0.00171f
C916 _1056_/a_27_47# acc0.A\[10\] 0.00364f
C917 _0181_ clknet_1_1__leaf__0461_ 0.0266f
C918 clk _0970_/a_285_47# 0
C919 _0153_ _0510_/a_109_297# 0
C920 hold61/a_391_47# net209 0
C921 net157 _1048_/a_975_413# 0
C922 _1042_/a_193_47# hold51/a_391_47# 0
C923 _0174_ _1046_/a_27_47# 0
C924 acc0.A\[25\] _1008_/a_27_47# 0
C925 _0165_ clknet_1_0__leaf__0461_ 0.09059f
C926 VPWR pp[31] 0.45733f
C927 _0460_ _0373_ 0.04633f
C928 _0247_ acc0.A\[18\] 0.05018f
C929 _0677_/a_47_47# _0677_/a_129_47# 0.00369f
C930 VPWR _0764_/a_384_47# 0
C931 _0546_/a_240_47# _1040_/a_634_159# 0
C932 _0546_/a_149_47# _1040_/a_466_413# 0
C933 _0399_ _1014_/a_466_413# 0
C934 _0743_/a_51_297# _0360_ 0.03512f
C935 _0487_ _1063_/a_27_47# 0.00376f
C936 _0342_ _0345_ 0.12216f
C937 _0341_ _0219_ 0.51091f
C938 _1019_/a_634_159# clknet_1_0__leaf__0461_ 0
C939 _0258_ _0824_/a_59_75# 0.04506f
C940 _1004_/a_466_413# _0379_ 0
C941 _0645_/a_285_47# acc0.A\[13\] 0.04452f
C942 acc0.A\[8\] _0989_/a_891_413# 0.02828f
C943 clknet_1_0__leaf__0464_ _0270_ 0.00742f
C944 _0144_ _0473_ 0
C945 _0346_ _0991_/a_466_413# 0.01908f
C946 _0974_/a_448_47# _0487_ 0.04121f
C947 _0600_/a_103_199# acc0.A\[23\] 0.00141f
C948 _0994_/a_193_47# net80 0.01442f
C949 _0996_/a_891_413# net6 0
C950 _0982_/a_27_47# _0218_ 0
C951 clknet_1_0__leaf__0464_ _0987_/a_466_413# 0
C952 hold48/a_285_47# net9 0
C953 hold88/a_285_47# _0988_/a_891_413# 0.00677f
C954 hold88/a_391_47# _0988_/a_1059_315# 0.00126f
C955 _0811_/a_81_21# hold70/a_285_47# 0.00102f
C956 hold64/a_49_47# clknet_1_0__leaf__0459_ 0
C957 _0345_ _0737_/a_285_47# 0.00296f
C958 _0361_ _0317_ 0.00193f
C959 hold15/a_285_47# VPWR 0.30286f
C960 hold7/a_285_47# net73 0.0026f
C961 hold7/a_49_47# _0085_ 0
C962 hold74/a_285_47# clkbuf_1_1__f__0461_/a_110_47# 0
C963 _0730_/a_79_21# _0352_ 0.11615f
C964 _0313_ _0686_/a_27_53# 0.00172f
C965 hold44/a_391_47# acc0.A\[27\] 0
C966 _0334_ _0345_ 0.03607f
C967 net28 net29 0
C968 _1034_/a_193_47# _1034_/a_592_47# 0.00135f
C969 _1034_/a_466_413# _1034_/a_561_413# 0.00772f
C970 _1034_/a_634_159# _1034_/a_975_413# 0
C971 hold6/a_49_47# _0544_/a_149_47# 0
C972 _0796_/a_510_47# _0410_ 0.00567f
C973 _0796_/a_297_297# _0094_ 0.00172f
C974 _0462_ _0771_/a_298_297# 0
C975 _0313_ _1008_/a_891_413# 0
C976 _0607_/a_109_297# _0308_ 0
C977 net168 _1053_/a_592_47# 0
C978 _0559_/a_512_297# net205 0
C979 comp0.B\[15\] _0465_ 0.0053f
C980 input25/a_75_212# input27/a_75_212# 0
C981 _0621_/a_285_297# _0434_ 0
C982 _0924_/a_27_47# net247 0.04744f
C983 _0464_ _0498_/a_240_47# 0
C984 _0257_ _0269_ 0
C985 pp[6] net58 0.10187f
C986 hold25/a_391_47# net30 0
C987 hold25/a_285_47# _0172_ 0.00216f
C988 _0729_/a_68_297# _0350_ 0.18445f
C989 _0640_/a_215_297# clknet_0__0465_ 0.00878f
C990 _0183_ net234 0.00618f
C991 _0399_ _0781_/a_150_297# 0
C992 control0.state\[0\] _1066_/a_381_47# 0
C993 _0570_/a_109_297# net197 0.00908f
C994 _0416_ _0284_ 0
C995 clknet_0__0464_ _1045_/a_466_413# 0.00113f
C996 _0853_/a_68_297# _0350_ 0
C997 _0224_ _0379_ 0
C998 _1063_/a_1017_47# _0161_ 0
C999 _0225_ _0378_ 0.54631f
C1000 _0086_ _0988_/a_891_413# 0
C1001 control0.state\[0\] _1068_/a_381_47# 0
C1002 control0.state\[0\] net1 0.11946f
C1003 _0842_/a_59_75# _0445_ 0
C1004 clknet_0__0458_ _0266_ 0.0011f
C1005 _0455_ acc0.A\[18\] 0
C1006 VPWR _1026_/a_561_413# 0.00314f
C1007 output59/a_27_47# net56 0
C1008 net219 net47 0
C1009 _0483_ _1072_/a_381_47# 0
C1010 control0.count\[3\] _1072_/a_975_413# 0.00189f
C1011 _0848_/a_109_297# _0450_ 0.01041f
C1012 _0848_/a_27_47# _0446_ 0.04535f
C1013 net215 _0216_ 0.07881f
C1014 _0183_ net46 0.02846f
C1015 output43/a_27_47# pp[14] 0
C1016 pp[16] output41/a_27_47# 0.01817f
C1017 VPWR _0817_/a_81_21# 0.55515f
C1018 _0547_/a_68_297# _0206_ 0.11908f
C1019 _0793_/a_51_297# net42 0.16046f
C1020 hold27/a_49_47# net147 0.05158f
C1021 _0218_ _0446_ 0.00589f
C1022 hold66/a_391_47# VPWR 0.21736f
C1023 pp[15] _1013_/a_193_47# 0
C1024 _0585_/a_373_47# _0112_ 0
C1025 hold64/a_49_47# _0453_ 0
C1026 net242 hold95/a_391_47# 0.13105f
C1027 _1018_/a_193_47# _0242_ 0
C1028 _1071_/a_193_47# _0488_ 0
C1029 _1071_/a_27_47# _0466_ 0.03987f
C1030 clknet_0__0465_ _0465_ 0.26116f
C1031 net135 acc0.A\[15\] 0
C1032 hold8/a_49_47# _0739_/a_79_21# 0
C1033 _0770_/a_79_21# _0248_ 0
C1034 _0993_/a_27_47# _0283_ 0
C1035 VPWR net134 0.39118f
C1036 hold8/a_285_47# _0347_ 0
C1037 _0959_/a_80_21# net25 0
C1038 _0855_/a_81_21# _0117_ 0.00317f
C1039 _0519_/a_384_47# _0437_ 0
C1040 acc0.A\[28\] clknet_1_1__leaf__0462_ 0.05254f
C1041 _1017_/a_634_159# _1017_/a_381_47# 0
C1042 _0487_ _1062_/a_1059_315# 0.06553f
C1043 _0357_ _0727_/a_193_47# 0
C1044 _0430_ _0346_ 0
C1045 clknet_1_1__leaf__0460_ hold50/a_391_47# 0
C1046 _0753_/a_297_297# _0234_ 0.00114f
C1047 _1052_/a_634_159# net9 0.02059f
C1048 _0644_/a_47_47# _0346_ 0.00453f
C1049 net56 _0724_/a_113_297# 0
C1050 clknet_1_1__leaf__0462_ net209 0
C1051 _0984_/a_466_413# _0219_ 0
C1052 _1016_/a_27_47# _1060_/a_193_47# 0
C1053 net248 _0255_ 0.02467f
C1054 _0500_/a_27_47# net9 0.00131f
C1055 net197 hold50/a_285_47# 0.0072f
C1056 _1006_/a_466_413# net52 0
C1057 _0507_/a_27_297# acc0.A\[13\] 0.06316f
C1058 _1000_/a_27_47# net45 0.13755f
C1059 _1000_/a_1059_315# net86 0
C1060 _1000_/a_466_413# _0098_ 0
C1061 _0223_ clknet_1_0__leaf__0460_ 0.03279f
C1062 _0430_ net65 0
C1063 _1060_/a_1017_47# _0158_ 0
C1064 _0958_/a_109_47# _0161_ 0
C1065 _1056_/a_466_413# hold34/a_49_47# 0
C1066 _1056_/a_193_47# hold34/a_391_47# 0
C1067 _0621_/a_35_297# _0252_ 0.00125f
C1068 _0129_ _1013_/a_1059_315# 0
C1069 _0363_ _1010_/a_27_47# 0
C1070 _0168_ _0169_ 0
C1071 control0.count\[1\] net164 0
C1072 _0346_ _0401_ 0.50192f
C1073 _0151_ _0186_ 0.00607f
C1074 acc0.A\[5\] _0346_ 0.00111f
C1075 hold46/a_391_47# _0200_ 0.05061f
C1076 net184 net154 0
C1077 VPWR _0084_ 0.2997f
C1078 _0959_/a_80_21# _0477_ 0.08801f
C1079 _0555_/a_51_297# _0174_ 0
C1080 _0210_ VPWR 1.09727f
C1081 _1033_/a_27_47# _1033_/a_634_159# 0.14092f
C1082 _0536_/a_240_47# _1046_/a_193_47# 0
C1083 output55/a_27_47# _0219_ 0.01693f
C1084 clknet_1_1__leaf__0458_ _0431_ 0.00174f
C1085 acc0.A\[5\] net65 0
C1086 _0463_ _0207_ 0
C1087 net55 _0734_/a_47_47# 0
C1088 _1012_/a_27_47# _1012_/a_634_159# 0.14145f
C1089 _0293_ _0817_/a_585_47# 0.00128f
C1090 _0331_ net57 0
C1091 hold96/a_391_47# net215 0
C1092 _0346_ net222 0.00115f
C1093 net211 _0247_ 0
C1094 _0401_ _0992_/a_466_413# 0
C1095 _0347_ _1007_/a_891_413# 0
C1096 _0352_ _1007_/a_634_159# 0
C1097 _1056_/a_193_47# _0510_/a_27_297# 0
C1098 _1056_/a_27_47# _0510_/a_109_297# 0
C1099 net158 hold36/a_391_47# 0
C1100 _0195_ _1031_/a_466_413# 0.03155f
C1101 _0216_ _1031_/a_193_47# 0.00235f
C1102 _0363_ _1009_/a_193_47# 0.00235f
C1103 hold66/a_391_47# net48 0
C1104 _0171_ clknet_1_1__leaf__0457_ 0
C1105 _0375_ _0374_ 0.0562f
C1106 control0.count\[3\] _0217_ 0.01659f
C1107 output55/a_27_47# _0728_/a_59_75# 0.0048f
C1108 _0476_ _0957_/a_32_297# 0.37434f
C1109 clkbuf_0__0458_/a_110_47# _0843_/a_68_297# 0.0135f
C1110 clkbuf_1_0__f__0457_/a_110_47# net211 0
C1111 clknet_0__0457_ _0579_/a_373_47# 0.0022f
C1112 hold27/a_49_47# net125 0.00228f
C1113 _0109_ _0700_/a_113_47# 0
C1114 _0161_ _0160_ 0.00344f
C1115 _0130_ _0457_ 0.01503f
C1116 _0637_/a_56_297# net47 0
C1117 net149 net223 0
C1118 _1072_/a_1059_315# clknet_0_clk 0.00284f
C1119 _1050_/a_193_47# _1050_/a_592_47# 0
C1120 _1050_/a_466_413# _1050_/a_561_413# 0.00772f
C1121 _1050_/a_634_159# _1050_/a_975_413# 0
C1122 hold27/a_391_47# _0953_/a_32_297# 0.00721f
C1123 hold59/a_285_47# _0454_ 0
C1124 hold59/a_49_47# _0455_ 0.01532f
C1125 _0990_/a_193_47# _0181_ 0.0349f
C1126 _0476_ net23 0.05314f
C1127 _0717_/a_80_21# acc0.A\[29\] 0
C1128 net36 _0854_/a_510_47# 0
C1129 _1041_/a_193_47# _0546_/a_51_297# 0
C1130 _1014_/a_193_47# _0345_ 0
C1131 clknet_1_0__leaf__0464_ _1051_/a_27_47# 0
C1132 _1024_/a_634_159# net50 0.00213f
C1133 _0179_ net135 0.00187f
C1134 net36 _0498_/a_51_297# 0
C1135 _0768_/a_109_297# _0462_ 0
C1136 hold29/a_285_47# _0122_ 0
C1137 _0428_ _0425_ 0
C1138 _0183_ _0996_/a_27_47# 0
C1139 _0339_ acc0.A\[29\] 0.0038f
C1140 _0465_ _0849_/a_215_47# 0
C1141 _0278_ _0218_ 0.1406f
C1142 _0565_/a_245_297# _0565_/a_240_47# 0
C1143 _0180_ _0527_/a_27_297# 0.1443f
C1144 net54 _0319_ 0.1893f
C1145 _0178_ _0208_ 0.45443f
C1146 _0680_/a_300_47# VPWR 0.00164f
C1147 net242 acc0.A\[28\] 0
C1148 _0595_/a_109_297# _0227_ 0.01129f
C1149 _0582_/a_109_297# _0774_/a_68_297# 0
C1150 _0998_/a_381_47# net43 0
C1151 _0662_/a_81_21# clknet_0__0465_ 0
C1152 _0218_ _0245_ 0.06677f
C1153 _1054_/a_466_413# _1052_/a_1059_315# 0
C1154 _0852_/a_285_47# _0399_ 0
C1155 pp[26] net156 0
C1156 _0409_ _0794_/a_110_297# 0.00193f
C1157 _0795_/a_81_21# _0300_ 0
C1158 _0982_/a_891_413# net149 0.00259f
C1159 _0176_ _1040_/a_466_413# 0.02829f
C1160 _1014_/a_193_47# hold2/a_49_47# 0
C1161 _1014_/a_27_47# hold2/a_285_47# 0
C1162 _0179_ _1054_/a_27_47# 0.01128f
C1163 net21 _1044_/a_27_47# 0.0218f
C1164 net183 _1044_/a_193_47# 0
C1165 _1056_/a_891_413# _0179_ 0.04957f
C1166 clkbuf_0__0465_/a_110_47# net72 0.00528f
C1167 _0748_/a_81_21# _0371_ 0
C1168 hold46/a_391_47# net193 0.15922f
C1169 _0995_/a_27_47# _0797_/a_27_413# 0.00106f
C1170 net25 _0173_ 0.00465f
C1171 _1056_/a_193_47# _0181_ 0
C1172 net205 _1036_/a_193_47# 0
C1173 _0973_/a_27_297# net240 0.11602f
C1174 _0555_/a_149_47# _0173_ 0.02212f
C1175 _0555_/a_51_297# _0208_ 0.18938f
C1176 _0236_ clknet_1_0__leaf__0457_ 0
C1177 _1024_/a_27_47# _1023_/a_27_47# 0.00164f
C1178 comp0.B\[13\] _1046_/a_27_47# 0
C1179 _0533_/a_109_47# _0465_ 0
C1180 hold10/a_49_47# _0199_ 0.00268f
C1181 hold10/a_391_47# net8 0
C1182 _0817_/a_266_47# clknet_1_1__leaf__0465_ 0
C1183 _0180_ _1061_/a_27_47# 0
C1184 _0343_ _1000_/a_592_47# 0
C1185 _0465_ hold71/a_285_47# 0.02245f
C1186 _1012_/a_193_47# clknet_1_1__leaf__0461_ 0.00205f
C1187 _1046_/a_27_47# _1046_/a_193_47# 0.96588f
C1188 hold86/a_49_47# hold100/a_285_47# 0.03505f
C1189 hold86/a_285_47# hold100/a_49_47# 0.03505f
C1190 _1058_/a_27_47# net66 0
C1191 clknet_1_1__leaf__0463_ input24/a_75_212# 0.00318f
C1192 _1050_/a_466_413# clkbuf_1_0__f__0464_/a_110_47# 0
C1193 _0772_/a_215_47# _0099_ 0.00256f
C1194 _0377_ _0103_ 0.00169f
C1195 net61 _0642_/a_27_413# 0
C1196 _0629_/a_59_75# _0182_ 0
C1197 _1054_/a_381_47# net12 0
C1198 _1016_/a_1059_315# net221 0.02842f
C1199 net204 _0473_ 0
C1200 net168 A[4] 0.05628f
C1201 _0752_/a_300_297# _0375_ 0.04187f
C1202 acc0.A\[2\] hold71/a_285_47# 0
C1203 net215 _1024_/a_193_47# 0.00589f
C1204 hold91/a_49_47# _0219_ 0
C1205 _0732_/a_209_297# _0732_/a_303_47# 0
C1206 net44 net43 0.14572f
C1207 _0724_/a_113_297# _0345_ 0.01247f
C1208 VPWR _0542_/a_149_47# 0.00483f
C1209 _0118_ net202 0.01525f
C1210 pp[8] A[11] 0.00425f
C1211 _0996_/a_27_47# acc0.A\[15\] 0.01268f
C1212 _0996_/a_193_47# net42 0
C1213 clkbuf_1_1__f__0463_/a_110_47# _0175_ 0.0943f
C1214 _0200_ net153 0
C1215 _0536_/a_240_47# comp0.B\[9\] 0
C1216 _1043_/a_27_47# net19 0
C1217 _1043_/a_193_47# net195 0.00607f
C1218 _1043_/a_466_413# _0203_ 0.00212f
C1219 _0211_ _1036_/a_27_47# 0
C1220 B[9] _0140_ 0
C1221 _0458_ _0186_ 0.33696f
C1222 clkbuf_1_0__f__0458_/a_110_47# hold75/a_391_47# 0.0061f
C1223 _0323_ clkbuf_0__0460_/a_110_47# 0.0553f
C1224 acc0.A\[12\] _1057_/a_27_47# 0.00334f
C1225 hold27/a_49_47# _0473_ 0
C1226 _1033_/a_891_413# net17 0.01093f
C1227 net63 _0518_/a_27_297# 0
C1228 _1019_/a_27_47# _0208_ 0
C1229 net44 _0999_/a_27_47# 0
C1230 _0246_ _0775_/a_79_21# 0
C1231 _1030_/a_466_413# _0333_ 0
C1232 _0206_ net127 0.00282f
C1233 comp0.B\[8\] net153 0
C1234 net129 net20 0
C1235 _1052_/a_193_47# _0522_/a_27_297# 0
C1236 _1052_/a_27_47# _0522_/a_109_297# 0
C1237 pp[26] acc0.A\[26\] 0
C1238 _0375_ _0249_ 0.01663f
C1239 _0761_/a_113_47# _0460_ 0
C1240 _0518_/a_109_297# net15 0.00919f
C1241 _0614_/a_183_297# _0246_ 0
C1242 hold86/a_391_47# _0446_ 0.00959f
C1243 _0856_/a_79_21# _0219_ 0
C1244 hold41/a_49_47# VPWR 0.29614f
C1245 hold100/a_285_47# acc0.A\[14\] 0.00113f
C1246 _0712_/a_465_47# _0195_ 0
C1247 _0985_/a_381_47# _0985_/a_561_413# 0.00123f
C1248 _0985_/a_891_413# _0985_/a_975_413# 0.00851f
C1249 _0504_/a_27_47# clknet_1_1__leaf__0457_ 0
C1250 _0217_ net176 0.28507f
C1251 clkbuf_1_0__f__0463_/a_110_47# _1040_/a_193_47# 0.00233f
C1252 _0688_/a_109_297# acc0.A\[25\] 0
C1253 net61 _0218_ 0.04303f
C1254 _0326_ _1007_/a_466_413# 0
C1255 net240 net17 0.01661f
C1256 _1018_/a_634_159# _1018_/a_592_47# 0
C1257 net36 _1014_/a_1059_315# 0
C1258 hold85/a_391_47# _0967_/a_215_297# 0
C1259 hold19/a_391_47# _1016_/a_193_47# 0.00107f
C1260 hold19/a_285_47# _1016_/a_634_159# 0
C1261 hold19/a_49_47# _1016_/a_466_413# 0.01453f
C1262 hold11/a_391_47# _0464_ 0
C1263 comp0.B\[14\] _1046_/a_891_413# 0.00437f
C1264 _0789_/a_75_199# _0409_ 0.02218f
C1265 _0404_ _0795_/a_81_21# 0.00538f
C1266 output58/a_27_47# _0642_/a_215_297# 0
C1267 _0195_ hold2/a_285_47# 0
C1268 _1021_/a_27_47# _1032_/a_27_47# 0
C1269 _0982_/a_634_159# _0982_/a_381_47# 0
C1270 net45 net165 0
C1271 _1011_/a_634_159# clknet_1_1__leaf__0462_ 0
C1272 _1049_/a_193_47# _1049_/a_381_47# 0.09799f
C1273 _1049_/a_634_159# _1049_/a_891_413# 0.03684f
C1274 _1049_/a_27_47# _1049_/a_561_413# 0.0027f
C1275 _0353_ _0335_ 0.01163f
C1276 _0983_/a_561_413# acc0.A\[15\] 0
C1277 _0349_ _0354_ 0
C1278 net12 _0522_/a_27_297# 0.01947f
C1279 net148 _0522_/a_373_47# 0
C1280 _0524_/a_27_297# net13 0
C1281 _0115_ net206 0
C1282 _0645_/a_47_47# _0303_ 0
C1283 _0172_ _0540_/a_240_47# 0.02343f
C1284 _0369_ _0345_ 0.69063f
C1285 _0462_ _0366_ 0
C1286 _0465_ _0529_/a_109_47# 0
C1287 _0305_ clknet_1_1__leaf__0465_ 0
C1288 clknet_0__0457_ _0345_ 0.05227f
C1289 _0467_ clkbuf_1_1__f_clk/a_110_47# 0.04516f
C1290 _0399_ _0841_/a_297_297# 0.00321f
C1291 _0397_ acc0.A\[17\] 0.0019f
C1292 _0413_ net6 0
C1293 comp0.B\[6\] net28 0.00549f
C1294 _1019_/a_634_159# _0218_ 0
C1295 hold56/a_391_47# _0133_ 0
C1296 hold98/a_285_47# net245 0.01139f
C1297 net193 net153 0
C1298 _0313_ _0320_ 0.05896f
C1299 hold16/a_285_47# _0195_ 0.02941f
C1300 _1066_/a_193_47# _1066_/a_381_47# 0.09972f
C1301 _1066_/a_634_159# _1066_/a_891_413# 0.03684f
C1302 _1066_/a_27_47# _1066_/a_561_413# 0.0027f
C1303 _0269_ clknet_1_1__leaf__0458_ 0.14942f
C1304 hold37/a_49_47# _1050_/a_1059_315# 0
C1305 net56 _1010_/a_381_47# 0
C1306 clknet_0__0459_ hold74/a_285_47# 0
C1307 _0343_ acc0.A\[17\] 0.00225f
C1308 net1 _1066_/a_193_47# 0
C1309 net45 acc0.A\[19\] 0.00405f
C1310 net89 _0382_ 0
C1311 net45 _0999_/a_561_413# 0
C1312 VPWR _1052_/a_975_413# 0.00477f
C1313 output64/a_27_47# _0253_ 0
C1314 _0852_/a_117_297# _0345_ 0
C1315 _0833_/a_79_21# net235 0.12013f
C1316 _1031_/a_381_47# acc0.A\[30\] 0
C1317 _1023_/a_466_413# _1022_/a_891_413# 0
C1318 _1068_/a_193_47# _1068_/a_381_47# 0.09799f
C1319 _1068_/a_634_159# _1068_/a_891_413# 0.03684f
C1320 _1068_/a_27_47# _1068_/a_561_413# 0.00163f
C1321 _0346_ hold70/a_49_47# 0.00815f
C1322 _0290_ _0809_/a_81_21# 0
C1323 net109 _0103_ 0
C1324 input1/a_27_47# net1 0.10965f
C1325 _1030_/a_27_47# _1030_/a_634_159# 0.13646f
C1326 _0557_/a_149_47# comp0.B\[4\] 0.00104f
C1327 _0217_ hold68/a_49_47# 0.00964f
C1328 net105 clknet_1_0__leaf__0461_ 0.2183f
C1329 _0294_ net219 0.0286f
C1330 VPWR net22 1.73304f
C1331 _0298_ net81 0
C1332 clkbuf_1_1__f_clk/a_110_47# comp0.B\[0\] 0.07463f
C1333 _1034_/a_193_47# clknet_1_1__leaf_clk 0
C1334 net49 net51 0
C1335 clkbuf_0__0460_/a_110_47# net237 0
C1336 net239 _0350_ 0.08095f
C1337 VPWR hold40/a_391_47# 0.18626f
C1338 _0415_ _0279_ 0.08979f
C1339 _1032_/a_381_47# net23 0.01048f
C1340 _0346_ _0089_ 0.66613f
C1341 _1035_/a_634_159# clknet_1_1__leaf__0463_ 0.00493f
C1342 _1035_/a_27_47# net122 0.00169f
C1343 _0992_/a_193_47# hold70/a_391_47# 0
C1344 _0992_/a_634_159# hold70/a_285_47# 0.00139f
C1345 clknet_1_0__leaf__0464_ _0085_ 0
C1346 VPWR net75 0.37914f
C1347 pp[27] _0221_ 0.04923f
C1348 hold53/a_285_47# _0123_ 0.00491f
C1349 comp0.B\[10\] hold5/a_391_47# 0.07195f
C1350 net198 net18 0.53844f
C1351 _0598_/a_79_21# _0598_/a_382_297# 0.00145f
C1352 _1015_/a_27_47# _0181_ 0.00844f
C1353 _0454_ _0219_ 0
C1354 _0718_/a_47_47# acc0.A\[29\] 0
C1355 net248 _0830_/a_215_47# 0
C1356 hold47/a_285_47# _1051_/a_193_47# 0
C1357 hold47/a_391_47# _1051_/a_27_47# 0
C1358 _0343_ net60 0.26456f
C1359 pp[8] net66 0.04811f
C1360 clknet_0__0458_ _0399_ 0.01605f
C1361 _0269_ _0263_ 0.13573f
C1362 _1051_/a_891_413# _0186_ 0.01795f
C1363 _1034_/a_1059_315# comp0.B\[2\] 0.13583f
C1364 _0765_/a_510_47# _0346_ 0
C1365 clkbuf_1_1__f__0458_/a_110_47# _0186_ 0.10596f
C1366 clknet_1_0__leaf__0463_ VPWR 3.42856f
C1367 _0343_ net5 0.08189f
C1368 _0125_ _1008_/a_27_47# 0
C1369 acc0.A\[27\] _1008_/a_466_413# 0.01691f
C1370 _0992_/a_27_47# net67 0.00111f
C1371 _1000_/a_27_47# VPWR 0.53865f
C1372 VPWR _0513_/a_299_297# 0.22953f
C1373 hold64/a_391_47# _0399_ 0
C1374 _1072_/a_634_159# _0466_ 0
C1375 _0254_ clknet_0__0465_ 0.06223f
C1376 net45 clkload3/a_268_47# 0
C1377 _0975_/a_59_75# clkbuf_1_0__f_clk/a_110_47# 0
C1378 net232 _0477_ 0.03032f
C1379 hold89/a_391_47# clkbuf_0_clk/a_110_47# 0
C1380 _0219_ _0505_/a_27_297# 0.04754f
C1381 _0100_ _0219_ 0
C1382 control0.state\[0\] control0.sh 0
C1383 clknet_0__0464_ net184 0.01001f
C1384 _0346_ _1006_/a_891_413# 0.0458f
C1385 comp0.B\[11\] _0545_/a_68_297# 0
C1386 _0247_ _0611_/a_150_297# 0
C1387 _0756_/a_129_47# net50 0.00383f
C1388 _0961_/a_113_297# _0478_ 0.03393f
C1389 net39 _0803_/a_68_297# 0.10065f
C1390 hold52/a_49_47# _0216_ 0.00788f
C1391 net168 hold21/a_285_47# 0.00853f
C1392 pp[30] _1031_/a_975_413# 0
C1393 _0407_ _0406_ 0.12514f
C1394 _0596_/a_59_75# clknet_1_0__leaf__0460_ 0.05207f
C1395 _0227_ _0606_/a_215_297# 0
C1396 _0686_/a_27_53# _0321_ 0
C1397 _0258_ _0432_ 0.26017f
C1398 _0973_/a_373_47# _0487_ 0.00305f
C1399 net175 _0530_/a_81_21# 0.06322f
C1400 _0343_ _0998_/a_634_159# 0.00253f
C1401 net138 VPWR 0.52372f
C1402 _0510_/a_27_297# clknet_1_1__leaf__0465_ 0
C1403 _0645_/a_47_47# _0996_/a_634_159# 0
C1404 _1017_/a_381_47# net103 0.02262f
C1405 _0467_ VPWR 1.48575f
C1406 acc0.A\[12\] _0672_/a_297_297# 0.00604f
C1407 hold13/a_285_47# net204 0
C1408 pp[28] _0327_ 0
C1409 _1017_/a_27_47# _1016_/a_1059_315# 0
C1410 _1017_/a_466_413# _1016_/a_193_47# 0.00297f
C1411 _1017_/a_193_47# _1016_/a_466_413# 0.00332f
C1412 _1017_/a_634_159# _1016_/a_634_159# 0
C1413 _0231_ _0375_ 0.53432f
C1414 _0661_/a_27_297# _0661_/a_205_297# 0.00412f
C1415 net178 _0516_/a_27_297# 0
C1416 _0280_ acc0.A\[14\] 0
C1417 _0822_/a_109_297# _0254_ 0.00174f
C1418 _0346_ _0616_/a_78_199# 0
C1419 _0998_/a_193_47# acc0.A\[17\] 0
C1420 _0578_/a_27_297# acc0.A\[20\] 0.00187f
C1421 input25/a_75_212# B[2] 0.19774f
C1422 _0849_/a_79_21# net47 0
C1423 output64/a_27_47# net74 0
C1424 _0506_/a_81_21# _0219_ 0
C1425 _0461_ acc0.A\[16\] 0
C1426 acc0.A\[13\] _0185_ 0
C1427 _0465_ _0986_/a_27_47# 0
C1428 _0555_/a_51_297# _0555_/a_245_297# 0.01218f
C1429 _0645_/a_285_47# VPWR 0
C1430 clkload0/a_27_47# _1071_/a_891_413# 0
C1431 _0733_/a_544_297# VPWR 0.01074f
C1432 _0415_ _0416_ 0.13354f
C1433 net85 clkbuf_1_1__f__0461_/a_110_47# 0.00131f
C1434 acc0.A\[30\] _0219_ 0.44802f
C1435 _0299_ _0797_/a_27_413# 0.10603f
C1436 hold47/a_49_47# clknet_1_0__leaf__0465_ 0.0035f
C1437 _0298_ _0797_/a_207_413# 0
C1438 _0476_ _0213_ 0.00289f
C1439 _0521_/a_384_47# _0151_ 0
C1440 _0248_ _0617_/a_68_297# 0.13363f
C1441 _1033_/a_891_413# _1033_/a_975_413# 0.00851f
C1442 _1033_/a_27_47# net119 0.26732f
C1443 _1033_/a_381_47# _1033_/a_561_413# 0.00123f
C1444 net149 clkbuf_0__0457_/a_110_47# 0.00104f
C1445 _0216_ _0329_ 0
C1446 net63 _0987_/a_27_47# 0.00425f
C1447 _0221_ _0724_/a_199_47# 0.01064f
C1448 VPWR comp0.B\[0\] 0.66614f
C1449 _1012_/a_891_413# _1012_/a_975_413# 0.00851f
C1450 _1012_/a_381_47# _1012_/a_561_413# 0.00123f
C1451 _1039_/a_381_47# _0176_ 0.01627f
C1452 VPWR _0780_/a_117_297# 0.00792f
C1453 _0130_ _1033_/a_193_47# 0.00282f
C1454 _1056_/a_1017_47# acc0.A\[10\] 0.00181f
C1455 _0545_/a_68_297# _0202_ 0
C1456 net58 _0264_ 0
C1457 _0344_ _0704_/a_68_297# 0
C1458 _0216_ clknet_1_0__leaf__0460_ 0.22939f
C1459 clknet_1_1__leaf__0460_ _0726_/a_245_297# 0
C1460 _0846_/a_240_47# _0345_ 0
C1461 _0846_/a_51_297# _0219_ 0.13692f
C1462 _0985_/a_193_47# _0636_/a_59_75# 0
C1463 _0529_/a_27_297# _0261_ 0.01322f
C1464 _0529_/a_109_297# _0262_ 0
C1465 hold79/a_391_47# _0162_ 0
C1466 _1056_/a_193_47# _0187_ 0
C1467 _0352_ net93 0.18164f
C1468 _0284_ net246 0
C1469 _0107_ _1009_/a_592_47# 0
C1470 _0805_/a_181_47# _0345_ 0
C1471 hold27/a_391_47# _0174_ 0.00702f
C1472 _1054_/a_27_47# hold83/a_49_47# 0.06616f
C1473 _1009_/a_466_413# _0219_ 0.01748f
C1474 _0181_ clknet_1_1__leaf__0465_ 0.38279f
C1475 hold86/a_391_47# net61 0
C1476 hold86/a_49_47# net233 0.00248f
C1477 _0220_ hold95/a_285_47# 0
C1478 _0259_ _0991_/a_466_413# 0
C1479 net44 _0677_/a_129_47# 0.00309f
C1480 _1050_/a_1059_315# acc0.A\[4\] 0.12817f
C1481 _0369_ net52 0
C1482 net15 _0987_/a_193_47# 0
C1483 clknet_1_1__leaf__0464_ hold51/a_391_47# 0
C1484 _1055_/a_891_413# acc0.A\[9\] 0.00762f
C1485 net178 _0399_ 0
C1486 _0257_ clkbuf_0__0458_/a_110_47# 0
C1487 _1041_/a_466_413# net152 0
C1488 pp[25] VPWR 0.26959f
C1489 net110 net50 0.21328f
C1490 _0854_/a_215_47# _0346_ 0
C1491 _0946_/a_30_53# _0484_ 0
C1492 _0216_ _0221_ 0.00849f
C1493 _0181_ _0215_ 0
C1494 _0163_ _0175_ 0
C1495 _1033_/a_891_413# _0165_ 0
C1496 _0350_ _0988_/a_891_413# 0
C1497 _0794_/a_27_47# acc0.A\[15\] 0
C1498 hold26/a_391_47# _0138_ 0
C1499 VPWR _0442_ 0.46042f
C1500 net161 net28 0
C1501 clkbuf_1_0__f__0463_/a_110_47# _0207_ 0.03093f
C1502 _0836_/a_68_297# _0369_ 0
C1503 net158 hold26/a_285_47# 0
C1504 _0476_ _0212_ 0.06275f
C1505 _0357_ _0350_ 0.05913f
C1506 VPWR _0544_/a_245_297# 0.00503f
C1507 _0983_/a_193_47# _1018_/a_634_159# 0
C1508 _0983_/a_27_47# _1018_/a_466_413# 0
C1509 hold96/a_285_47# net52 0.00905f
C1510 control0.state\[0\] _0483_ 0
C1511 _0294_ _0352_ 0.03321f
C1512 VPWR _1034_/a_634_159# 0.17968f
C1513 clknet_1_0__leaf__0460_ _1067_/a_27_47# 0.00138f
C1514 _0204_ _1043_/a_193_47# 0
C1515 _0369_ net212 0.13428f
C1516 _1004_/a_466_413# _0575_/a_27_297# 0
C1517 hold34/a_285_47# hold35/a_49_47# 0.00643f
C1518 hold34/a_49_47# hold35/a_285_47# 0.00643f
C1519 net58 net170 0
C1520 net169 _1052_/a_1059_315# 0.01079f
C1521 _0183_ _0902_/a_27_47# 0
C1522 _0465_ _0845_/a_193_297# 0
C1523 clknet_1_0__leaf__0458_ _0465_ 1.0493f
C1524 acc0.A\[14\] net103 0
C1525 VPWR _0374_ 0.71025f
C1526 hold6/a_285_47# _1043_/a_634_159# 0
C1527 hold6/a_49_47# _1043_/a_466_413# 0
C1528 _0176_ net174 0.22824f
C1529 _1053_/a_27_47# A[5] 0.00849f
C1530 _0998_/a_27_47# _0998_/a_466_413# 0.26005f
C1531 _0998_/a_193_47# _0998_/a_634_159# 0.12126f
C1532 hold32/a_49_47# VPWR 0.26229f
C1533 _0956_/a_114_297# _0208_ 0.00771f
C1534 _0337_ net208 0
C1535 clknet_1_0__leaf__0458_ acc0.A\[2\] 0.27667f
C1536 net64 _0988_/a_1059_315# 0.10597f
C1537 net45 _1018_/a_975_413# 0
C1538 net26 net28 0.00209f
C1539 _1059_/a_193_47# _0459_ 0.01099f
C1540 _1031_/a_975_413# _0339_ 0
C1541 hold96/a_391_47# clknet_1_0__leaf__0460_ 0.00116f
C1542 hold64/a_49_47# _0345_ 0
C1543 _0498_/a_51_297# _1061_/a_27_47# 0
C1544 _0796_/a_79_21# _0400_ 0.00526f
C1545 hold58/a_391_47# comp0.B\[4\] 0.07035f
C1546 net240 _0165_ 0.03401f
C1547 net85 _0998_/a_1059_315# 0
C1548 _0662_/a_81_21# _0986_/a_27_47# 0
C1549 _0769_/a_81_21# clknet_1_0__leaf__0461_ 0
C1550 net193 _1046_/a_592_47# 0
C1551 A[14] net5 0
C1552 _0574_/a_27_297# _0105_ 0.0012f
C1553 comp0.B\[1\] _0208_ 0.31903f
C1554 _0310_ _0776_/a_27_47# 0
C1555 hold87/a_49_47# clknet_1_0__leaf__0461_ 0.00157f
C1556 VPWR _0507_/a_27_297# 0.26358f
C1557 net118 _0584_/a_27_297# 0
C1558 _1001_/a_891_413# _0350_ 0.00913f
C1559 _1046_/a_466_413# _1046_/a_592_47# 0.00553f
C1560 _1046_/a_634_159# _1046_/a_1017_47# 0
C1561 _1019_/a_27_47# _1019_/a_193_47# 0.96965f
C1562 net233 acc0.A\[14\] 0
C1563 _0991_/a_381_47# _0263_ 0
C1564 _1019_/a_634_159# _0099_ 0.00176f
C1565 _1019_/a_891_413# net223 0
C1566 _0481_ _0162_ 0
C1567 _0227_ hold3/a_49_47# 0.00797f
C1568 acc0.A\[21\] hold3/a_285_47# 0.0772f
C1569 _1000_/a_27_47# clknet_1_0__leaf__0459_ 0.00387f
C1570 _0557_/a_240_47# _0549_/a_68_297# 0
C1571 _1056_/a_634_159# _0153_ 0
C1572 _0458_ net62 0
C1573 _0458_ _0450_ 0
C1574 _1032_/a_1017_47# clknet_1_0__leaf__0457_ 0
C1575 _1016_/a_1017_47# _0115_ 0
C1576 control0.state\[0\] control0.count\[1\] 0
C1577 VPWR _0317_ 0.42866f
C1578 net154 _0525_/a_299_297# 0.10014f
C1579 _1051_/a_891_413# _1050_/a_634_159# 0
C1580 _1051_/a_634_159# _1050_/a_891_413# 0
C1581 _1051_/a_1059_315# _1050_/a_466_413# 0
C1582 _1051_/a_466_413# _1050_/a_1059_315# 0
C1583 _1039_/a_1059_315# clkbuf_1_0__f__0463_/a_110_47# 0.01696f
C1584 _0716_/a_27_47# VPWR 0.43467f
C1585 _0949_/a_59_75# _1063_/a_27_47# 0
C1586 VPWR net165 1.75649f
C1587 _0218_ _0431_ 0.20098f
C1588 _0985_/a_381_47# net175 0
C1589 _0310_ _0219_ 0
C1590 _0462_ acc0.A\[24\] 0
C1591 _0982_/a_466_413# clkbuf_0__0457_/a_110_47# 0
C1592 _0559_/a_240_47# clknet_0__0463_ 0
C1593 _0452_ _0181_ 0.04964f
C1594 net45 clkbuf_1_1__f__0461_/a_110_47# 0.07307f
C1595 net196 _0203_ 0
C1596 _0556_/a_150_297# comp0.B\[4\] 0
C1597 net9 _1049_/a_27_47# 0.00622f
C1598 net175 _1049_/a_466_413# 0
C1599 _0217_ acc0.A\[18\] 0.0641f
C1600 _0133_ _0496_/a_27_47# 0
C1601 hold34/a_285_47# A[9] 0.00167f
C1602 hold87/a_285_47# net47 0.03086f
C1603 _0275_ _0840_/a_68_297# 0.04864f
C1604 _0259_ _0401_ 0.33686f
C1605 _0293_ _0816_/a_68_297# 0
C1606 _0576_/a_109_297# _0216_ 0
C1607 control0.sh _0565_/a_51_297# 0
C1608 _0775_/a_297_297# _0352_ 0
C1609 net48 _0374_ 0
C1610 net63 _0191_ 0.00236f
C1611 _0457_ _1032_/a_975_413# 0
C1612 _1041_/a_634_159# net10 0
C1613 control0.state\[1\] clkbuf_1_0__f_clk/a_110_47# 0
C1614 _0143_ _0180_ 0.03218f
C1615 _0279_ _0347_ 0.42113f
C1616 _1000_/a_1017_47# net46 0
C1617 clknet_0__0463_ net29 0
C1618 _0384_ _0346_ 0.02352f
C1619 _0758_/a_79_21# _0758_/a_215_47# 0.04584f
C1620 VPWR acc0.A\[19\] 1.25597f
C1621 _1024_/a_27_47# net52 0.00675f
C1622 VPWR _0999_/a_561_413# 0.00312f
C1623 _1052_/a_381_47# acc0.A\[6\] 0.00159f
C1624 _1052_/a_193_47# _0193_ 0
C1625 _0757_/a_68_297# net51 0.00154f
C1626 _0752_/a_300_297# VPWR 0.24266f
C1627 _0984_/a_1059_315# _0465_ 0.00207f
C1628 _0581_/a_109_297# net219 0.00164f
C1629 _0990_/a_27_47# _0990_/a_634_159# 0.13601f
C1630 clkbuf_0__0463_/a_110_47# _0213_ 0
C1631 _0289_ acc0.A\[13\] 0
C1632 _1039_/a_27_47# _0498_/a_51_297# 0
C1633 hold22/a_391_47# A[8] 0
C1634 _0534_/a_299_297# net149 0.06935f
C1635 _0733_/a_79_199# clkbuf_0__0462_/a_110_47# 0.01359f
C1636 _1039_/a_1017_47# net8 0
C1637 _0344_ _0216_ 0.00497f
C1638 _0985_/a_1017_47# _0083_ 0
C1639 _0984_/a_466_413# net58 0
C1640 hold27/a_49_47# comp0.B\[8\] 0
C1641 _0240_ _0394_ 0
C1642 _0326_ _0105_ 0.00234f
C1643 _0734_/a_285_47# _0350_ 0
C1644 _0369_ _0394_ 0
C1645 _0672_/a_79_21# acc0.A\[15\] 0.00253f
C1646 _0672_/a_297_297# net42 0
C1647 _0850_/a_150_297# _0350_ 0
C1648 _0343_ _0990_/a_561_413# 0
C1649 _0985_/a_1059_315# acc0.A\[3\] 0
C1650 _0463_ _0472_ 0.3782f
C1651 hold19/a_49_47# net166 0
C1652 hold56/a_49_47# _0132_ 0
C1653 _0346_ _1014_/a_466_413# 0.00199f
C1654 _0484_ _0487_ 0.09138f
C1655 _0343_ _0793_/a_245_297# 0
C1656 comp0.B\[10\] _0546_/a_51_297# 0.0146f
C1657 _0409_ _0345_ 0.02643f
C1658 _1053_/a_891_413# _0191_ 0
C1659 VPWR hold83/a_285_47# 0.29834f
C1660 _0982_/a_891_413# _0080_ 0
C1661 _0982_/a_381_47# net68 0
C1662 hold88/a_391_47# net235 0.13581f
C1663 net97 clknet_1_1__leaf__0462_ 0.00207f
C1664 _1049_/a_193_47# acc0.A\[3\] 0
C1665 _1049_/a_1059_315# _0147_ 0.04233f
C1666 _1049_/a_891_413# net135 0
C1667 net38 acc0.A\[11\] 0.31352f
C1668 hold25/a_285_47# _1040_/a_193_47# 0
C1669 hold25/a_49_47# _1040_/a_634_159# 0
C1670 hold25/a_391_47# _1040_/a_27_47# 0
C1671 _1011_/a_193_47# hold80/a_285_47# 0
C1672 _1011_/a_27_47# hold80/a_391_47# 0
C1673 clknet_0__0464_ _0176_ 0
C1674 net12 _0193_ 0.0293f
C1675 hold9/a_49_47# _0347_ 0
C1676 _0747_/a_215_47# _0371_ 0.00549f
C1677 _0747_/a_79_21# _0104_ 0.05052f
C1678 net248 _0989_/a_27_47# 0
C1679 _0237_ net159 0
C1680 _0949_/a_59_75# _1062_/a_1059_315# 0
C1681 VPWR _0249_ 0.60249f
C1682 _0551_/a_27_47# _0173_ 0
C1683 _1070_/a_193_47# _1070_/a_381_47# 0.10164f
C1684 _1070_/a_634_159# _1070_/a_891_413# 0.03684f
C1685 _1070_/a_27_47# _1070_/a_561_413# 0.0027f
C1686 clkbuf_1_0__f__0459_/a_110_47# acc0.A\[17\] 0
C1687 _1052_/a_27_47# _0150_ 0.1213f
C1688 _0172_ acc0.A\[15\] 0.28763f
C1689 _1053_/a_634_159# _1053_/a_592_47# 0
C1690 hold42/a_391_47# acc0.A\[10\] 0
C1691 pp[17] _1030_/a_27_47# 0.00252f
C1692 net44 _1030_/a_634_159# 0.0391f
C1693 _0575_/a_109_47# net199 0.00305f
C1694 hold98/a_285_47# VPWR 0.29389f
C1695 _0552_/a_68_297# control0.sh 0.00118f
C1696 net53 clkbuf_0__0462_/a_110_47# 0.00888f
C1697 clknet_1_0__leaf__0465_ _1050_/a_891_413# 0.00441f
C1698 _0532_/a_299_297# _0465_ 0.00209f
C1699 net45 _0998_/a_1059_315# 0.00837f
C1700 _0198_ _1061_/a_634_159# 0
C1701 _1032_/a_634_159# _0208_ 0
C1702 _1032_/a_891_413# _0173_ 0
C1703 _0183_ _1023_/a_193_47# 0
C1704 acc0.A\[22\] _1023_/a_634_159# 0.00281f
C1705 hold43/a_391_47# _0195_ 0.00845f
C1706 hold43/a_49_47# _0216_ 0.01153f
C1707 _1066_/a_891_413# clknet_1_1__leaf_clk 0
C1708 _1066_/a_193_47# control0.sh 0.01232f
C1709 _0179_ _0523_/a_299_297# 0.04802f
C1710 _0217_ hold59/a_49_47# 0.05199f
C1711 hold75/a_391_47# acc0.A\[15\] 0.00564f
C1712 _0314_ _1007_/a_891_413# 0.01599f
C1713 _0313_ _1007_/a_1059_315# 0
C1714 _0756_/a_47_47# _0345_ 0
C1715 _0082_ _0263_ 0
C1716 _0262_ net170 0
C1717 _0309_ _0777_/a_285_47# 0.03974f
C1718 hold10/a_391_47# _0492_/a_27_47# 0
C1719 acc0.A\[2\] _0532_/a_299_297# 0
C1720 net109 _1022_/a_381_47# 0.00141f
C1721 net177 _1022_/a_891_413# 0.00721f
C1722 net203 net185 0
C1723 _1068_/a_1059_315# _0166_ 0
C1724 clkbuf_1_1__f__0464_/a_110_47# _1044_/a_381_47# 0
C1725 _1030_/a_891_413# _1030_/a_975_413# 0.00851f
C1726 _1030_/a_381_47# _1030_/a_561_413# 0.00123f
C1727 clknet_0__0461_ clknet_1_0__leaf__0461_ 0.00411f
C1728 _0997_/a_27_47# net83 0.2243f
C1729 hold78/a_285_47# _0339_ 0.00585f
C1730 _1038_/a_466_413# _0552_/a_68_297# 0
C1731 _0476_ _0161_ 0
C1732 _0966_/a_27_47# _0975_/a_59_75# 0.00116f
C1733 _0461_ _0247_ 0.03774f
C1734 _0152_ net11 0
C1735 clknet_1_0__leaf__0462_ _0758_/a_215_47# 0
C1736 _0375_ _0225_ 0.05547f
C1737 _0330_ _0355_ 0
C1738 _0432_ net72 0.02437f
C1739 hold27/a_285_47# _1046_/a_634_159# 0
C1740 hold27/a_391_47# _1046_/a_193_47# 0
C1741 hold27/a_49_47# _1046_/a_466_413# 0
C1742 _0429_ _0152_ 0
C1743 _1014_/a_1059_315# hold60/a_391_47# 0.00126f
C1744 _1014_/a_891_413# hold60/a_285_47# 0.00677f
C1745 acc0.A\[14\] _0637_/a_311_297# 0.00151f
C1746 VPWR net197 0.30935f
C1747 clkbuf_1_0__f__0457_/a_110_47# _0461_ 0.00578f
C1748 net121 clknet_1_1__leaf__0463_ 0.35545f
C1749 _0233_ net46 0.35953f
C1750 _1056_/a_27_47# _1056_/a_634_159# 0.14145f
C1751 _0416_ _0347_ 0.01869f
C1752 _1032_/a_193_47# net17 0.01828f
C1753 _0389_ _0242_ 0.24272f
C1754 _0390_ acc0.A\[19\] 0.00246f
C1755 _0310_ _0746_/a_81_21# 0
C1756 _0229_ _0226_ 0.12977f
C1757 _0320_ _0321_ 0.00572f
C1758 output49/a_27_47# pp[21] 0.15655f
C1759 _0987_/a_634_159# _0987_/a_975_413# 0
C1760 _0987_/a_466_413# _0987_/a_561_413# 0.00772f
C1761 clknet_0__0459_ acc0.A\[13\] 0.19284f
C1762 clkbuf_1_0__f__0459_/a_110_47# net5 0.0047f
C1763 net194 _1051_/a_381_47# 0
C1764 net227 _0333_ 0
C1765 net211 _0217_ 0.1856f
C1766 pp[15] net81 0.00945f
C1767 _0312_ _0366_ 0
C1768 _0305_ _0398_ 0
C1769 _0290_ _0186_ 0
C1770 clknet_1_1__leaf__0459_ hold81/a_49_47# 0.01089f
C1771 _0855_/a_81_21# _0855_/a_384_47# 0.00138f
C1772 acc0.A\[1\] _1047_/a_1059_315# 0.10073f
C1773 _0182_ _1047_/a_466_413# 0.01305f
C1774 net1 clkbuf_1_1__f_clk/a_110_47# 0
C1775 _0608_/a_27_47# _0306_ 0.00704f
C1776 hold15/a_285_47# _0345_ 0
C1777 _1004_/a_27_47# _1004_/a_561_413# 0.0027f
C1778 _1004_/a_634_159# _1004_/a_891_413# 0.03684f
C1779 _1004_/a_193_47# _1004_/a_381_47# 0.09503f
C1780 _0729_/a_150_297# net57 0
C1781 _0195_ _0729_/a_68_297# 0.0015f
C1782 clknet_1_0__leaf__0459_ _0507_/a_27_297# 0.00876f
C1783 _1027_/a_193_47# _1008_/a_193_47# 0
C1784 _0094_ net41 0
C1785 pp[16] _0341_ 0.00172f
C1786 _0557_/a_240_47# _1035_/a_27_47# 0
C1787 _0557_/a_51_297# _1035_/a_1059_315# 0
C1788 clknet_0__0464_ net130 0.15955f
C1789 _0665_/a_109_297# acc0.A\[13\] 0
C1790 net157 _1049_/a_193_47# 0
C1791 acc0.A\[30\] hold61/a_49_47# 0.33062f
C1792 _0788_/a_150_297# _0399_ 0
C1793 _1021_/a_1059_315# _0382_ 0
C1794 hold18/a_49_47# _0465_ 0.01285f
C1795 _0528_/a_81_21# _0186_ 0
C1796 _0219_ _0184_ 0.05441f
C1797 _0179_ _0172_ 0.02202f
C1798 _0239_ _0219_ 0.00121f
C1799 _0447_ _0843_/a_68_297# 0.10534f
C1800 _0172_ B[14] 0
C1801 clknet_1_0__leaf__0465_ _1053_/a_27_47# 0.01301f
C1802 net63 clkbuf_1_0__f__0465_/a_110_47# 0.01779f
C1803 _1029_/a_193_47# _1029_/a_592_47# 0.00135f
C1804 _1029_/a_466_413# _1029_/a_561_413# 0.00772f
C1805 _1029_/a_634_159# _1029_/a_975_413# 0
C1806 acc0.A\[16\] _0582_/a_27_297# 0
C1807 clknet_1_0__leaf__0459_ net165 0
C1808 _0482_ net226 0.0013f
C1809 input24/a_75_212# input28/a_75_212# 0
C1810 _0577_/a_27_297# clknet_1_0__leaf__0460_ 0
C1811 _0390_ _0249_ 0
C1812 comp0.B\[11\] hold51/a_285_47# 0.02212f
C1813 _0254_ _0986_/a_27_47# 0
C1814 _0268_ _0446_ 0.09968f
C1815 acc0.A\[4\] _0256_ 0.01032f
C1816 _0343_ net84 0.00631f
C1817 _0817_/a_81_21# _0345_ 0.15491f
C1818 _0817_/a_81_21# _0814_/a_27_47# 0
C1819 _0187_ clknet_1_1__leaf__0465_ 0.66899f
C1820 _0462_ _0610_/a_59_75# 0.00317f
C1821 _0313_ clkbuf_1_0__f__0462_/a_110_47# 0.2287f
C1822 _0430_ _0253_ 0.03042f
C1823 hold67/a_285_47# clkbuf_1_1__f__0465_/a_110_47# 0
C1824 _0621_/a_285_47# _0253_ 0.00297f
C1825 comp0.B\[13\] _1045_/a_592_47# 0
C1826 acc0.A\[4\] _0987_/a_1059_315# 0.00482f
C1827 _0218_ _0269_ 0.27518f
C1828 _1015_/a_1059_315# _0565_/a_240_47# 0
C1829 _0716_/a_27_47# _0283_ 0.00196f
C1830 _0984_/a_193_47# _0263_ 0
C1831 _1004_/a_193_47# _0225_ 0
C1832 _1020_/a_27_47# net150 0
C1833 _1046_/a_891_413# _1045_/a_891_413# 0
C1834 clknet_1_0__leaf__0463_ net30 0.18569f
C1835 acc0.A\[29\] _0701_/a_303_47# 0
C1836 acc0.A\[1\] _0186_ 0
C1837 net178 _0190_ 0.24996f
C1838 _1017_/a_193_47# net166 0
C1839 net103 _1016_/a_634_159# 0.01689f
C1840 hold15/a_285_47# hold16/a_49_47# 0
C1841 _0661_/a_277_297# _0287_ 0.00106f
C1842 _0554_/a_150_297# comp0.B\[4\] 0
C1843 _0440_ acc0.A\[6\] 0
C1844 _0462_ _0691_/a_68_297# 0.00181f
C1845 clknet_1_0__leaf__0459_ acc0.A\[19\] 0.02957f
C1846 clknet_1_0__leaf__0462_ net108 0.28152f
C1847 _0856_/a_297_297# _0465_ 0.00105f
C1848 A[10] A[11] 0
C1849 _0275_ _0255_ 0
C1850 _0483_ _1068_/a_193_47# 0.00743f
C1851 control0.count\[3\] _1068_/a_466_413# 0
C1852 _0782_/a_27_47# _0182_ 0
C1853 hold81/a_285_47# hold81/a_391_47# 0.41909f
C1854 _1028_/a_1059_315# _1028_/a_891_413# 0.31086f
C1855 _1028_/a_193_47# _1028_/a_975_413# 0
C1856 _1028_/a_466_413# _1028_/a_381_47# 0.03733f
C1857 _0555_/a_149_47# net204 0.01083f
C1858 net63 input11/a_75_212# 0
C1859 _1030_/a_193_47# _0354_ 0
C1860 net58 _0856_/a_79_21# 0
C1861 _0343_ _0996_/a_634_159# 0.00144f
C1862 _0369_ _0989_/a_891_413# 0.00511f
C1863 net96 _0219_ 0
C1864 _0441_ _0835_/a_215_47# 0.00228f
C1865 _0453_ net165 0
C1866 _0812_/a_79_21# _0812_/a_297_297# 0.01735f
C1867 _0464_ clknet_1_1__leaf__0457_ 0.04146f
C1868 _0765_/a_297_297# clknet_1_0__leaf__0457_ 0
C1869 _0853_/a_68_297# _0852_/a_35_297# 0
C1870 _0238_ _0245_ 0
C1871 _0369_ _0992_/a_891_413# 0
C1872 hold57/a_391_47# _0549_/a_68_297# 0
C1873 _0985_/a_592_47# VPWR 0
C1874 hold27/a_391_47# comp0.B\[9\] 0
C1875 _0553_/a_149_47# _0176_ 0
C1876 _0174_ _0496_/a_27_47# 0
C1877 pp[30] hold61/a_391_47# 0.00719f
C1878 _0084_ _0345_ 0.02622f
C1879 _0483_ _0478_ 0.07747f
C1880 VPWR _1018_/a_975_413# 0.00436f
C1881 output45/a_27_47# net45 0.17206f
C1882 hold55/a_49_47# comp0.B\[1\] 0
C1883 _0351_ _0720_/a_68_297# 0.10687f
C1884 acc0.A\[11\] _0282_ 0
C1885 _0722_/a_510_47# net239 0
C1886 clknet_0__0463_ _0137_ 0.01748f
C1887 _0192_ clknet_1_0__leaf__0465_ 0.01689f
C1888 _0557_/a_51_297# _1037_/a_193_47# 0
C1889 VPWR _1049_/a_381_47# 0.07542f
C1890 _0802_/a_59_75# _0647_/a_285_47# 0
C1891 net149 _0350_ 0.29556f
C1892 _0581_/a_27_297# _0774_/a_68_297# 0.01998f
C1893 _0556_/a_68_297# input24/a_75_212# 0.00745f
C1894 _0231_ VPWR 0.58303f
C1895 _0812_/a_215_47# net228 0
C1896 _0263_ clkbuf_0__0458_/a_110_47# 0.01795f
C1897 _0796_/a_79_21# clkbuf_0__0459_/a_110_47# 0
C1898 _0575_/a_109_47# VPWR 0
C1899 _0202_ hold51/a_285_47# 0
C1900 _1041_/a_1059_315# net31 0.06081f
C1901 pp[15] _0797_/a_207_413# 0.00243f
C1902 _0460_ _1006_/a_193_47# 0.04143f
C1903 _0113_ comp0.B\[0\] 0
C1904 _0259_ _0089_ 0.00509f
C1905 hold97/a_49_47# _1008_/a_1059_315# 0.00791f
C1906 hold97/a_391_47# _1008_/a_634_159# 0
C1907 _0751_/a_111_297# _0460_ 0
C1908 VPWR _1066_/a_381_47# 0.09508f
C1909 _0490_ _1072_/a_27_47# 0
C1910 _0453_ acc0.A\[19\] 0
C1911 _1010_/a_27_47# clknet_1_1__leaf__0462_ 0
C1912 _0968_/a_193_297# _0488_ 0
C1913 VPWR _1068_/a_381_47# 0.06961f
C1914 VPWR net1 1.91898f
C1915 _0081_ _0853_/a_68_297# 0
C1916 _1053_/a_891_413# input11/a_75_212# 0.00342f
C1917 _0152_ clknet_1_1__leaf__0458_ 0.0016f
C1918 _0349_ _0353_ 0.00134f
C1919 _0218_ hold72/a_49_47# 0.08537f
C1920 _0315_ _0219_ 0.05269f
C1921 _0257_ net248 0.43471f
C1922 _0993_/a_381_47# _0417_ 0
C1923 _0993_/a_634_159# _0091_ 0.002f
C1924 VPWR clkbuf_1_1__f__0461_/a_110_47# 1.23151f
C1925 comp0.B\[14\] net184 0
C1926 A[7] A[8] 0
C1927 _0661_/a_109_297# clknet_1_1__leaf__0465_ 0
C1928 acc0.A\[17\] clkbuf_0__0461_/a_110_47# 0.0076f
C1929 _0769_/a_81_21# _0218_ 0
C1930 hold32/a_391_47# A[9] 0.05822f
C1931 net18 _1043_/a_592_47# 0.00131f
C1932 net198 _1043_/a_1017_47# 0
C1933 hold76/a_285_47# _0771_/a_298_297# 0
C1934 hold76/a_391_47# _0771_/a_215_297# 0
C1935 _0478_ control0.count\[1\] 0.00537f
C1936 clknet_1_0__leaf__0464_ net170 0.27541f
C1937 clknet_1_0__leaf__0465_ _1046_/a_381_47# 0.00194f
C1938 net103 _0116_ 0.00169f
C1939 hold87/a_49_47# _0218_ 0.01916f
C1940 _0343_ _0983_/a_592_47# 0
C1941 VPWR _0426_ 0.42879f
C1942 _1057_/a_381_47# _0181_ 0
C1943 net187 _0460_ 0
C1944 hold25/a_391_47# net171 0
C1945 hold25/a_285_47# _0207_ 0.0011f
C1946 _0996_/a_1059_315# acc0.A\[13\] 0
C1947 _0996_/a_193_47# net5 0.10913f
C1948 acc0.A\[21\] _0760_/a_285_47# 0.03054f
C1949 control0.sh _0493_/a_27_47# 0.12184f
C1950 _1019_/a_891_413# clkbuf_0__0457_/a_110_47# 0
C1951 _1002_/a_1017_47# acc0.A\[20\] 0
C1952 _0998_/a_193_47# net84 0.0535f
C1953 _0998_/a_1059_315# _0998_/a_1017_47# 0
C1954 _0710_/a_381_47# _0220_ 0
C1955 net45 _0793_/a_149_47# 0
C1956 _1020_/a_27_47# control0.add 0
C1957 _0430_ net74 0
C1958 clknet_1_0__leaf__0460_ _0756_/a_377_297# 0
C1959 net38 _0281_ 0
C1960 acc0.A\[12\] hold45/a_391_47# 0
C1961 _1003_/a_1017_47# _0369_ 0
C1962 _0101_ _0762_/a_215_47# 0
C1963 _0961_/a_113_297# VPWR 0.17936f
C1964 _0410_ _0408_ 0
C1965 net7 _1061_/a_193_47# 0.03057f
C1966 net150 _0219_ 0.00807f
C1967 _1024_/a_891_413# acc0.A\[23\] 0
C1968 net203 _1033_/a_634_159# 0
C1969 _0398_ _0181_ 0
C1970 clknet_0__0463_ comp0.B\[6\] 0.03906f
C1971 _0984_/a_634_159# net47 0.00739f
C1972 net190 _0569_/a_27_297# 0.0613f
C1973 control0.state\[1\] _0966_/a_27_47# 0
C1974 _0968_/a_109_297# net236 0
C1975 hold38/a_49_47# _0474_ 0
C1976 hold38/a_391_47# comp0.B\[6\] 0.01426f
C1977 VPWR _0185_ 0.32961f
C1978 _0174_ _1044_/a_975_413# 0
C1979 _0496_/a_27_47# _0208_ 0
C1980 _1019_/a_466_413# _1019_/a_592_47# 0.00553f
C1981 _1019_/a_634_159# _1019_/a_1017_47# 0
C1982 _0714_/a_51_297# _0714_/a_512_297# 0.0116f
C1983 _1058_/a_466_413# net37 0
C1984 net187 _0457_ 0
C1985 _0965_/a_47_47# _0965_/a_129_47# 0.00369f
C1986 hold42/a_391_47# _0188_ 0.03926f
C1987 net48 net1 0
C1988 _0467_ comp0.B\[3\] 0
C1989 net72 _0986_/a_381_47# 0
C1990 _0441_ _0172_ 0.07944f
C1991 VPWR _1012_/a_592_47# 0
C1992 _0730_/a_79_21# acc0.A\[27\] 0.03383f
C1993 _0172_ _0544_/a_51_297# 0.13487f
C1994 _0096_ _0307_ 0
C1995 _1051_/a_193_47# acc0.A\[4\] 0
C1996 _0149_ _1050_/a_1059_315# 0.00323f
C1997 _1030_/a_193_47# _0567_/a_27_297# 0
C1998 clk _0468_ 0.07843f
C1999 net173 _1040_/a_1059_315# 0
C2000 _0726_/a_245_297# _0726_/a_240_47# 0
C2001 acc0.A\[4\] _1045_/a_466_413# 0
C2002 pp[30] clknet_1_1__leaf__0462_ 0.04339f
C2003 _0183_ hold2/a_285_47# 0.00451f
C2004 _0291_ net62 0
C2005 hold9/a_391_47# net114 0
C2006 hold24/a_285_47# net171 0.04876f
C2007 _1058_/a_891_413# net67 0.00792f
C2008 hold24/a_49_47# _0207_ 0.00486f
C2009 _0535_/a_68_297# net152 0.00151f
C2010 _1033_/a_891_413# _1032_/a_1059_315# 0.01007f
C2011 _1033_/a_1059_315# _1032_/a_891_413# 0.01007f
C2012 _0346_ net229 0
C2013 net242 _1010_/a_27_47# 0
C2014 _0729_/a_68_297# _1010_/a_891_413# 0
C2015 A[10] net66 0.04415f
C2016 hold100/a_391_47# _0350_ 0.02174f
C2017 net175 _0147_ 0.2719f
C2018 _1013_/a_634_159# _0220_ 0
C2019 hold5/a_49_47# hold5/a_285_47# 0.22264f
C2020 _0326_ _0359_ 0.00818f
C2021 hold55/a_391_47# _1032_/a_27_47# 0
C2022 clknet_1_0__leaf__0465_ _0271_ 0.00407f
C2023 hold26/a_391_47# net22 0.04689f
C2024 _0536_/a_51_297# _0176_ 0
C2025 comp0.B\[3\] comp0.B\[0\] 0
C2026 VPWR _0998_/a_1059_315# 0.39441f
C2027 acc0.A\[29\] hold50/a_49_47# 0
C2028 clknet_1_0__leaf__0465_ _0987_/a_891_413# 0.00862f
C2029 _0347_ _0739_/a_79_21# 0.1471f
C2030 _0351_ net116 0
C2031 net208 _0333_ 0.00149f
C2032 _0990_/a_891_413# _0990_/a_975_413# 0.00851f
C2033 _0990_/a_381_47# _0990_/a_561_413# 0.00123f
C2034 hold81/a_285_47# _0281_ 0
C2035 clknet_1_0__leaf__0465_ A[5] 0.02002f
C2036 _1002_/a_891_413# _0460_ 0.01095f
C2037 _0294_ _0392_ 0.08967f
C2038 _1032_/a_193_47# _0165_ 0
C2039 _0174_ _0180_ 0.00162f
C2040 _0361_ _0462_ 0.02307f
C2041 _0793_/a_51_297# _0793_/a_245_297# 0.01218f
C2042 net16 acc0.A\[10\] 0
C2043 _0537_/a_150_297# _1043_/a_193_47# 0
C2044 _0343_ _0617_/a_68_297# 0.01369f
C2045 clknet_1_0__leaf__0463_ hold26/a_391_47# 0.00163f
C2046 _0172_ _0141_ 0.41545f
C2047 _0371_ _0352_ 0.16119f
C2048 _0174_ net152 0.66328f
C2049 _1050_/a_27_47# _0180_ 0.01694f
C2050 net61 _0268_ 0.05815f
C2051 _0518_/a_109_297# acc0.A\[5\] 0
C2052 hold86/a_391_47# _0269_ 0.01904f
C2053 _0967_/a_215_297# _0476_ 0.17744f
C2054 _0798_/a_113_297# _0405_ 0
C2055 _0770_/a_382_297# net46 0.00114f
C2056 hold55/a_285_47# _0721_/a_27_47# 0
C2057 _0466_ _0486_ 0.05678f
C2058 hold24/a_49_47# _1039_/a_1059_315# 0
C2059 _0312_ acc0.A\[24\] 0
C2060 net44 pp[17] 0.01256f
C2061 hold75/a_285_47# net165 0
C2062 net200 _1025_/a_634_159# 0.04161f
C2063 _0123_ _1025_/a_1059_315# 0.0131f
C2064 clknet_1_1__leaf__0463_ _1062_/a_1017_47# 0
C2065 _0124_ net113 0
C2066 clkload4/a_110_47# _0369_ 0
C2067 _1034_/a_27_47# comp0.B\[5\] 0
C2068 _0465_ _0846_/a_245_297# 0
C2069 _0832_/a_113_47# _0439_ 0.00937f
C2070 _1051_/a_27_47# _1051_/a_1059_315# 0.04875f
C2071 _1051_/a_193_47# _1051_/a_466_413# 0.07855f
C2072 hold9/a_391_47# _0365_ 0
C2073 hold9/a_49_47# _0106_ 0
C2074 _1056_/a_193_47# clknet_1_1__leaf__0465_ 0.00109f
C2075 VPWR _0832_/a_113_47# 0
C2076 _0742_/a_81_21# _0219_ 0.0065f
C2077 _0218_ clknet_0__0461_ 0.20411f
C2078 acc0.A\[14\] _0849_/a_297_297# 0
C2079 _0612_/a_59_75# _0242_ 0.03057f
C2080 net58 _0846_/a_51_297# 0
C2081 net106 _1033_/a_1059_315# 0
C2082 _1070_/a_1059_315# _0168_ 0
C2083 _1045_/a_634_159# _1045_/a_381_47# 0
C2084 _1070_/a_381_47# VPWR 0.07905f
C2085 _1070_/a_193_47# control0.count\[1\] 0.00113f
C2086 _1003_/a_27_47# hold66/a_285_47# 0
C2087 clknet_0__0458_ _0346_ 0.0115f
C2088 VPWR _1043_/a_193_47# 0.30605f
C2089 _0678_/a_68_297# _0306_ 0.01251f
C2090 _0217_ net177 0.09601f
C2091 acc0.A\[22\] net109 0.02634f
C2092 hold28/a_49_47# net170 0
C2093 hold23/a_285_47# acc0.A\[4\] 0
C2094 _0472_ clkbuf_1_0__f__0463_/a_110_47# 0
C2095 VPWR _1030_/a_592_47# 0
C2096 _1029_/a_27_47# _0106_ 0
C2097 _1043_/a_634_159# _1043_/a_381_47# 0
C2098 clknet_1_0__leaf__0459_ net1 0.04167f
C2099 hold46/a_49_47# _0176_ 0.00119f
C2100 clknet_1_1__leaf__0459_ _0654_/a_207_413# 0.02699f
C2101 hold20/a_49_47# _1005_/a_27_47# 0
C2102 _0554_/a_68_297# input24/a_75_212# 0
C2103 net82 acc0.A\[16\] 0
C2104 _0261_ _0449_ 0
C2105 _0309_ _0219_ 0.02536f
C2106 net236 _0486_ 0.05097f
C2107 clknet_1_0__leaf__0459_ clkbuf_1_1__f__0461_/a_110_47# 0
C2108 clknet_1_1__leaf__0460_ _0777_/a_47_47# 0
C2109 _1004_/a_381_47# VPWR 0.07961f
C2110 _0153_ A[9] 0.08019f
C2111 _1021_/a_1059_315# _1002_/a_1059_315# 0
C2112 hold89/a_391_47# _0487_ 0.05683f
C2113 _0518_/a_27_297# _0180_ 0.09966f
C2114 _1054_/a_27_47# _1054_/a_466_413# 0.27314f
C2115 _1054_/a_193_47# _1054_/a_634_159# 0.11105f
C2116 _0736_/a_139_47# clknet_1_1__leaf__0460_ 0
C2117 _1071_/a_634_159# clknet_1_0__leaf_clk 0
C2118 _0290_ net62 0
C2119 hold100/a_49_47# acc0.A\[1\] 0
C2120 _0983_/a_27_47# VPWR 0.40351f
C2121 acc0.A\[0\] hold60/a_49_47# 0.00295f
C2122 _0730_/a_79_21# _1010_/a_193_47# 0
C2123 _1056_/a_381_47# _1056_/a_561_413# 0.00123f
C2124 _0180_ _0208_ 0.03682f
C2125 _0982_/a_193_47# acc0.A\[1\] 0
C2126 _0339_ clknet_1_1__leaf__0462_ 0.00614f
C2127 comp0.B\[10\] _1042_/a_891_413# 0.00313f
C2128 output55/a_27_47# _0108_ 0
C2129 _0792_/a_209_297# _0792_/a_209_47# 0
C2130 _0792_/a_80_21# _0792_/a_303_47# 0.01146f
C2131 _0345_ hold40/a_391_47# 0
C2132 _0783_/a_79_21# clkbuf_1_1__f__0461_/a_110_47# 0.01349f
C2133 _0282_ _0281_ 0.0712f
C2134 _1038_/a_27_47# _1038_/a_193_47# 0.97371f
C2135 net194 acc0.A\[5\] 0
C2136 acc0.A\[9\] net47 0.00173f
C2137 net235 acc0.A\[8\] 0.1894f
C2138 net234 _0456_ 0.00401f
C2139 _0289_ VPWR 1.33042f
C2140 _0849_/a_510_47# _0451_ 0.00404f
C2141 net222 _0446_ 0.00169f
C2142 _0182_ _0145_ 0.24751f
C2143 _0476_ _0131_ 0
C2144 hold65/a_49_47# _0255_ 0
C2145 _1041_/a_1059_315# _0548_/a_240_47# 0
C2146 _0218_ _0082_ 0
C2147 _0972_/a_256_47# _0471_ 0.00361f
C2148 clknet_1_0__leaf__0459_ _0185_ 0
C2149 _0557_/a_245_297# _0133_ 0
C2150 _0557_/a_512_297# net121 0
C2151 _0727_/a_193_47# _0356_ 0
C2152 _0157_ _1060_/a_1059_315# 0
C2153 _1059_/a_1059_315# _0158_ 0
C2154 _0983_/a_193_47# _0983_/a_891_413# 0.19229f
C2155 _0983_/a_27_47# _0983_/a_381_47# 0.05761f
C2156 _0983_/a_634_159# _0983_/a_1059_315# 0
C2157 _0820_/a_79_21# hold67/a_391_47# 0
C2158 _0285_ net67 0.0018f
C2159 clknet_1_0__leaf__0465_ _1051_/a_634_159# 0.00364f
C2160 _0225_ VPWR 1.05921f
C2161 clknet_1_0__leaf__0465_ _1045_/a_1059_315# 0
C2162 _0758_/a_79_21# _0350_ 0.01375f
C2163 _0576_/a_27_297# net110 0.01974f
C2164 output45/a_27_47# VPWR 0.32185f
C2165 hold98/a_285_47# _0995_/a_634_159# 0.0135f
C2166 hold98/a_391_47# _0995_/a_193_47# 0.01053f
C2167 acc0.A\[16\] _0115_ 0
C2168 clkbuf_1_0__f__0461_/a_110_47# _0245_ 0.0048f
C2169 hold37/a_285_47# net131 0.01427f
C2170 hold37/a_49_47# net184 0
C2171 _0399_ _0507_/a_109_47# 0
C2172 net183 _0954_/a_32_297# 0
C2173 _0120_ clknet_1_0__leaf__0460_ 0
C2174 _0770_/a_297_47# VPWR 0.0058f
C2175 VPWR _0436_ 0.23459f
C2176 net55 hold95/a_391_47# 0
C2177 comp0.B\[13\] _1044_/a_975_413# 0
C2178 _0182_ _0446_ 0.00159f
C2179 comp0.B\[14\] _0176_ 0.13647f
C2180 _0422_ net143 0
C2181 _0437_ output63/a_27_47# 0.00149f
C2182 _0337_ _0221_ 0.00576f
C2183 _1015_/a_193_47# _0566_/a_27_47# 0.00103f
C2184 clknet_0__0463_ net26 0.00234f
C2185 _0606_/a_215_297# _0237_ 0
C2186 _1056_/a_27_47# hold35/a_49_47# 0
C2187 _1003_/a_634_159# _0217_ 0.00525f
C2188 _1003_/a_27_47# _0183_ 0
C2189 _0648_/a_27_297# _0276_ 0.20558f
C2190 _0956_/a_32_297# _0956_/a_304_297# 0.00167f
C2191 net162 _0129_ 0.48636f
C2192 acc0.A\[31\] net163 0
C2193 _1013_/a_466_413# _0218_ 0.00682f
C2194 _0317_ _0697_/a_80_21# 0.01839f
C2195 _1016_/a_634_159# _1016_/a_592_47# 0
C2196 net248 clknet_1_1__leaf__0458_ 0.02111f
C2197 _0251_ hold31/a_285_47# 0
C2198 net56 _0317_ 0
C2199 _0521_/a_81_21# _0180_ 0
C2200 pp[30] hold92/a_49_47# 0.01341f
C2201 net59 hold92/a_391_47# 0.13392f
C2202 control0.count\[3\] _0166_ 0
C2203 net242 _0339_ 0
C2204 clkbuf_0__0464_/a_110_47# net7 0
C2205 _0379_ net109 0
C2206 comp0.B\[1\] _0956_/a_220_297# 0.00805f
C2207 clknet_1_1__leaf__0462_ _1026_/a_193_47# 0.00845f
C2208 _1028_/a_466_413# acc0.A\[28\] 0
C2209 _0211_ net171 0
C2210 _0297_ acc0.A\[13\] 0.17029f
C2211 _1057_/a_381_47# _0187_ 0.01628f
C2212 _0399_ _0242_ 0
C2213 _0225_ net48 0.00224f
C2214 _0176_ _0543_/a_68_297# 0.13534f
C2215 _0173_ _0560_/a_150_297# 0
C2216 _0812_/a_215_47# _0090_ 0.00299f
C2217 VPWR _0990_/a_592_47# 0.001f
C2218 _0999_/a_592_47# _0399_ 0
C2219 _0327_ _0701_/a_80_21# 0.07939f
C2220 _0343_ _0725_/a_209_297# 0.00622f
C2221 input20/a_75_212# clknet_1_1__leaf__0464_ 0.0117f
C2222 hold97/a_49_47# clknet_1_1__leaf__0462_ 0
C2223 VPWR _0793_/a_149_47# 0.00327f
C2224 _1011_/a_27_47# _1029_/a_27_47# 0
C2225 _0749_/a_81_21# _0346_ 0.05204f
C2226 clkbuf_1_0__f__0462_/a_110_47# _0321_ 0.00126f
C2227 clknet_0__0459_ VPWR 2.60181f
C2228 _0397_ _0777_/a_129_47# 0.00341f
C2229 net64 net235 0
C2230 net39 _0994_/a_466_413# 0.03097f
C2231 clkbuf_0__0460_/a_110_47# clkbuf_1_0__f__0462_/a_110_47# 0.00125f
C2232 hold45/a_285_47# _0179_ 0.04047f
C2233 VPWR acc0.A\[3\] 1.63746f
C2234 _1032_/a_27_47# _0352_ 0
C2235 _1059_/a_1059_315# acc0.A\[14\] 0.06445f
C2236 _0584_/a_109_297# net157 0.0022f
C2237 _0116_ _0774_/a_68_297# 0.00141f
C2238 _0538_/a_51_297# net20 0.01348f
C2239 _1041_/a_1059_315# net7 0.05583f
C2240 _0211_ net24 0.0976f
C2241 _0403_ _0417_ 0
C2242 _1057_/a_27_47# acc0.A\[11\] 0
C2243 hold4/a_49_47# _1022_/a_891_413# 0
C2244 hold4/a_391_47# _1022_/a_466_413# 0
C2245 _0978_/a_27_297# clknet_1_0__leaf_clk 0
C2246 _0984_/a_193_47# _0218_ 0
C2247 net36 _0181_ 0.82516f
C2248 hold31/a_285_47# net58 0
C2249 VPWR control0.sh 2.09846f
C2250 _0198_ _1047_/a_1059_315# 0
C2251 _0146_ _1047_/a_193_47# 0
C2252 _1015_/a_27_47# _0215_ 0
C2253 _1056_/a_27_47# A[9] 0
C2254 comp0.B\[13\] net152 0
C2255 hold46/a_285_47# _0139_ 0.00182f
C2256 clknet_1_0__leaf__0462_ _0350_ 0.00514f
C2257 _0170_ _1072_/a_561_413# 0
C2258 _0665_/a_109_297# VPWR 0.00461f
C2259 _1056_/a_634_159# _1056_/a_1017_47# 0
C2260 hold29/a_49_47# hold29/a_391_47# 0.00188f
C2261 hold20/a_285_47# _0468_ 0
C2262 comp0.B\[14\] net130 0
C2263 _0398_ clknet_1_1__leaf__0461_ 0.06144f
C2264 _1054_/a_1059_315# VPWR 0.4014f
C2265 _0153_ _0516_/a_27_297# 0
C2266 _0305_ _0308_ 0.21469f
C2267 _0357_ _0195_ 0.04287f
C2268 _0358_ net57 0.0047f
C2269 acc0.A\[5\] _0987_/a_193_47# 0.00692f
C2270 _1051_/a_1059_315# _0085_ 0.01018f
C2271 _1051_/a_891_413# net73 0.00205f
C2272 clknet_1_0__leaf__0462_ _1025_/a_561_413# 0
C2273 net231 hold84/a_391_47# 0.1341f
C2274 hold34/a_391_47# _0515_/a_81_21# 0.00198f
C2275 clknet_1_1__leaf__0459_ _0286_ 0.14903f
C2276 _0770_/a_297_47# _0390_ 0
C2277 _0512_/a_109_297# net3 0.00625f
C2278 _1038_/a_466_413# VPWR 0.25652f
C2279 net154 _0524_/a_109_47# 0.00126f
C2280 _1041_/a_466_413# A[15] 0
C2281 net1 _0113_ 0.00232f
C2282 hold45/a_285_47# _0513_/a_81_21# 0
C2283 _0323_ _0368_ 0
C2284 VPWR _0655_/a_109_93# 0.08989f
C2285 _0767_/a_59_75# _0352_ 0
C2286 _1018_/a_891_413# acc0.A\[18\] 0.04296f
C2287 hold39/a_391_47# net23 0
C2288 _0183_ _0576_/a_373_47# 0.00196f
C2289 _0329_ _0319_ 0.32123f
C2290 hold74/a_391_47# _0219_ 0
C2291 net166 net219 0.00239f
C2292 _0131_ clkbuf_0__0463_/a_110_47# 0
C2293 clknet_0_clk _1068_/a_1017_47# 0
C2294 _0369_ clknet_1_0__leaf__0457_ 0.24209f
C2295 net120 _1065_/a_466_413# 0
C2296 _0983_/a_27_47# clknet_1_0__leaf__0459_ 0
C2297 clknet_0__0457_ clknet_1_0__leaf__0457_ 0.0325f
C2298 _0343_ acc0.A\[18\] 0.03295f
C2299 _0695_/a_80_21# _0250_ 0.14179f
C2300 _0627_/a_109_93# _0346_ 0.04548f
C2301 _0804_/a_79_21# _0276_ 0
C2302 _0374_ _0345_ 0.28447f
C2303 _0218_ clkbuf_0__0458_/a_110_47# 0.09666f
C2304 hold30/a_285_47# _0121_ 0.00407f
C2305 net247 net147 0
C2306 VPWR _0851_/a_113_47# 0
C2307 net44 _0567_/a_109_297# 0
C2308 _0369_ _0988_/a_1059_315# 0
C2309 net203 net119 0.21658f
C2310 VPWR _0418_ 0.20267f
C2311 VPWR _0785_/a_384_47# 0
C2312 net70 net47 0.0283f
C2313 _0430_ net61 0
C2314 _1019_/a_891_413# _0350_ 0
C2315 net190 _0127_ 0
C2316 _0842_/a_59_75# _0842_/a_145_75# 0.00658f
C2317 clknet_1_1__leaf__0459_ _0794_/a_27_47# 0
C2318 net145 _0218_ 0
C2319 _0157_ _0294_ 0
C2320 _0405_ net41 0.03711f
C2321 _1019_/a_1017_47# net105 0
C2322 _1031_/a_27_47# _1030_/a_27_47# 0
C2323 _0714_/a_51_297# _0111_ 0.10241f
C2324 _0817_/a_368_297# _0346_ 0.00226f
C2325 net35 _1071_/a_891_413# 0.0045f
C2326 _1008_/a_27_47# net244 0.00126f
C2327 net51 _1005_/a_592_47# 0
C2328 _0221_ _0319_ 0
C2329 _0325_ _0326_ 0.06116f
C2330 _0179_ _0437_ 0
C2331 net40 _0300_ 0
C2332 net245 _0297_ 0
C2333 net61 acc0.A\[5\] 0
C2334 _0180_ _0987_/a_27_47# 0
C2335 VPWR net157 0.98742f
C2336 _0237_ hold3/a_49_47# 0.06828f
C2337 _0381_ hold3/a_285_47# 0.0661f
C2338 _0343_ _0995_/a_891_413# 0.00111f
C2339 _1014_/a_381_47# clknet_1_0__leaf__0461_ 0.00291f
C2340 _1025_/a_27_47# _1025_/a_193_47# 0.97057f
C2341 _0726_/a_149_47# _0109_ 0
C2342 acc0.A\[4\] net184 0
C2343 _0668_/a_382_297# net6 0.00138f
C2344 _0339_ hold92/a_49_47# 0
C2345 _0479_ clkbuf_1_0__f_clk/a_110_47# 0.00205f
C2346 _0317_ _0345_ 0
C2347 net206 _0350_ 0.02728f
C2348 _0232_ net51 0.00377f
C2349 _0716_/a_27_47# _0345_ 0.01428f
C2350 net8 _0178_ 0
C2351 _0289_ _0283_ 0.22592f
C2352 control0.state\[2\] clknet_1_0__leaf__0460_ 0
C2353 _0343_ _0605_/a_109_297# 0
C2354 _0465_ _0448_ 0.00843f
C2355 _0800_/a_240_47# clknet_1_1__leaf__0459_ 0.00952f
C2356 net34 _1064_/a_381_47# 0.01649f
C2357 _1056_/a_592_47# acc0.A\[10\] 0.00143f
C2358 net165 _0345_ 0.03183f
C2359 clknet_1_0__leaf__0458_ net146 0.00172f
C2360 _1033_/a_381_47# clknet_1_1__leaf__0463_ 0
C2361 _0983_/a_27_47# _0453_ 0
C2362 net61 net222 0
C2363 B[7] A[1] 0.22703f
C2364 _1015_/a_466_413# net157 0.0011f
C2365 _0217_ _0461_ 0.03181f
C2366 hold58/a_49_47# _0133_ 0
C2367 _1050_/a_891_413# _0148_ 0
C2368 _0080_ _0350_ 0
C2369 net245 _0412_ 0.01406f
C2370 _1059_/a_634_159# net228 0
C2371 _0244_ _0393_ 0.05455f
C2372 _0739_/a_215_47# _0365_ 0.00735f
C2373 _0739_/a_79_21# _0106_ 0.05113f
C2374 acc0.A\[2\] _0448_ 0
C2375 _1046_/a_27_47# net10 0.44142f
C2376 clknet_0__0457_ _1001_/a_1059_315# 0
C2377 net77 net62 0.0024f
C2378 hold77/a_49_47# clknet_1_1__leaf__0461_ 0
C2379 _0515_/a_81_21# _0181_ 0
C2380 _0467_ _1065_/a_1059_315# 0.02098f
C2381 _0352_ _0365_ 0.07562f
C2382 _0119_ net187 0
C2383 _0089_ _0446_ 0
C2384 net77 _0450_ 0
C2385 hold95/a_49_47# hold95/a_285_47# 0.22264f
C2386 hold58/a_49_47# _0558_/a_68_297# 0
C2387 _0465_ _1048_/a_1017_47# 0
C2388 _0996_/a_27_47# _0996_/a_466_413# 0.27314f
C2389 _0996_/a_193_47# _0996_/a_634_159# 0.11072f
C2390 control0.count\[3\] _0168_ 0
C2391 _0483_ VPWR 0.92403f
C2392 acc0.A\[14\] _0264_ 0
C2393 _1054_/a_592_47# net9 0
C2394 _0238_ _0326_ 0
C2395 net67 _0218_ 0.07932f
C2396 _0555_/a_51_297# net8 0
C2397 _0174_ _0498_/a_51_297# 0.08607f
C2398 _0514_/a_373_47# net66 0
C2399 _0990_/a_1017_47# _0088_ 0
C2400 net36 _1018_/a_27_47# 0
C2401 _0473_ clknet_1_1__leaf__0464_ 0.00186f
C2402 _0386_ _0246_ 0
C2403 net125 net247 0.02654f
C2404 net152 comp0.B\[9\] 0
C2405 _0139_ net127 0
C2406 comp0.B\[3\] _1066_/a_381_47# 0
C2407 acc0.A\[19\] _0345_ 0.09186f
C2408 _0999_/a_466_413# _0219_ 0
C2409 _0793_/a_240_47# _0407_ 0.01246f
C2410 _0260_ _0261_ 0
C2411 _0646_/a_377_297# acc0.A\[13\] 0.00289f
C2412 acc0.A\[16\] _1017_/a_891_413# 0.02225f
C2413 _0234_ _0754_/a_149_47# 0.0021f
C2414 _0537_/a_68_297# net129 0.00181f
C2415 _1060_/a_466_413# _0505_/a_27_297# 0
C2416 hold55/a_285_47# _0182_ 0
C2417 _0195_ _0850_/a_150_297# 0
C2418 _0226_ _0382_ 0
C2419 acc0.A\[15\] _0301_ 0
C2420 _0559_/a_51_297# _0175_ 0.10947f
C2421 _0313_ _0324_ 0.32557f
C2422 net61 _0182_ 0.00134f
C2423 net237 _0368_ 0.17198f
C2424 VPWR _0996_/a_1059_315# 0.40143f
C2425 _0691_/a_150_297# _0219_ 0
C2426 _1065_/a_1059_315# comp0.B\[0\] 0.0133f
C2427 _0647_/a_285_47# _0414_ 0
C2428 _0698_/a_113_297# _1008_/a_466_413# 0
C2429 _0465_ _0444_ 0.00147f
C2430 comp0.B\[7\] _1039_/a_1017_47# 0
C2431 clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ 1.62938f
C2432 hold68/a_391_47# net199 0
C2433 net215 _0575_/a_373_47# 0
C2434 _1037_/a_381_47# net28 0
C2435 _1034_/a_1017_47# comp0.B\[6\] 0
C2436 clknet_1_0__leaf__0461_ _0771_/a_215_297# 0
C2437 hold33/a_391_47# _1041_/a_27_47# 0
C2438 _0331_ clkbuf_1_1__f__0462_/a_110_47# 0.11791f
C2439 _1051_/a_891_413# _1051_/a_1017_47# 0.00617f
C2440 _1051_/a_193_47# _0149_ 0.21099f
C2441 hold65/a_391_47# _0830_/a_79_21# 0
C2442 _1051_/a_634_159# net137 0
C2443 clknet_0__0459_ clknet_1_0__leaf__0459_ 0.21263f
C2444 _1045_/a_193_47# _1044_/a_381_47# 0
C2445 net247 _0635_/a_109_297# 0
C2446 net162 hold61/a_285_47# 0
C2447 _0992_/a_193_47# acc0.A\[10\] 0.07833f
C2448 _1051_/a_1059_315# net131 0
C2449 _0294_ acc0.A\[9\] 0.09812f
C2450 _0210_ net171 0
C2451 net160 _0207_ 0.00263f
C2452 net62 _0986_/a_1059_315# 0.14242f
C2453 VPWR control0.count\[1\] 0.81746f
C2454 _1045_/a_381_47# net131 0
C2455 _1045_/a_891_413# net184 0
C2456 clkbuf_1_0__f__0464_/a_110_47# net170 0.01283f
C2457 net78 net217 0.15846f
C2458 net23 _1067_/a_381_47# 0.01918f
C2459 _1003_/a_891_413# net213 0
C2460 net61 _0443_ 0.00344f
C2461 _1072_/a_1059_315# clknet_1_0__leaf_clk 0
C2462 _0399_ _0990_/a_27_47# 0.42673f
C2463 _0249_ _0345_ 0
C2464 _0643_/a_337_297# _0465_ 0
C2465 _1028_/a_592_47# _0350_ 0
C2466 clknet_1_1__leaf__0464_ _0186_ 0.03933f
C2467 _1002_/a_193_47# net240 0.00178f
C2468 clknet_1_1__leaf__0459_ _0673_/a_103_199# 0
C2469 _0984_/a_466_413# _0158_ 0
C2470 _0227_ _0223_ 0
C2471 _1043_/a_381_47# net129 0
C2472 _1043_/a_891_413# net196 0
C2473 _1060_/a_634_159# _0506_/a_299_297# 0
C2474 VPWR _0568_/a_373_47# 0
C2475 VPWR _1015_/a_975_413# 0.0048f
C2476 hold49/a_49_47# clknet_1_1__leaf__0464_ 0.01395f
C2477 clknet_1_1__leaf__0459_ _0672_/a_79_21# 0.0021f
C2478 clknet_0__0459_ _0283_ 0
C2479 _0195_ hold19/a_391_47# 0
C2480 _0181_ _0308_ 0.00579f
C2481 clknet_1_1__leaf__0460_ _0743_/a_240_47# 0
C2482 _0788_/a_150_297# _0346_ 0
C2483 _0458_ _0529_/a_27_297# 0.00896f
C2484 _0361_ _0312_ 0
C2485 _0594_/a_113_47# net150 0
C2486 _0210_ net24 0.5277f
C2487 _0628_/a_109_297# _0186_ 0.00158f
C2488 _0479_ control0.count\[2\] 0.11999f
C2489 clknet_1_0__leaf__0463_ _1040_/a_27_47# 0.02653f
C2490 control0.state\[1\] hold84/a_391_47# 0
C2491 hold3/a_49_47# _1005_/a_27_47# 0
C2492 net58 output47/a_27_47# 0.00101f
C2493 _0984_/a_193_47# hold86/a_391_47# 0
C2494 pp[25] net52 0
C2495 _1021_/a_381_47# net88 0.00676f
C2496 _0233_ _0601_/a_68_297# 0.11124f
C2497 _1032_/a_634_159# _1032_/a_466_413# 0.23992f
C2498 _1032_/a_193_47# _1032_/a_1059_315# 0.03405f
C2499 _1032_/a_27_47# _1032_/a_891_413# 0.03224f
C2500 _0191_ _0180_ 0.13401f
C2501 _1054_/a_27_47# net169 0.10769f
C2502 _1054_/a_193_47# net140 0.01516f
C2503 _1054_/a_1059_315# _1054_/a_1017_47# 0
C2504 _0568_/a_27_297# _0568_/a_109_297# 0.17136f
C2505 _1015_/a_634_159# _1015_/a_592_47# 0
C2506 _0712_/a_79_21# _1030_/a_27_47# 0
C2507 _0717_/a_80_21# hold80/a_49_47# 0
C2508 _1038_/a_27_47# net29 0.0049f
C2509 _0748_/a_299_297# _0369_ 0.00453f
C2510 net78 _0744_/a_27_47# 0
C2511 _0824_/a_59_75# _0824_/a_145_75# 0.00658f
C2512 _0991_/a_891_413# _0347_ 0
C2513 _0557_/a_240_47# _0173_ 0.01223f
C2514 _0357_ _1010_/a_891_413# 0
C2515 _0108_ _1010_/a_634_159# 0.00197f
C2516 _0439_ pp[4] 0
C2517 _0753_/a_79_21# clknet_1_0__leaf__0460_ 0.0136f
C2518 clknet_1_1__leaf__0462_ _1027_/a_592_47# 0
C2519 _0335_ hold80/a_391_47# 0
C2520 VPWR pp[4] 0.58089f
C2521 _0252_ output63/a_27_47# 0.0099f
C2522 _1056_/a_27_47# _0399_ 0
C2523 _0234_ _0228_ 0.00599f
C2524 _0376_ _0605_/a_109_297# 0
C2525 _0989_/a_193_47# pp[5] 0
C2526 _0343_ _1031_/a_891_413# 0.00106f
C2527 _1014_/a_27_47# net149 0.05963f
C2528 _0216_ clknet_0__0462_ 0
C2529 VPWR _0550_/a_240_47# 0.00407f
C2530 _0217_ _0465_ 0.00217f
C2531 net247 _1047_/a_1059_315# 0
C2532 _1038_/a_466_413# _1038_/a_592_47# 0.00553f
C2533 _1038_/a_634_159# _1038_/a_1017_47# 0
C2534 _1039_/a_1059_315# net160 0
C2535 _0211_ _1037_/a_466_413# 0
C2536 _0855_/a_81_21# _0399_ 0
C2537 _0442_ _0836_/a_68_297# 0.11268f
C2538 _0172_ _1043_/a_27_47# 0.00797f
C2539 _1067_/a_1059_315# clknet_1_0__leaf__0461_ 0.0056f
C2540 _0461_ _0248_ 0
C2541 hold19/a_285_47# _0369_ 0.00198f
C2542 _0655_/a_215_53# _0286_ 0.00195f
C2543 _0655_/a_109_93# _0283_ 0.1266f
C2544 net40 _0646_/a_285_47# 0.07106f
C2545 net59 _0336_ 0.00186f
C2546 _0134_ net121 0.00203f
C2547 clknet_1_0__leaf__0465_ _1044_/a_466_413# 0.00145f
C2548 _0983_/a_1059_315# net69 0
C2549 clknet_1_0__leaf__0465_ net137 0.01329f
C2550 net154 _0142_ 0.06086f
C2551 _1011_/a_193_47# _0347_ 0
C2552 clkbuf_1_1__f__0465_/a_110_47# _0990_/a_891_413# 0
C2553 _0661_/a_27_297# _0295_ 0
C2554 _1034_/a_891_413# net33 0
C2555 hold86/a_391_47# clkbuf_0__0458_/a_110_47# 0
C2556 _0102_ _0380_ 0
C2557 _0263_ _0447_ 0
C2558 net40 _0995_/a_592_47# 0
C2559 _0245_ _1006_/a_891_413# 0
C2560 _0283_ _0418_ 0
C2561 _0172_ _0171_ 0.00522f
C2562 _0659_/a_150_297# _0291_ 0
C2563 _0143_ comp0.B\[12\] 0
C2564 output62/a_27_47# pp[4] 0.33841f
C2565 hold64/a_49_47# clknet_1_0__leaf__0457_ 0.0099f
C2566 _0550_/a_51_297# _0550_/a_149_47# 0.02487f
C2567 _0997_/a_466_413# net42 0.03125f
C2568 _0230_ _0600_/a_337_297# 0.00758f
C2569 _0116_ hold72/a_391_47# 0
C2570 net106 _1032_/a_27_47# 0.00661f
C2571 _0229_ _0765_/a_79_21# 0
C2572 _0466_ _1068_/a_975_413# 0.00109f
C2573 acc0.A\[12\] _1058_/a_193_47# 0.02569f
C2574 _1031_/a_1059_315# net60 0
C2575 _0268_ _0269_ 0.3227f
C2576 _0851_/a_113_47# _0453_ 0.00954f
C2577 net89 _0217_ 0
C2578 _0101_ net150 0.02042f
C2579 _0280_ _0276_ 0.12495f
C2580 _1054_/a_634_159# acc0.A\[6\] 0.00203f
C2581 _0117_ hold60/a_285_47# 0.00107f
C2582 _0316_ _0313_ 0.00157f
C2583 _0330_ _0322_ 0.00374f
C2584 clknet_1_0__leaf__0462_ _1005_/a_1059_315# 0.00219f
C2585 VPWR _0955_/a_32_297# 0.39677f
C2586 _0553_/a_149_47# net28 0
C2587 _0244_ net206 0.00657f
C2588 _1061_/a_1059_315# acc0.A\[15\] 0.1292f
C2589 hold31/a_391_47# _0254_ 0
C2590 clknet_0__0459_ _0996_/a_1017_47# 0
C2591 net158 net147 0
C2592 _0330_ _0327_ 0.04845f
C2593 clknet_0__0458_ _0259_ 0.00514f
C2594 _0534_/a_299_297# hold71/a_285_47# 0
C2595 _0998_/a_381_47# _0399_ 0.00869f
C2596 _0998_/a_891_413# _0096_ 0.00415f
C2597 net84 _0783_/a_215_47# 0
C2598 _0313_ _0347_ 0
C2599 _0329_ _0333_ 0.02517f
C2600 hold22/a_285_47# VPWR 0.27975f
C2601 hold11/a_391_47# clknet_1_0__leaf__0464_ 0
C2602 clknet_0__0465_ net66 0.03576f
C2603 acc0.A\[10\] net142 0
C2604 _0186_ _0825_/a_68_297# 0.02341f
C2605 _1036_/a_27_47# control0.sh 0
C2606 _0356_ _0350_ 0
C2607 _0773_/a_35_297# _0773_/a_285_297# 0.02504f
C2608 hold68/a_391_47# VPWR 0.18194f
C2609 _0490_ _0467_ 0
C2610 net150 hold4/a_285_47# 0
C2611 _0217_ hold4/a_49_47# 0.03883f
C2612 acc0.A\[20\] _0749_/a_299_297# 0
C2613 _0328_ _1026_/a_466_413# 0
C2614 _1008_/a_634_159# hold50/a_391_47# 0.00158f
C2615 _1008_/a_466_413# hold50/a_285_47# 0
C2616 _1052_/a_634_159# net11 0.00179f
C2617 _1052_/a_891_413# net154 0
C2618 VPWR _0462_ 1.66398f
C2619 _0195_ net149 0.55386f
C2620 _0645_/a_129_47# _0301_ 0
C2621 _0982_/a_27_47# _1014_/a_466_413# 0.00287f
C2622 _0985_/a_891_413# _0219_ 0
C2623 _0195_ _1017_/a_466_413# 0.02358f
C2624 hold64/a_49_47# _1001_/a_1059_315# 0
C2625 clk _0978_/a_109_297# 0.00111f
C2626 hold48/a_391_47# net21 0
C2627 hold4/a_391_47# net151 0.14562f
C2628 net70 _0294_ 0
C2629 acc0.A\[0\] _0263_ 0
C2630 hold39/a_285_47# _0173_ 0.04048f
C2631 hold39/a_391_47# _0213_ 0.01847f
C2632 net55 _0702_/a_113_47# 0
C2633 hold42/a_49_47# VPWR 0.25594f
C2634 _0677_/a_47_47# _0306_ 0.0015f
C2635 hold17/a_391_47# clkbuf_1_0__f_clk/a_110_47# 0
C2636 _0752_/a_384_47# clknet_1_0__leaf__0460_ 0
C2637 _1057_/a_466_413# VPWR 0.24415f
C2638 _1048_/a_466_413# _0186_ 0
C2639 _0221_ _0333_ 1.14936f
C2640 _0732_/a_80_21# clknet_1_0__leaf__0460_ 0
C2641 hold24/a_285_47# _0135_ 0
C2642 hold29/a_49_47# net50 0.0575f
C2643 clkbuf_1_1__f__0462_/a_110_47# _1008_/a_27_47# 0
C2644 _0231_ _0345_ 0
C2645 _0343_ net241 0
C2646 _0647_/a_285_47# _0404_ 0
C2647 _0241_ _0216_ 0.04398f
C2648 _0464_ net135 0.1632f
C2649 _0179_ _0252_ 0.15464f
C2650 _0179_ _0989_/a_381_47# 0
C2651 _0275_ _0257_ 0
C2652 _0272_ _0258_ 0
C2653 net44 _0399_ 0
C2654 _0362_ _1009_/a_27_47# 0
C2655 _0153_ _0190_ 0.07956f
C2656 _0222_ _0606_/a_215_297# 0
C2657 _0249_ net52 0
C2658 net1 _0345_ 0
C2659 acc0.A\[12\] _0787_/a_80_21# 0
C2660 _0647_/a_47_47# _0304_ 0
C2661 _0315_ _1007_/a_193_47# 0
C2662 _0367_ _1007_/a_27_47# 0
C2663 _0366_ _1007_/a_634_159# 0.0569f
C2664 _0971_/a_299_297# control0.reset 0
C2665 clkbuf_1_1__f__0459_/a_110_47# _0277_ 0.0098f
C2666 net172 VPWR 0.30128f
C2667 hold5/a_285_47# net152 0.00969f
C2668 hold5/a_49_47# net32 0
C2669 _0338_ _0220_ 0.24669f
C2670 _0335_ _0336_ 0
C2671 net45 hold59/a_391_47# 0
C2672 net64 pp[6] 0.08048f
C2673 _0343_ output42/a_27_47# 0.06466f
C2674 _0805_/a_27_47# _0402_ 0.225f
C2675 hold69/a_49_47# hold69/a_285_47# 0.22264f
C2676 _0522_/a_27_297# _0522_/a_109_47# 0.00393f
C2677 net118 clknet_1_0__leaf__0460_ 0
C2678 net117 _0352_ 0
C2679 _0989_/a_891_413# net75 0
C2680 _0179_ _1061_/a_1059_315# 0
C2681 _1001_/a_27_47# _0580_/a_27_297# 0
C2682 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# 1.66421f
C2683 _0323_ clknet_0__0460_ 0.3652f
C2684 net35 _1072_/a_561_413# 0
C2685 _1067_/a_975_413# _0460_ 0
C2686 _1067_/a_1017_47# clknet_1_0__leaf__0457_ 0
C2687 _0690_/a_68_297# _0364_ 0
C2688 net78 _0350_ 0
C2689 _0401_ _0659_/a_68_297# 0.0014f
C2690 _1017_/a_634_159# _0369_ 0.01832f
C2691 _0225_ _1023_/a_27_47# 0
C2692 clknet_0__0465_ _0350_ 0.09186f
C2693 _0152_ net15 0
C2694 net44 _1031_/a_27_47# 0
C2695 clknet_1_0__leaf__0460_ _0250_ 0.20634f
C2696 _0426_ _0345_ 0.16053f
C2697 _0672_/a_297_297# _0303_ 0
C2698 _0607_/a_109_47# _0347_ 0
C2699 _0432_ clkbuf_1_0__f__0465_/a_110_47# 0.02957f
C2700 _0426_ _0814_/a_27_47# 0.00782f
C2701 _1059_/a_891_413# net41 0
C2702 _0965_/a_377_297# _0488_ 0
C2703 _0965_/a_47_47# _0466_ 0.04017f
C2704 hold100/a_391_47# hold18/a_391_47# 0.00216f
C2705 net48 _0462_ 0.05039f
C2706 _0275_ _0818_/a_109_47# 0
C2707 _1020_/a_381_47# net118 0.00119f
C2708 _0760_/a_129_47# _0237_ 0.00164f
C2709 _0760_/a_47_47# _0382_ 0.14737f
C2710 _0760_/a_285_47# _0381_ 0.07042f
C2711 _0428_ _0181_ 0.35855f
C2712 net178 _0988_/a_634_159# 0.04005f
C2713 _0217_ _0582_/a_27_297# 0.10556f
C2714 net248 _0218_ 0.12026f
C2715 _0982_/a_1059_315# hold18/a_285_47# 0
C2716 _0982_/a_891_413# hold18/a_49_47# 0
C2717 _0815_/a_113_297# _0991_/a_193_47# 0
C2718 _1053_/a_1059_315# _0152_ 0
C2719 _1012_/a_27_47# _0306_ 0
C2720 _1012_/a_193_47# _0308_ 0
C2721 _0983_/a_634_159# _0399_ 0.03727f
C2722 net225 _0111_ 0.13548f
C2723 output51/a_27_47# _1022_/a_1059_315# 0
C2724 net51 _1022_/a_193_47# 0.00473f
C2725 net150 net23 0
C2726 net133 _0159_ 0
C2727 _0981_/a_109_297# _0478_ 0
C2728 _0181_ hold60/a_391_47# 0
C2729 hold58/a_49_47# _0208_ 0
C2730 VPWR _0297_ 0.63663f
C2731 _0328_ _0315_ 0.02555f
C2732 net36 _0531_/a_27_297# 0
C2733 clknet_1_0__leaf__0463_ _1061_/a_466_413# 0.00184f
C2734 acc0.A\[21\] _0384_ 0
C2735 hold21/a_285_47# acc0.A\[8\] 0
C2736 _0185_ _0345_ 0
C2737 net247 _0497_/a_68_297# 0.00369f
C2738 _1038_/a_1059_315# net180 0
C2739 _1038_/a_27_47# _0137_ 0
C2740 _1038_/a_466_413# net30 0
C2741 clknet_1_0__leaf__0463_ net171 0.00139f
C2742 _0712_/a_561_47# net60 0
C2743 hold7/a_285_47# _0194_ 0
C2744 net160 _1037_/a_1059_315# 0.00292f
C2745 acc0.A\[0\] clknet_1_0__leaf__0461_ 0.04299f
C2746 _1025_/a_466_413# _1025_/a_592_47# 0.00553f
C2747 _1025_/a_634_159# _1025_/a_1017_47# 0
C2748 acc0.A\[13\] _0669_/a_183_297# 0
C2749 _1012_/a_592_47# _0345_ 0
C2750 _0390_ _0462_ 0.00123f
C2751 _0764_/a_81_21# _0460_ 0.00307f
C2752 _0984_/a_27_47# _0347_ 0
C2753 comp0.B\[1\] net202 0
C2754 hold25/a_49_47# _0136_ 0.29021f
C2755 _0369_ _0973_/a_109_47# 0
C2756 comp0.B\[1\] clknet_1_1__leaf__0463_ 0
C2757 net69 _0266_ 0
C2758 _0113_ net157 0
C2759 VPWR net13 0.69246f
C2760 _0247_ net223 0
C2761 _1070_/a_592_47# _0488_ 0
C2762 control0.count\[1\] _0976_/a_535_374# 0
C2763 clkbuf_0_clk/a_110_47# _0972_/a_250_297# 0
C2764 _0412_ VPWR 0.35864f
C2765 net236 _0965_/a_47_47# 0
C2766 net145 net228 0
C2767 _0955_/a_304_297# _0215_ 0
C2768 comp0.B\[6\] _0564_/a_150_297# 0
C2769 clknet_1_1__leaf__0459_ net79 0.14732f
C2770 clknet_1_1__leaf__0459_ _0808_/a_585_47# 0
C2771 clknet_1_0__leaf__0463_ net24 0
C2772 clknet_0__0463_ _0465_ 0.00219f
C2773 hold17/a_391_47# control0.count\[2\] 0.04972f
C2774 _0403_ _0994_/a_891_413# 0
C2775 net150 net35 0
C2776 hold86/a_285_47# _0449_ 0.00228f
C2777 _0116_ _0264_ 0
C2778 acc0.A\[14\] _0670_/a_297_297# 0
C2779 clkload4/a_268_47# acc0.A\[15\] 0
C2780 hold18/a_285_47# _0451_ 0
C2781 _0539_/a_68_297# net19 0.00298f
C2782 _0996_/a_1059_315# _0996_/a_1017_47# 0
C2783 _1055_/a_891_413# _0517_/a_299_297# 0
C2784 _0715_/a_27_47# _0181_ 0.01297f
C2785 _0998_/a_27_47# _0219_ 0
C2786 _0443_ _0431_ 0.10956f
C2787 hold57/a_391_47# _0173_ 0.05484f
C2788 _0388_ _0352_ 0.1541f
C2789 _0314_ _1025_/a_193_47# 0
C2790 hold5/a_49_47# net10 0.00911f
C2791 A[8] net11 0
C2792 clkload2/a_110_47# clknet_1_0__leaf__0465_ 0
C2793 _0218_ _0771_/a_215_297# 0
C2794 _0753_/a_561_47# acc0.A\[23\] 0
C2795 _0849_/a_215_47# _0350_ 0.00858f
C2796 net99 _0220_ 0
C2797 comp0.B\[3\] control0.sh 0.00864f
C2798 net158 _0473_ 0
C2799 comp0.B\[1\] net8 0
C2800 _0159_ comp0.B\[10\] 0
C2801 _0518_/a_373_47# _0369_ 0
C2802 _0298_ clkbuf_1_1__f__0459_/a_110_47# 0
C2803 _0376_ net241 0
C2804 _0158_ _0505_/a_27_297# 0.0122f
C2805 net146 _0505_/a_109_297# 0.00374f
C2806 _1060_/a_466_413# _0184_ 0
C2807 _1060_/a_891_413# net6 0
C2808 acc0.A\[16\] _1016_/a_193_47# 0.02088f
C2809 _0559_/a_149_47# _0559_/a_240_47# 0.06872f
C2810 _0701_/a_303_47# clknet_1_1__leaf__0462_ 0
C2811 clknet_1_0__leaf__0463_ _1039_/a_466_413# 0
C2812 _1057_/a_381_47# clknet_1_1__leaf__0465_ 0.01248f
C2813 net58 clknet_1_1__leaf__0457_ 0
C2814 VPWR _1036_/a_891_413# 0.19241f
C2815 A[13] output40/a_27_47# 0.00541f
C2816 net237 clknet_0__0460_ 0
C2817 clknet_0__0457_ _0982_/a_634_159# 0
C2818 clknet_1_1__leaf__0461_ _0308_ 0.03826f
C2819 _1044_/a_634_159# _1044_/a_1059_315# 0
C2820 _1044_/a_27_47# _1044_/a_381_47# 0.06222f
C2821 _1044_/a_193_47# _1044_/a_891_413# 0.19489f
C2822 _0596_/a_145_75# acc0.A\[21\] 0
C2823 _0596_/a_59_75# _0227_ 0.04176f
C2824 net227 acc0.A\[29\] 0.23925f
C2825 _0296_ clkbuf_1_1__f__0459_/a_110_47# 0.00626f
C2826 _0274_ _0640_/a_465_297# 0
C2827 hold46/a_285_47# _0954_/a_32_297# 0
C2828 _1038_/a_27_47# comp0.B\[6\] 0.00351f
C2829 _0815_/a_113_297# _0423_ 0.00758f
C2830 _0174_ A[15] 0
C2831 _1056_/a_27_47# _0190_ 0
C2832 _1051_/a_592_47# acc0.A\[5\] 0
C2833 net131 _1044_/a_891_413# 0
C2834 _0222_ hold3/a_49_47# 0
C2835 clknet_0__0458_ _0253_ 0.02272f
C2836 hold59/a_285_47# net234 0
C2837 clknet_1_0__leaf__0462_ _0592_/a_68_297# 0.00449f
C2838 net67 net228 0.13624f
C2839 _0386_ _0774_/a_68_297# 0
C2840 _0580_/a_109_297# clknet_1_0__leaf__0461_ 0.00415f
C2841 _0753_/a_79_21# hold94/a_285_47# 0
C2842 clk _0480_ 0.0084f
C2843 _0358_ clkbuf_1_1__f__0460_/a_110_47# 0.00413f
C2844 net23 control0.add 0
C2845 net46 _1023_/a_1059_315# 0.04204f
C2846 _0699_/a_68_297# net227 0
C2847 _1067_/a_193_47# net17 0.0356f
C2848 output66/a_27_47# acc0.A\[10\] 0
C2849 hold56/a_391_47# clknet_1_1__leaf__0463_ 0.01075f
C2850 _1051_/a_1059_315# net170 0
C2851 _1051_/a_891_413# _0196_ 0
C2852 _1057_/a_27_47# _1057_/a_193_47# 0.96543f
C2853 _0259_ _0627_/a_109_93# 0
C2854 VPWR _0754_/a_245_297# 0.00558f
C2855 _1039_/a_381_47# clknet_0__0463_ 0.00136f
C2856 _0324_ _0321_ 0.03477f
C2857 hold54/a_285_47# net106 0
C2858 _0158_ _0506_/a_81_21# 0.12289f
C2859 _0552_/a_68_297# _0549_/a_68_297# 0.01117f
C2860 _0231_ net52 0
C2861 _0839_/a_109_297# clknet_0__0465_ 0
C2862 clkbuf_0__0460_/a_110_47# _0324_ 0.00205f
C2863 _1059_/a_27_47# _1059_/a_193_47# 0.9735f
C2864 _0575_/a_27_297# pp[24] 0
C2865 _0575_/a_109_47# net52 0.00103f
C2866 _1003_/a_1017_47# _0467_ 0
C2867 B[6] net29 0.00532f
C2868 acc0.A\[14\] _0454_ 0
C2869 clknet_0__0464_ _0142_ 0.49293f
C2870 net166 hold72/a_285_47# 0
C2871 _1030_/a_592_47# _0345_ 0
C2872 acc0.A\[4\] _0525_/a_299_297# 0
C2873 _0662_/a_81_21# _0424_ 0.01116f
C2874 hold100/a_49_47# net247 0
C2875 acc0.A\[12\] pp[9] 0
C2876 _0500_/a_27_47# _1047_/a_27_47# 0.00897f
C2877 _0310_ _0775_/a_79_21# 0
C2878 _1032_/a_634_159# net202 0
C2879 _0430_ _0269_ 0
C2880 _0568_/a_109_297# _0128_ 0.00169f
C2881 _0146_ _0178_ 0
C2882 _1032_/a_634_159# clknet_1_1__leaf__0463_ 0
C2883 _0569_/a_109_297# acc0.A\[29\] 0.0219f
C2884 _0108_ net96 0.00108f
C2885 _0374_ hold94/a_391_47# 0.07467f
C2886 net9 net71 0
C2887 _0179_ _1058_/a_27_47# 0
C2888 _0487_ net91 0
C2889 acc0.A\[14\] _0505_/a_27_297# 0.12279f
C2890 _0820_/a_215_47# _0990_/a_1059_315# 0
C2891 hold46/a_391_47# _0540_/a_51_297# 0
C2892 _1014_/a_381_47# _0112_ 0.11469f
C2893 _0244_ _0773_/a_35_297# 0.04409f
C2894 _0210_ _0553_/a_51_297# 0
C2895 _0218_ _0339_ 0.00633f
C2896 _0310_ _0614_/a_183_297# 0
C2897 _0679_/a_68_297# _0245_ 0
C2898 _0211_ _0135_ 0
C2899 _0783_/a_215_47# _0783_/a_510_47# 0.00529f
C2900 _1038_/a_592_47# net172 0
C2901 hold39/a_391_47# _0161_ 0
C2902 _0223_ _0352_ 0.19787f
C2903 net33 _1066_/a_592_47# 0.00258f
C2904 net193 clknet_1_1__leaf__0464_ 0.00269f
C2905 _0573_/a_27_47# net149 0.02367f
C2906 hold44/a_391_47# VPWR 0.18842f
C2907 _0328_ _0689_/a_150_297# 0
C2908 _0765_/a_215_47# _0352_ 0.04233f
C2909 net55 net97 0
C2910 _0427_ _0816_/a_68_297# 0
C2911 hold86/a_49_47# _0846_/a_51_297# 0
C2912 _0343_ _1055_/a_466_413# 0
C2913 acc0.A\[27\] _1028_/a_634_159# 0.00516f
C2914 comp0.B\[14\] _0954_/a_114_297# 0.00249f
C2915 _0646_/a_377_297# VPWR 0.00381f
C2916 hold25/a_391_47# _0206_ 0
C2917 _0289_ _0345_ 0.09029f
C2918 clknet_0__0463_ net174 0
C2919 _0289_ _0814_/a_27_47# 0.00667f
C2920 _0292_ _0814_/a_109_47# 0
C2921 _0268_ _0082_ 0.00209f
C2922 _0269_ net222 0
C2923 control0.count\[2\] _0976_/a_218_47# 0
C2924 input30/a_75_212# clkbuf_1_0__f__0463_/a_110_47# 0
C2925 acc0.A\[20\] hold73/a_49_47# 0.00633f
C2926 _0274_ _0988_/a_27_47# 0
C2927 hold27/a_391_47# net10 0
C2928 _0129_ _1030_/a_1059_315# 0
C2929 _1020_/a_561_413# net1 0
C2930 net163 _1030_/a_634_159# 0
C2931 _0293_ _0295_ 0
C2932 _0287_ _0304_ 0.00836f
C2933 net168 _1052_/a_1059_315# 0.00304f
C2934 _0140_ hold51/a_391_47# 0
C2935 _0267_ _0841_/a_510_47# 0
C2936 _0352_ _1006_/a_1059_315# 0.01588f
C2937 acc0.A\[21\] _0383_ 0.0261f
C2938 _0570_/a_27_297# clknet_1_1__leaf__0462_ 0.0183f
C2939 VPWR _0995_/a_561_413# 0.00318f
C2940 _0284_ _0993_/a_1059_315# 0.00118f
C2941 net101 _1015_/a_193_47# 0.00358f
C2942 _0641_/a_113_47# _0437_ 0
C2943 _0769_/a_81_21# clkbuf_1_0__f__0461_/a_110_47# 0.00176f
C2944 _0343_ _0799_/a_80_21# 0.13135f
C2945 _0346_ _0242_ 0
C2946 net23 net231 0
C2947 clkbuf_1_1__f__0464_/a_110_47# net148 0
C2948 hold78/a_49_47# net45 0.00758f
C2949 net247 _0450_ 0
C2950 _0225_ _0345_ 0.07808f
C2951 _0663_/a_27_413# _0290_ 0.09411f
C2952 clknet_1_0__leaf__0465_ _0148_ 0.00276f
C2953 acc0.A\[14\] _0506_/a_81_21# 0
C2954 _1051_/a_466_413# _0525_/a_299_297# 0
C2955 _0216_ _0747_/a_215_47# 0.00638f
C2956 _0550_/a_240_47# net30 0.05957f
C2957 _0550_/a_245_297# _0137_ 0.00276f
C2958 _0550_/a_149_47# _0172_ 0.00103f
C2959 _0126_ _1008_/a_1059_315# 0
C2960 _0104_ _1006_/a_561_413# 0
C2961 _0432_ _0824_/a_145_75# 0.00139f
C2962 _0533_/a_27_297# acc0.A\[1\] 0.05719f
C2963 _0951_/a_209_311# _1062_/a_27_47# 0
C2964 _0951_/a_109_93# _1062_/a_193_47# 0
C2965 _0354_ _0353_ 0.16578f
C2966 _0349_ _0730_/a_510_47# 0
C2967 _0183_ _1060_/a_27_47# 0.06273f
C2968 _0174_ comp0.B\[12\] 0
C2969 net178 _0253_ 0
C2970 _0723_/a_207_413# _0334_ 0.22001f
C2971 hold24/a_285_47# _0206_ 0
C2972 net140 acc0.A\[6\] 0.10687f
C2973 B[12] _0542_/a_245_297# 0
C2974 hold64/a_285_47# _0241_ 0
C2975 _1000_/a_975_413# _0461_ 0
C2976 hold53/a_49_47# _1024_/a_193_47# 0
C2977 hold53/a_285_47# _1024_/a_27_47# 0
C2978 _0218_ net6 0.0214f
C2979 _0186_ net148 0.16709f
C2980 _0280_ _0369_ 0
C2981 _0262_ clknet_1_1__leaf__0457_ 0.00251f
C2982 VPWR _0474_ 0.66333f
C2983 net14 net12 0.04159f
C2984 _0275_ clknet_1_1__leaf__0458_ 0.06922f
C2985 _0272_ net72 0.00197f
C2986 hold33/a_285_47# comp0.B\[10\] 0
C2987 hold45/a_391_47# acc0.A\[11\] 0.04835f
C2988 input21/a_75_212# _0176_ 0
C2989 net55 _0707_/a_201_297# 0
C2990 _0216_ hold9/a_391_47# 0
C2991 _0240_ _0246_ 0.4539f
C2992 VPWR _1023_/a_891_413# 0.18788f
C2993 _1047_/a_466_413# clkbuf_1_1__f__0457_/a_110_47# 0.01042f
C2994 hold100/a_285_47# _0846_/a_240_47# 0
C2995 _1036_/a_1017_47# _0175_ 0
C2996 hold59/a_391_47# VPWR 0.18001f
C2997 hold38/a_285_47# net23 0
C2998 _0446_ _0844_/a_297_47# 0.0481f
C2999 _0369_ _0246_ 0
C3000 _0313_ _0106_ 0
C3001 clknet_1_1__leaf__0462_ hold50/a_49_47# 0.01445f
C3002 net45 _0129_ 0.00123f
C3003 _0991_/a_1059_315# _0991_/a_891_413# 0.31086f
C3004 _0991_/a_193_47# _0991_/a_975_413# 0
C3005 _0991_/a_466_413# _0991_/a_381_47# 0.03733f
C3006 _0726_/a_245_297# _0219_ 0.00125f
C3007 output36/a_27_47# VPWR 0.2556f
C3008 _0627_/a_215_53# _0186_ 0
C3009 _0837_/a_585_47# clknet_1_1__leaf__0458_ 0
C3010 acc0.A\[12\] _0402_ 0.11082f
C3011 _0218_ _0447_ 0
C3012 net21 net195 0.02287f
C3013 net23 clknet_1_1__leaf__0457_ 0
C3014 _0443_ _0269_ 0
C3015 _1014_/a_27_47# net206 0
C3016 output66/a_27_47# _0510_/a_109_297# 0
C3017 _0461_ _0565_/a_512_297# 0
C3018 _0216_ _1029_/a_634_159# 0.00779f
C3019 hold26/a_391_47# net157 0
C3020 net160 _0472_ 0.00402f
C3021 _0793_/a_149_47# _0345_ 0.00156f
C3022 _0080_ _1014_/a_27_47# 0
C3023 net68 _1014_/a_193_47# 0
C3024 _0982_/a_193_47# net100 0
C3025 _1004_/a_27_47# acc0.A\[23\] 0
C3026 net235 _0369_ 0.11147f
C3027 _0736_/a_311_297# _0462_ 0
C3028 _0316_ _0321_ 0.06979f
C3029 clknet_0__0459_ _0345_ 0.00226f
C3030 net7 _1046_/a_634_159# 0
C3031 _1001_/a_891_413# _0183_ 0
C3032 net123 _1037_/a_193_47# 0.00759f
C3033 clknet_1_0__leaf__0462_ _0195_ 0
C3034 _0250_ hold94/a_285_47# 0
C3035 _0249_ hold94/a_391_47# 0
C3036 _0399_ _0996_/a_381_47# 0.00376f
C3037 net186 _0132_ 0
C3038 acc0.A\[3\] _0345_ 0
C3039 net189 VPWR 0.33839f
C3040 _0984_/a_193_47# _0268_ 0
C3041 _0530_/a_81_21# _0465_ 0.00229f
C3042 _0800_/a_51_297# _0277_ 0
C3043 _0230_ _0762_/a_215_47# 0
C3044 _0598_/a_297_47# _0383_ 0.01213f
C3045 _0808_/a_266_47# _0418_ 0.04052f
C3046 acc0.A\[20\] _0181_ 0.00149f
C3047 _1021_/a_634_159# _0183_ 0
C3048 _1021_/a_891_413# net150 0.0093f
C3049 _1021_/a_1059_315# _0217_ 0.0064f
C3050 _1041_/a_381_47# clknet_1_0__leaf__0463_ 0.01223f
C3051 _0347_ _0321_ 0
C3052 _1002_/a_1059_315# _0760_/a_47_47# 0
C3053 _1060_/a_27_47# acc0.A\[15\] 0.01137f
C3054 net62 _0841_/a_79_21# 0
C3055 clkbuf_1_1__f__0461_/a_110_47# _0394_ 0
C3056 net31 hold5/a_391_47# 0
C3057 _0450_ _0841_/a_79_21# 0
C3058 _0348_ _0220_ 0.03103f
C3059 clknet_0__0457_ _0858_/a_27_47# 0
C3060 clkbuf_1_1__f__0463_/a_110_47# clknet_1_0__leaf__0461_ 0
C3061 _1058_/a_381_47# acc0.A\[10\] 0
C3062 acc0.A\[2\] _0530_/a_81_21# 0.05822f
C3063 _0391_ _0771_/a_382_47# 0
C3064 _0099_ _0771_/a_215_297# 0
C3065 _0366_ net93 0.03488f
C3066 acc0.A\[10\] _0420_ 0
C3067 comp0.B\[10\] net20 0
C3068 clknet_1_0__leaf__0465_ _0525_/a_384_47# 0
C3069 _0239_ _0775_/a_79_21# 0
C3070 _0522_/a_109_47# _0193_ 0.00325f
C3071 _0661_/a_27_297# _0346_ 0.09841f
C3072 _0351_ _0347_ 0
C3073 _0976_/a_76_199# _0488_ 0.06155f
C3074 hold87/a_285_47# acc0.A\[1\] 0
C3075 _0244_ _0387_ 0
C3076 net103 _0240_ 0
C3077 _0800_/a_149_47# _0412_ 0.01815f
C3078 pp[8] _0179_ 0.00245f
C3079 _0800_/a_512_297# _0413_ 0.0018f
C3080 acc0.A\[29\] net208 0
C3081 pp[27] _0723_/a_27_413# 0
C3082 _0461_ _1018_/a_891_413# 0
C3083 _0463_ _0176_ 0.02076f
C3084 net103 _0369_ 0.19772f
C3085 _0224_ net177 0
C3086 _0655_/a_109_93# _0345_ 0.01031f
C3087 _1011_/a_27_47# _1011_/a_193_47# 0.96574f
C3088 net201 _0563_/a_512_297# 0
C3089 _0170_ _1068_/a_634_159# 0
C3090 _0500_/a_27_47# net133 0.01774f
C3091 VPWR _0830_/a_297_297# 0.00835f
C3092 _0402_ _0650_/a_68_297# 0
C3093 hold86/a_285_47# _0260_ 0
C3094 VPWR _0312_ 0.76752f
C3095 _0343_ _0461_ 0.02881f
C3096 _1004_/a_381_47# net52 0.00398f
C3097 clkbuf_1_0__f__0461_/a_110_47# clknet_0__0461_ 0.31131f
C3098 VPWR _1031_/a_561_413# 0.00311f
C3099 _0504_/a_27_47# hold2/a_285_47# 0.02308f
C3100 _0350_ _1006_/a_27_47# 0.04599f
C3101 clknet_0__0465_ _0986_/a_634_159# 0.00427f
C3102 _0195_ _1019_/a_891_413# 0
C3103 _0268_ clkbuf_0__0458_/a_110_47# 0.11882f
C3104 _0714_/a_51_297# _0195_ 0.0176f
C3105 net46 _0219_ 0.04073f
C3106 net178 net74 0.13106f
C3107 acc0.A\[12\] _0648_/a_205_297# 0
C3108 _0217_ _0115_ 0
C3109 _0458_ _0449_ 0.00744f
C3110 _0425_ _0991_/a_891_413# 0
C3111 clkbuf_0_clk/a_110_47# _0971_/a_81_21# 0
C3112 _0572_/a_109_297# _1025_/a_27_47# 0
C3113 _1043_/a_1059_315# hold51/a_49_47# 0.0037f
C3114 _1043_/a_634_159# hold51/a_391_47# 0
C3115 net69 _0399_ 0.03166f
C3116 clknet_1_0__leaf__0462_ hold96/a_49_47# 0.01699f
C3117 _0372_ _0460_ 0.01586f
C3118 _0350_ _0986_/a_27_47# 0.00424f
C3119 _1020_/a_193_47# VPWR 0.31148f
C3120 _0851_/a_113_47# _0345_ 0
C3121 _0345_ _0418_ 0.01789f
C3122 _0820_/a_215_47# VPWR 0.00199f
C3123 clknet_0__0458_ _0446_ 0.0276f
C3124 _0835_/a_292_297# _0255_ 0
C3125 output66/a_27_47# _0188_ 0
C3126 _0955_/a_32_297# comp0.B\[3\] 0.16805f
C3127 acc0.A\[31\] _0220_ 0.01096f
C3128 _0159_ _0177_ 0
C3129 net172 net30 0
C3130 _0789_/a_75_199# _0297_ 0.22244f
C3131 _0150_ _0522_/a_109_297# 0.00149f
C3132 _0251_ hold65/a_391_47# 0
C3133 _0429_ hold65/a_49_47# 0
C3134 net49 _1022_/a_27_47# 0.00151f
C3135 _0837_/a_81_21# _0186_ 0
C3136 _0195_ net206 0.07078f
C3137 _0216_ net219 0
C3138 _1025_/a_381_47# acc0.A\[25\] 0.01613f
C3139 _0292_ _0819_/a_299_297# 0
C3140 net55 _1010_/a_27_47# 0.00848f
C3141 _1020_/a_193_47# _1015_/a_466_413# 0
C3142 _1020_/a_466_413# _1015_/a_193_47# 0
C3143 _0971_/a_299_297# _0460_ 0.00272f
C3144 _0181_ _0880_/a_27_47# 0.03527f
C3145 A[14] _0799_/a_80_21# 0
C3146 control0.reset _0565_/a_149_47# 0
C3147 hold101/a_49_47# clknet_1_0__leaf__0465_ 0
C3148 net240 _1067_/a_1059_315# 0
C3149 _0165_ _1067_/a_193_47# 0.39319f
C3150 net54 _0686_/a_219_297# 0
C3151 _0179_ _1060_/a_27_47# 0
C3152 clknet_1_0__leaf__0458_ _0991_/a_27_47# 0.01075f
C3153 _0080_ _0195_ 0
C3154 clknet_1_0__leaf__0457_ hold40/a_391_47# 0.00206f
C3155 control0.state\[2\] _0974_/a_222_93# 0.02558f
C3156 net54 _1008_/a_1059_315# 0.17834f
C3157 _0486_ _0974_/a_79_199# 0.08763f
C3158 clknet_1_1__leaf__0463_ _0496_/a_27_47# 0.00132f
C3159 control0.state\[1\] net23 0
C3160 _0183_ _0586_/a_27_47# 0
C3161 _0179_ _0988_/a_891_413# 0
C3162 _1019_/a_1059_315# _0369_ 0
C3163 hold20/a_285_47# _1072_/a_891_413# 0.00163f
C3164 hold20/a_391_47# _1072_/a_1059_315# 0.00124f
C3165 _0225_ net52 0
C3166 hold10/a_391_47# net201 0
C3167 clknet_0__0457_ _1019_/a_1059_315# 0
C3168 _0559_/a_240_47# comp0.B\[5\] 0
C3169 hold91/a_285_47# net41 0.08665f
C3170 _0972_/a_93_21# _0161_ 0
C3171 _0080_ _0856_/a_510_47# 0
C3172 _0531_/a_27_297# _1061_/a_27_47# 0
C3173 pp[27] _0352_ 0
C3174 _0800_/a_51_297# _0298_ 0
C3175 _0412_ _0789_/a_75_199# 0
C3176 _1021_/a_891_413# control0.add 0
C3177 net55 _1009_/a_193_47# 0.00241f
C3178 _1045_/a_193_47# clknet_1_1__leaf__0464_ 0
C3179 VPWR _0417_ 0.19994f
C3180 _1036_/a_634_159# _1036_/a_466_413# 0.23992f
C3181 _1036_/a_193_47# _1036_/a_1059_315# 0.03405f
C3182 _1036_/a_27_47# _1036_/a_891_413# 0.03224f
C3183 _1056_/a_634_159# _1056_/a_592_47# 0
C3184 _0422_ net37 0.00196f
C3185 _0346_ _0990_/a_27_47# 0.00128f
C3186 _0857_/a_27_47# _0181_ 0
C3187 _1047_/a_381_47# acc0.A\[15\] 0
C3188 _1030_/a_1059_315# hold61/a_285_47# 0.0129f
C3189 _0769_/a_384_47# _0386_ 0.00921f
C3190 _0769_/a_299_297# _0388_ 0.05973f
C3191 _0472_ acc0.A\[15\] 0.0014f
C3192 clknet_1_1__leaf_clk hold84/a_391_47# 0.00138f
C3193 _0984_/a_27_47# _1059_/a_27_47# 0
C3194 _1012_/a_27_47# _0778_/a_68_297# 0.00128f
C3195 hold90/a_285_47# _0319_ 0
C3196 _0183_ hold19/a_391_47# 0
C3197 _0993_/a_891_413# _0218_ 0
C3198 _0578_/a_27_297# _0578_/a_109_297# 0.17136f
C3199 _0644_/a_47_47# _0644_/a_285_47# 0.01755f
C3200 _1049_/a_27_47# net11 0
C3201 comp0.B\[5\] net29 0
C3202 comp0.B\[6\] B[6] 0
C3203 _0466_ clknet_0_clk 0.29731f
C3204 _0725_/a_80_21# _0725_/a_209_297# 0.06257f
C3205 _0158_ _0184_ 0.00579f
C3206 net43 _0459_ 0.00429f
C3207 net226 _0978_/a_373_47# 0.00131f
C3208 _0111_ _0340_ 0
C3209 clknet_1_0__leaf__0463_ _0553_/a_51_297# 0.00121f
C3210 _0090_ net67 0.02682f
C3211 _1041_/a_1059_315# _0544_/a_149_47# 0
C3212 output67/a_27_47# _0181_ 0
C3213 _0845_/a_193_297# _0350_ 0
C3214 clknet_1_0__leaf__0458_ _0350_ 0.72677f
C3215 clknet_1_0__leaf__0464_ clknet_1_1__leaf__0457_ 0
C3216 control0.state\[1\] net35 0.00251f
C3217 _0675_/a_68_297# net221 0
C3218 _0227_ _0577_/a_27_297# 0
C3219 _0437_ _0435_ 0.36216f
C3220 clknet_0__0457_ net68 0.02688f
C3221 clknet_1_0__leaf__0463_ _0953_/a_304_297# 0
C3222 net44 _0306_ 0.22268f
C3223 _1065_/a_193_47# _0215_ 0.00189f
C3224 _0403_ _0787_/a_303_47# 0
C3225 _0654_/a_27_413# _0417_ 0.00168f
C3226 _1065_/a_466_413# _0175_ 0
C3227 comp0.B\[13\] comp0.B\[12\] 0.24933f
C3228 hold11/a_285_47# _0144_ 0.08052f
C3229 net158 _0200_ 0
C3230 _0606_/a_465_297# _0383_ 0
C3231 _1041_/a_193_47# hold6/a_285_47# 0
C3232 _1041_/a_27_47# hold6/a_391_47# 0
C3233 _0852_/a_35_297# net206 0
C3234 net188 _1058_/a_466_413# 0
C3235 _0996_/a_27_47# _0219_ 0
C3236 _0343_ _0997_/a_1059_315# 0
C3237 clknet_1_0__leaf__0462_ net90 0.00458f
C3238 _0181_ _1062_/a_27_47# 0
C3239 _0314_ _0313_ 0.48709f
C3240 _0995_/a_634_159# _0297_ 0
C3241 input20/a_75_212# B[11] 0.01581f
C3242 _0804_/a_510_47# net39 0
C3243 _0804_/a_215_47# acc0.A\[12\] 0
C3244 _0402_ net42 0
C3245 net3 net67 0.08459f
C3246 _1052_/a_27_47# _0518_/a_27_297# 0
C3247 _0346_ _0671_/a_113_297# 0
C3248 clknet_0__0460_ _0320_ 0
C3249 clknet_1_1__leaf_clk _1065_/a_975_413# 0
C3250 _0777_/a_47_47# _0777_/a_285_47# 0.01755f
C3251 _1049_/a_466_413# _0465_ 0
C3252 net36 _1038_/a_381_47# 0.01572f
C3253 pp[0] _1038_/a_1059_315# 0
C3254 net61 _0825_/a_150_297# 0
C3255 hold47/a_285_47# _0142_ 0.09458f
C3256 _0985_/a_891_413# net58 0
C3257 _0428_ _0990_/a_193_47# 0.02654f
C3258 net61 _0844_/a_297_47# 0.0063f
C3259 _0467_ _0974_/a_544_297# 0
C3260 _0414_ _0399_ 0
C3261 _0760_/a_47_47# net91 0
C3262 _0722_/a_297_297# _0350_ 0
C3263 _0670_/a_215_47# net41 0.00837f
C3264 _0216_ _1028_/a_561_413# 0
C3265 _0467_ clknet_1_0__leaf__0457_ 0.0598f
C3266 _0736_/a_56_297# _0363_ 0.12949f
C3267 _1057_/a_466_413# _1057_/a_592_47# 0.00553f
C3268 _1057_/a_634_159# _1057_/a_1017_47# 0
C3269 _0553_/a_149_47# clknet_0__0463_ 0
C3270 B[13] _1042_/a_891_413# 0
C3271 clknet_1_1__leaf__0459_ _0301_ 0.0349f
C3272 _0269_ _0986_/a_891_413# 0
C3273 net211 net87 0.21041f
C3274 _0111_ _1013_/a_381_47# 0.13423f
C3275 VPWR _1064_/a_975_413# 0.00453f
C3276 _0081_ net206 0.00483f
C3277 _0454_ _0116_ 0
C3278 _0607_/a_27_297# clknet_0__0461_ 0.03375f
C3279 net236 clknet_0_clk 0
C3280 _0369_ net143 0.00136f
C3281 _1001_/a_1059_315# _1000_/a_27_47# 0
C3282 _1001_/a_27_47# _1000_/a_1059_315# 0
C3283 _1059_/a_634_159# _1059_/a_1017_47# 0
C3284 _1059_/a_466_413# _1059_/a_592_47# 0.00553f
C3285 VPWR _0669_/a_183_297# 0
C3286 hold78/a_49_47# VPWR 0.29316f
C3287 VPWR _0728_/a_145_75# 0
C3288 hold13/a_391_47# _0210_ 0.02068f
C3289 hold19/a_391_47# acc0.A\[15\] 0
C3290 hold76/a_285_47# net45 0
C3291 hold41/a_285_47# _0186_ 0.0054f
C3292 net36 _0452_ 0.07602f
C3293 _0528_/a_81_21# _0196_ 0.17319f
C3294 net222 _0082_ 0.00118f
C3295 _0568_/a_373_47# _0345_ 0.00108f
C3296 hold23/a_285_47# _0195_ 0.00497f
C3297 acc0.A\[7\] _0834_/a_109_297# 0
C3298 _0399_ net102 0
C3299 _0981_/a_109_297# VPWR 0.19326f
C3300 _0433_ _0989_/a_193_47# 0
C3301 _0433_ hold1/a_285_47# 0
C3302 _0181_ _1047_/a_634_159# 0
C3303 _0630_/a_109_297# _0219_ 0
C3304 comp0.B\[0\] clknet_1_0__leaf__0457_ 0
C3305 _0673_/a_103_199# _0673_/a_253_47# 0.06061f
C3306 _0515_/a_81_21# clknet_1_1__leaf__0465_ 0
C3307 acc0.A\[14\] _0184_ 0.01563f
C3308 _1002_/a_27_47# _0578_/a_27_297# 0
C3309 _0478_ _0489_ 0
C3310 _0388_ _0392_ 0.58356f
C3311 _0672_/a_79_21# _0672_/a_510_47# 0.00844f
C3312 _0672_/a_297_297# _0672_/a_215_47# 0
C3313 acc0.A\[0\] _0112_ 0
C3314 _0363_ net224 0.0993f
C3315 output43/a_27_47# hold98/a_391_47# 0
C3316 clknet_1_1__leaf__0459_ _0994_/a_193_47# 0
C3317 _1030_/a_466_413# clknet_1_1__leaf__0462_ 0
C3318 pp[17] net163 0
C3319 hold65/a_49_47# clknet_1_1__leaf__0458_ 0.00472f
C3320 _0984_/a_1059_315# _0350_ 0.02025f
C3321 _0349_ _0336_ 0
C3322 _0302_ net228 0.04487f
C3323 net158 net193 0
C3324 net233 _0846_/a_240_47# 0.08819f
C3325 _0715_/a_27_47# _0990_/a_193_47# 0
C3326 _0324_ _1026_/a_27_47# 0
C3327 acc0.A\[27\] net114 0.22873f
C3328 _0343_ net179 0
C3329 _1054_/a_193_47# _0087_ 0
C3330 VPWR _1008_/a_466_413# 0.26038f
C3331 _0129_ VPWR 0.36757f
C3332 net158 _1046_/a_466_413# 0.00203f
C3333 _0467_ _1062_/a_466_413# 0
C3334 _0464_ _0172_ 0
C3335 _0201_ net18 0
C3336 _0362_ _0685_/a_68_297# 0
C3337 _0216_ _0352_ 0.75306f
C3338 acc0.A\[13\] _0668_/a_79_21# 0
C3339 _0126_ clknet_1_1__leaf__0462_ 0.05893f
C3340 _0785_/a_299_297# _0819_/a_299_297# 0.06921f
C3341 net101 _0713_/a_27_47# 0.00297f
C3342 _0624_/a_59_75# _0624_/a_145_75# 0.00658f
C3343 clkload1/Y VPWR 0.43946f
C3344 _0368_ clkbuf_1_0__f__0462_/a_110_47# 0.00754f
C3345 _0183_ net149 0.05611f
C3346 hold38/a_49_47# _0173_ 0
C3347 hold38/a_285_47# _0213_ 0.00193f
C3348 _0399_ _0300_ 0.05159f
C3349 _0149_ _0525_/a_299_297# 0.00103f
C3350 _0637_/a_56_297# net247 0
C3351 _0467_ _0561_/a_149_47# 0
C3352 clknet_0__0462_ _0319_ 0.0091f
C3353 acc0.A\[1\] _0199_ 0.00161f
C3354 _0180_ net8 0.24635f
C3355 net34 clkbuf_0_clk/a_110_47# 0
C3356 comp0.B\[0\] _1062_/a_466_413# 0
C3357 net200 _1026_/a_193_47# 0
C3358 _0982_/a_27_47# clkbuf_1_1__f__0457_/a_110_47# 0
C3359 clknet_0__0458_ net61 0.00225f
C3360 hold28/a_49_47# clknet_1_1__leaf__0457_ 0
C3361 pp[18] hold78/a_285_47# 0.00151f
C3362 _0181_ net107 0
C3363 acc0.A\[24\] net93 0.03388f
C3364 _0469_ _0950_/a_75_212# 0.29289f
C3365 input31/a_75_212# _0546_/a_240_47# 0
C3366 net31 _0546_/a_51_297# 0
C3367 VPWR _0563_/a_51_297# 0.47208f
C3368 _0457_ _1034_/a_27_47# 0
C3369 net16 A[9] 0.04465f
C3370 control0.state\[1\] _1063_/a_466_413# 0.03261f
C3371 net105 _1014_/a_466_413# 0.00147f
C3372 clknet_1_0__leaf__0462_ _1022_/a_561_413# 0
C3373 _1005_/a_193_47# _1005_/a_891_413# 0.19489f
C3374 _1005_/a_27_47# _1005_/a_381_47# 0.06222f
C3375 _1005_/a_634_159# _1005_/a_1059_315# 0
C3376 _1067_/a_27_47# _0352_ 0
C3377 net55 _0339_ 0
C3378 VPWR _0511_/a_384_47# 0
C3379 _0519_/a_81_21# _0519_/a_384_47# 0.00138f
C3380 _0559_/a_51_297# comp0.B\[4\] 0
C3381 net152 net32 0.54097f
C3382 _0145_ clkbuf_1_1__f__0457_/a_110_47# 0.01075f
C3383 _0984_/a_193_47# net222 0
C3384 _0195_ _0405_ 0
C3385 _1013_/a_27_47# _1013_/a_466_413# 0.27314f
C3386 _1013_/a_193_47# _1013_/a_634_159# 0.11897f
C3387 comp0.B\[14\] _0142_ 0.02782f
C3388 acc0.A\[27\] _0365_ 0.31209f
C3389 _0991_/a_381_47# _0089_ 0.13435f
C3390 _0991_/a_466_413# net67 0
C3391 VPWR _0541_/a_68_297# 0.16193f
C3392 net185 clknet_0__0463_ 0
C3393 VPWR _0746_/a_299_297# 0.28199f
C3394 _0195_ _0356_ 0.00551f
C3395 net185 hold38/a_391_47# 0.13554f
C3396 _0212_ hold38/a_285_47# 0
C3397 _0891_/a_27_47# _0566_/a_27_47# 0
C3398 _0309_ _0775_/a_79_21# 0
C3399 hold96/a_391_47# _0352_ 0
C3400 hold96/a_285_47# _0102_ 0
C3401 _1000_/a_891_413# clknet_1_0__leaf__0461_ 0.00141f
C3402 _0462_ _0743_/a_149_47# 0
C3403 _0607_/a_27_297# _0607_/a_373_47# 0.01338f
C3404 _0985_/a_1059_315# _0261_ 0.02254f
C3405 _0985_/a_891_413# _0262_ 0
C3406 clknet_1_1__leaf__0459_ _0997_/a_634_159# 0.01443f
C3407 _0216_ net115 0.05156f
C3408 _0646_/a_47_47# _0995_/a_466_413# 0
C3409 _0574_/a_109_297# _0216_ 0.05362f
C3410 clknet_1_1__leaf__0459_ _0992_/a_381_47# 0.01109f
C3411 _0214_ _0171_ 0.00441f
C3412 _0291_ acc0.A\[9\] 0.16573f
C3413 _0559_/a_149_47# net26 0.00362f
C3414 _0274_ _0642_/a_215_297# 0.11896f
C3415 hold31/a_391_47# _0086_ 0.00386f
C3416 _1038_/a_634_159# _1040_/a_193_47# 0
C3417 _1038_/a_466_413# _1040_/a_27_47# 0
C3418 _1038_/a_193_47# _1040_/a_634_159# 0
C3419 VPWR _1065_/a_592_47# 0
C3420 _0260_ _0458_ 0.14902f
C3421 net228 net6 0
C3422 _0600_/a_253_297# _0223_ 0.00626f
C3423 _1012_/a_193_47# hold92/a_391_47# 0
C3424 net149 acc0.A\[15\] 0.06983f
C3425 _0217_ net223 0
C3426 _0764_/a_81_21# _0373_ 0.062f
C3427 _1018_/a_891_413# _0582_/a_27_297# 0
C3428 _1018_/a_1059_315# _0582_/a_109_297# 0
C3429 clknet_1_0__leaf__0463_ _0135_ 0.00334f
C3430 _0462_ _0345_ 0.04519f
C3431 _0766_/a_109_297# _0245_ 0.00107f
C3432 _1038_/a_975_413# comp0.B\[4\] 0
C3433 _0995_/a_1059_315# _0995_/a_891_413# 0.31086f
C3434 _0995_/a_193_47# _0995_/a_975_413# 0
C3435 _0995_/a_466_413# _0995_/a_381_47# 0.03733f
C3436 hold10/a_49_47# VPWR 0.28319f
C3437 hold76/a_49_47# net46 0.32453f
C3438 clknet_1_0__leaf__0457_ acc0.A\[19\] 0.12977f
C3439 _0365_ _0364_ 0.15708f
C3440 _0543_/a_68_297# _0142_ 0
C3441 _0343_ _0582_/a_27_297# 0.01958f
C3442 output56/a_27_47# _0350_ 0
C3443 _0983_/a_634_159# _0346_ 0
C3444 hold18/a_49_47# _0350_ 0.00136f
C3445 net59 hold95/a_285_47# 0
C3446 _1070_/a_193_47# _0489_ 0
C3447 VPWR _0549_/a_68_297# 0.16964f
C3448 _1034_/a_891_413# _0561_/a_51_297# 0
C3449 _1017_/a_27_47# _0675_/a_68_297# 0.00793f
C3450 net245 _0668_/a_79_21# 0.00133f
C3451 net40 _0668_/a_297_47# 0
C3452 output36/a_27_47# net30 0
C3453 net23 _1066_/a_634_159# 0
C3454 clknet_0_clk _1065_/a_634_159# 0.00827f
C3455 clknet_1_0__leaf__0465_ _1048_/a_27_47# 0
C3456 net152 _1042_/a_1059_315# 0
C3457 _0139_ _1042_/a_27_47# 0
C3458 net32 _1042_/a_466_413# 0.03302f
C3459 net165 _0635_/a_27_47# 0.04334f
C3460 _0123_ _0315_ 0
C3461 _1018_/a_193_47# _0459_ 0.00467f
C3462 hold85/a_285_47# control0.state\[2\] 0
C3463 hold57/a_391_47# net204 0.13065f
C3464 net53 _1007_/a_1017_47# 0
C3465 _1019_/a_27_47# _0580_/a_27_297# 0
C3466 VPWR _1069_/a_27_47# 0.56965f
C3467 _0293_ _0346_ 0.09087f
C3468 control0.state\[1\] _1062_/a_561_413# 0
C3469 control0.state\[0\] _1062_/a_975_413# 0.00256f
C3470 _0413_ _0093_ 0.00653f
C3471 _0982_/a_466_413# _0183_ 0.00608f
C3472 _0982_/a_891_413# _0217_ 0
C3473 pp[6] _0369_ 0
C3474 _0404_ _0399_ 0.51944f
C3475 _1034_/a_466_413# _0473_ 0
C3476 pp[28] hold95/a_391_47# 0
C3477 hold25/a_391_47# A[1] 0.00131f
C3478 acc0.A\[30\] hold62/a_391_47# 0
C3479 _0180_ net10 0.65254f
C3480 _1011_/a_466_413# _1011_/a_592_47# 0.00553f
C3481 _1011_/a_634_159# _1011_/a_1017_47# 0
C3482 _0133_ _1034_/a_891_413# 0.00222f
C3483 _0171_ _1061_/a_1059_315# 0
C3484 _1006_/a_27_47# _1006_/a_634_159# 0.14145f
C3485 pp[1] net62 0.12033f
C3486 comp0.B\[1\] _1067_/a_466_413# 0
C3487 net152 net10 0.03976f
C3488 _0247_ _0773_/a_285_297# 0
C3489 _0216_ net207 0.01945f
C3490 _0287_ _0992_/a_1059_315# 0
C3491 _0972_/a_250_297# _0487_ 0.02147f
C3492 net225 _0195_ 0.03071f
C3493 _0275_ _0218_ 0.00574f
C3494 _0964_/a_109_297# _0480_ 0.0019f
C3495 _0751_/a_29_53# _0751_/a_183_297# 0.00868f
C3496 net55 hold97/a_49_47# 0
C3497 _0401_ net67 0.04778f
C3498 _0124_ _1025_/a_193_47# 0
C3499 _1055_/a_891_413# VPWR 0.21738f
C3500 net196 hold51/a_285_47# 0
C3501 _1018_/a_634_159# clknet_1_0__leaf__0461_ 0.00398f
C3502 _0238_ _0771_/a_215_297# 0
C3503 _1001_/a_1059_315# acc0.A\[19\] 0
C3504 _0102_ _1024_/a_27_47# 0
C3505 _1003_/a_1059_315# VPWR 0.4068f
C3506 _0429_ _0828_/a_199_47# 0.00917f
C3507 clknet_0__0464_ _1049_/a_466_413# 0
C3508 _0837_/a_585_47# _0218_ 0
C3509 net54 clknet_1_1__leaf__0462_ 0.0589f
C3510 _0183_ _0094_ 0.00359f
C3511 comp0.B\[5\] comp0.B\[6\] 0.15906f
C3512 clkbuf_1_0__f__0463_/a_110_47# _0176_ 0.00309f
C3513 comp0.B\[3\] _0474_ 0.01881f
C3514 output67/a_27_47# _0187_ 0
C3515 hold74/a_49_47# _0218_ 0
C3516 _0959_/a_217_297# _0163_ 0
C3517 _0986_/a_27_47# _0986_/a_634_159# 0.14145f
C3518 _0299_ _0300_ 0.05755f
C3519 _0298_ _0277_ 0.17022f
C3520 _0089_ _0082_ 0
C3521 _0585_/a_109_47# _0181_ 0
C3522 net148 _0987_/a_634_159# 0
C3523 _0297_ _0345_ 0
C3524 _0311_ _0218_ 0
C3525 _0225_ hold94/a_391_47# 0.01753f
C3526 clkload4/Y _0114_ 0.00782f
C3527 net126 A[15] 0
C3528 _0252_ _0435_ 0
C3529 _0443_ clkbuf_0__0458_/a_110_47# 0.00946f
C3530 _1020_/a_193_47# _0113_ 0
C3531 _0118_ _1015_/a_193_47# 0
C3532 _0732_/a_80_21# hold90/a_285_47# 0
C3533 _1023_/a_27_47# _1023_/a_891_413# 0.03224f
C3534 _1023_/a_193_47# _1023_/a_1059_315# 0.03405f
C3535 _1023_/a_634_159# _1023_/a_466_413# 0.23992f
C3536 clkbuf_1_0__f__0461_/a_110_47# _0616_/a_215_47# 0
C3537 _0247_ _0350_ 0
C3538 _0170_ _0479_ 0
C3539 clkload2/Y _0180_ 0.00183f
C3540 clknet_1_0__leaf__0463_ _0497_/a_150_297# 0
C3541 _1042_/a_193_47# _1042_/a_381_47# 0.09503f
C3542 _1042_/a_634_159# _1042_/a_891_413# 0.03684f
C3543 _1042_/a_27_47# _1042_/a_561_413# 0.00163f
C3544 hold100/a_391_47# acc0.A\[15\] 0.01316f
C3545 _0296_ _0277_ 0
C3546 _0181_ _1060_/a_561_413# 0
C3547 control0.add _0391_ 0
C3548 _0516_/a_27_297# net16 0.18142f
C3549 _1010_/a_561_413# _0352_ 0
C3550 _0290_ acc0.A\[9\] 0.76683f
C3551 _0982_/a_466_413# acc0.A\[15\] 0
C3552 _0734_/a_129_47# _0317_ 0
C3553 clknet_1_1__leaf__0464_ _1044_/a_27_47# 0.05576f
C3554 _1011_/a_27_47# _0707_/a_75_199# 0
C3555 _0174_ _0181_ 0
C3556 _1045_/a_27_47# _0202_ 0
C3557 VPWR hold61/a_285_47# 0.28607f
C3558 _1017_/a_193_47# _0307_ 0
C3559 clknet_1_1__leaf__0460_ _0357_ 0.0628f
C3560 net231 _0161_ 0.21069f
C3561 _0412_ _0345_ 0.068f
C3562 _0800_/a_240_47# _0219_ 0.02833f
C3563 _0850_/a_68_297# net165 0
C3564 _0216_ _0551_/a_27_47# 0
C3565 _1021_/a_27_47# net118 0
C3566 _1036_/a_634_159# net161 0.00197f
C3567 _0997_/a_381_47# _0587_/a_27_47# 0
C3568 net10 _1042_/a_466_413# 0.00542f
C3569 _0229_ hold66/a_285_47# 0
C3570 _0153_ _0988_/a_634_159# 0
C3571 hold76/a_285_47# VPWR 0.28449f
C3572 _0248_ net223 0
C3573 net221 _0242_ 0
C3574 _1057_/a_27_47# _0511_/a_81_21# 0
C3575 VPWR _1040_/a_891_413# 0.18556f
C3576 _0992_/a_634_159# clknet_1_1__leaf__0465_ 0
C3577 hold52/a_391_47# hold68/a_285_47# 0
C3578 hold52/a_285_47# hold68/a_391_47# 0
C3579 control0.state\[2\] _0958_/a_27_47# 0.01261f
C3580 _0129_ _0567_/a_373_47# 0
C3581 hold27/a_285_47# _0159_ 0
C3582 net163 _0567_/a_109_297# 0
C3583 _0294_ _0583_/a_109_297# 0.00835f
C3584 _0218_ _0583_/a_27_297# 0
C3585 _1000_/a_193_47# _0241_ 0
C3586 _0997_/a_27_47# _0793_/a_240_47# 0
C3587 _0343_ _0254_ 0
C3588 _1050_/a_975_413# _0194_ 0
C3589 _0410_ _0406_ 0
C3590 _0094_ acc0.A\[15\] 0.00688f
C3591 hold31/a_49_47# clkbuf_1_1__f__0458_/a_110_47# 0
C3592 hold38/a_285_47# _0161_ 0
C3593 clknet_1_0__leaf__0462_ _1026_/a_381_47# 0
C3594 _1011_/a_1059_315# _0334_ 0
C3595 hold88/a_391_47# output47/a_27_47# 0
C3596 B[9] comp0.B\[10\] 0.00788f
C3597 _0455_ _0350_ 0
C3598 _0483_ _0490_ 0.19479f
C3599 hold49/a_391_47# _0141_ 0.05237f
C3600 clknet_1_0__leaf__0458_ _0986_/a_634_159# 0
C3601 _1002_/a_1059_315# _0765_/a_79_21# 0.01742f
C3602 _0271_ _0445_ 0
C3603 _0163_ _1062_/a_592_47# 0
C3604 clknet_1_0__leaf__0462_ _1024_/a_1017_47# 0
C3605 _0467_ _1063_/a_1017_47# 0
C3606 _0596_/a_59_75# _0237_ 0
C3607 _1058_/a_592_47# net4 0
C3608 _0368_ net51 0
C3609 _0511_/a_299_297# _0286_ 0
C3610 net61 _0627_/a_109_93# 0
C3611 _0428_ clknet_1_1__leaf__0465_ 0.00648f
C3612 _0399_ net16 0
C3613 _0195_ hold71/a_285_47# 0.00234f
C3614 _1032_/a_466_413# _1067_/a_634_159# 0
C3615 _1032_/a_634_159# _1067_/a_466_413# 0
C3616 _1032_/a_27_47# _1067_/a_891_413# 0
C3617 _1032_/a_891_413# _1067_/a_27_47# 0
C3618 _1052_/a_27_47# _0191_ 0
C3619 _0147_ _0465_ 0.00217f
C3620 _0615_/a_109_297# clknet_1_0__leaf__0461_ 0
C3621 _0660_/a_113_47# clknet_1_1__leaf__0465_ 0
C3622 clkload0/X clknet_0_clk 0.00174f
C3623 comp0.B\[11\] hold5/a_391_47# 0
C3624 hold68/a_391_47# net52 0
C3625 _0371_ _0366_ 0
C3626 _0999_/a_193_47# _0218_ 0.23703f
C3627 _0183_ _0393_ 0.08609f
C3628 _1054_/a_891_413# acc0.A\[7\] 0
C3629 _0258_ _0438_ 0
C3630 _0346_ _0655_/a_369_297# 0
C3631 _0618_/a_215_47# net51 0.00226f
C3632 net190 hold8/a_391_47# 0
C3633 _0777_/a_47_47# _0219_ 0
C3634 _0462_ net52 0.00738f
C3635 clknet_1_0__leaf__0464_ _1049_/a_634_159# 0.00198f
C3636 acc0.A\[2\] _0147_ 0.27393f
C3637 _1058_/a_193_47# acc0.A\[11\] 0.00238f
C3638 _0736_/a_139_47# _0219_ 0.01077f
C3639 _0457_ _0565_/a_149_47# 0
C3640 clknet_1_1__leaf__0459_ _0809_/a_384_47# 0
C3641 _0287_ _0421_ 0
C3642 hold64/a_285_47# _0352_ 0
C3643 VPWR _1035_/a_27_47# 0.67619f
C3644 _1053_/a_466_413# _1052_/a_466_413# 0
C3645 _1053_/a_193_47# _1052_/a_891_413# 0
C3646 _1053_/a_891_413# _1052_/a_193_47# 0
C3647 _0550_/a_149_47# _1040_/a_193_47# 0
C3648 _0550_/a_240_47# _1040_/a_27_47# 0
C3649 _0217_ _0758_/a_215_47# 0
C3650 _0358_ clkbuf_1_1__f__0462_/a_110_47# 0
C3651 hold22/a_49_47# _0437_ 0
C3652 _0404_ _0299_ 0.01136f
C3653 _0181_ _0208_ 0.12487f
C3654 _0224_ hold4/a_49_47# 0
C3655 _0643_/a_253_47# _0271_ 0
C3656 _0754_/a_245_297# _0345_ 0
C3657 control0.sh net171 0.00621f
C3658 _0230_ _0315_ 0
C3659 _0539_/a_150_297# VPWR 0.00165f
C3660 hold37/a_49_47# _0142_ 0
C3661 _1034_/a_27_47# net27 0
C3662 B[1] _0175_ 0
C3663 _0216_ net106 0
C3664 net4 _0186_ 0.0379f
C3665 _0314_ _0321_ 0
C3666 _0217_ _0487_ 0
C3667 _0313_ _0360_ 0.02285f
C3668 _0458_ _0643_/a_103_199# 0
C3669 _1055_/a_975_413# clknet_1_1__leaf__0465_ 0
C3670 _0314_ clkbuf_0__0460_/a_110_47# 0
C3671 net44 _0778_/a_68_297# 0.16398f
C3672 _0341_ _0342_ 0.16147f
C3673 net120 _0132_ 0
C3674 _0176_ _1042_/a_1017_47# 0
C3675 _0396_ _0347_ 0.00107f
C3676 _0508_/a_299_297# acc0.A\[15\] 0.00119f
C3677 clk _1068_/a_27_47# 0
C3678 clkbuf_0_clk/a_110_47# _1068_/a_466_413# 0.00204f
C3679 clknet_0__0457_ hold71/a_49_47# 0.00237f
C3680 _0555_/a_240_47# _0210_ 0
C3681 _0186_ hold83/a_391_47# 0.00213f
C3682 _1038_/a_634_159# _0207_ 0
C3683 _1026_/a_27_47# _1025_/a_27_47# 0.07618f
C3684 net24 control0.sh 0.02235f
C3685 _0959_/a_217_297# _1066_/a_27_47# 0
C3686 _0748_/a_81_21# _0250_ 0
C3687 B[12] net18 0
C3688 _0551_/a_27_47# net247 0
C3689 _0243_ hold76/a_391_47# 0.00371f
C3690 _0734_/a_285_47# clknet_1_1__leaf__0460_ 0
C3691 clknet_0__0458_ _0431_ 0.00367f
C3692 control0.state\[0\] net232 0.01252f
C3693 net247 _0849_/a_79_21# 0
C3694 _0329_ acc0.A\[29\] 0.00325f
C3695 VPWR _0994_/a_891_413# 0.18343f
C3696 _0343_ _1060_/a_634_159# 0
C3697 net159 _1068_/a_193_47# 0.00184f
C3698 net169 _0437_ 0
C3699 _0461_ clkbuf_0__0461_/a_110_47# 0.32323f
C3700 net167 clkbuf_1_0__f_clk/a_110_47# 0
C3701 output60/a_27_47# pp[14] 0
C3702 pp[31] output41/a_27_47# 0
C3703 net1 clknet_1_0__leaf__0457_ 0.0325f
C3704 _0486_ net17 0
C3705 _0230_ net150 0
C3706 _0229_ _0183_ 0
C3707 _0226_ _0217_ 0
C3708 net39 _0807_/a_68_297# 0
C3709 _0461_ _1015_/a_891_413# 0
C3710 net106 _1067_/a_27_47# 0
C3711 _1038_/a_466_413# net24 0
C3712 _0179_ A[10] 0.17026f
C3713 _1010_/a_466_413# _0350_ 0.0383f
C3714 pp[27] _1011_/a_466_413# 0
C3715 _0467_ _0160_ 0.3249f
C3716 hold75/a_391_47# _0219_ 0.05819f
C3717 _0557_/a_245_297# clknet_1_1__leaf__0463_ 0
C3718 _0646_/a_285_47# _0299_ 0
C3719 _0737_/a_35_297# _0737_/a_285_297# 0.02504f
C3720 net22 _0206_ 0
C3721 net86 net221 0
C3722 _0259_ _0990_/a_27_47# 0.00234f
C3723 net45 _0582_/a_109_47# 0
C3724 net89 _0166_ 0
C3725 _0216_ _0769_/a_299_297# 0
C3726 _0565_/a_51_297# _0173_ 0.116f
C3727 _0289_ _0809_/a_299_297# 0.00863f
C3728 _0287_ _0809_/a_81_21# 0.0613f
C3729 _0708_/a_68_297# _0220_ 0
C3730 _0341_ _1013_/a_592_47# 0
C3731 _0663_/a_207_413# _0369_ 0.00885f
C3732 net157 _1061_/a_466_413# 0.00433f
C3733 _0699_/a_68_297# _0329_ 0.01733f
C3734 _0961_/a_113_297# control0.count\[0\] 0.04938f
C3735 _0846_/a_245_297# _0350_ 0.00266f
C3736 hold70/a_285_47# hold70/a_391_47# 0.41909f
C3737 hold36/a_391_47# _0538_/a_51_297# 0.01217f
C3738 _0383_ _0381_ 0.02155f
C3739 _0221_ acc0.A\[29\] 0.14291f
C3740 _0995_/a_466_413# _0219_ 0
C3741 clkbuf_1_0__f__0462_/a_110_47# clknet_0__0460_ 0
C3742 _0174_ _0544_/a_240_47# 0.01381f
C3743 _0695_/a_217_297# _0312_ 0.01809f
C3744 _1009_/a_1059_315# _0350_ 0
C3745 net8 _0498_/a_51_297# 0
C3746 _0533_/a_27_297# net247 0
C3747 _0222_ _0223_ 0.15594f
C3748 _1034_/a_27_47# _1033_/a_193_47# 0
C3749 _1034_/a_193_47# _1033_/a_27_47# 0
C3750 _0217_ _1016_/a_193_47# 0
C3751 net108 _0217_ 0
C3752 clknet_1_0__leaf__0462_ _0183_ 0.10227f
C3753 clkbuf_1_0__f__0464_/a_110_47# clknet_1_1__leaf__0457_ 0
C3754 _0596_/a_59_75# _1005_/a_27_47# 0.00486f
C3755 _1031_/a_1059_315# _1031_/a_891_413# 0.31086f
C3756 _1031_/a_193_47# _1031_/a_975_413# 0
C3757 _1031_/a_466_413# _1031_/a_381_47# 0.03733f
C3758 _0531_/a_27_297# _1047_/a_634_159# 0
C3759 _0531_/a_109_297# _1047_/a_193_47# 0
C3760 comp0.B\[0\] _0160_ 0.00815f
C3761 _0240_ hold72/a_391_47# 0
C3762 clknet_1_0__leaf__0463_ _0206_ 0.06983f
C3763 net224 _0686_/a_219_297# 0
C3764 clknet_0__0462_ _0250_ 0
C3765 net67 hold70/a_49_47# 0.06285f
C3766 _0369_ hold72/a_391_47# 0.00404f
C3767 net82 _0343_ 0.00254f
C3768 hold30/a_285_47# _0756_/a_47_47# 0
C3769 _1041_/a_27_47# VPWR 0.41199f
C3770 comp0.B\[10\] hold6/a_285_47# 0
C3771 control0.state\[1\] _0161_ 0.15649f
C3772 _1000_/a_891_413# _0218_ 0
C3773 _1000_/a_381_47# _0294_ 0
C3774 _1005_/a_1059_315# net91 0
C3775 _1005_/a_466_413# _0103_ 0.03058f
C3776 _0179_ _0508_/a_299_297# 0.0826f
C3777 _0157_ _0656_/a_59_75# 0
C3778 _0465_ _0842_/a_59_75# 0.00208f
C3779 _0244_ _0247_ 0.58051f
C3780 _0481_ control0.state\[2\] 0.0016f
C3781 _0699_/a_68_297# _0221_ 0
C3782 comp0.B\[5\] net26 0.03779f
C3783 _0274_ net63 0
C3784 _0984_/a_592_47# _0082_ 0.00164f
C3785 _1060_/a_193_47# net5 0
C3786 net15 A[8] 0.02427f
C3787 _1013_/a_1059_315# _1013_/a_1017_47# 0
C3788 _0089_ net67 0
C3789 net1 _1062_/a_466_413# 0
C3790 _1002_/a_634_159# _1002_/a_975_413# 0
C3791 _1002_/a_466_413# _1002_/a_561_413# 0.00772f
C3792 _0770_/a_79_21# _0869_/a_27_47# 0
C3793 _1021_/a_193_47# net1 0.00235f
C3794 clknet_1_0__leaf__0465_ _0524_/a_373_47# 0
C3795 acc0.A\[21\] _0486_ 0.00462f
C3796 _0640_/a_297_297# VPWR 0
C3797 _0217_ clkbuf_0__0457_/a_110_47# 0.01528f
C3798 _0758_/a_297_297# _0379_ 0.00226f
C3799 _0319_ _0687_/a_59_75# 0.1308f
C3800 _0268_ _0447_ 0.0044f
C3801 _0984_/a_381_47# clknet_1_0__leaf__0458_ 0
C3802 net63 _0837_/a_266_47# 0
C3803 _0372_ _0373_ 0
C3804 _0087_ acc0.A\[6\] 0.02726f
C3805 net22 _1046_/a_1059_315# 0
C3806 _0965_/a_129_47# clknet_1_0__leaf_clk 0.00158f
C3807 hold28/a_391_47# _1049_/a_27_47# 0
C3808 hold28/a_285_47# _1049_/a_193_47# 0
C3809 acc0.A\[18\] _0611_/a_68_297# 0.02037f
C3810 _0552_/a_68_297# _0173_ 0
C3811 VPWR _0997_/a_381_47# 0.0874f
C3812 hold64/a_285_47# net207 0
C3813 net172 _1040_/a_27_47# 0
C3814 _1059_/a_1059_315# _0369_ 0.00396f
C3815 _0183_ _1019_/a_891_413# 0.00855f
C3816 _0217_ _1019_/a_561_413# 0
C3817 VPWR _0992_/a_1017_47# 0
C3818 _0316_ _0332_ 0
C3819 _1018_/a_891_413# _0115_ 0
C3820 net104 _0582_/a_373_47# 0
C3821 net248 acc0.A\[5\] 0.14212f
C3822 net227 clknet_1_1__leaf__0462_ 0
C3823 _0664_/a_79_21# clknet_1_1__leaf__0459_ 0.0029f
C3824 _0285_ _0653_/a_113_47# 0.00937f
C3825 _0765_/a_215_47# net220 0.0537f
C3826 _1035_/a_891_413# _0175_ 0
C3827 _0965_/a_47_47# _0974_/a_79_199# 0
C3828 _0230_ _0742_/a_81_21# 0
C3829 pp[28] _1011_/a_634_159# 0
C3830 net23 _0564_/a_68_297# 0
C3831 net55 _0685_/a_150_297# 0
C3832 _0316_ _0685_/a_68_297# 0
C3833 VPWR _1061_/a_975_413# 0.00494f
C3834 net77 acc0.A\[9\] 0
C3835 net67 _0656_/a_145_75# 0.00147f
C3836 _0343_ _0115_ 0.00594f
C3837 clknet_1_0__leaf__0463_ _1046_/a_1059_315# 0
C3838 _0332_ _0347_ 0.0023f
C3839 net69 _0346_ 0.20559f
C3840 clkbuf_1_0__f__0461_/a_110_47# _0771_/a_215_297# 0
C3841 output55/a_27_47# _0334_ 0.08271f
C3842 VPWR _0489_ 1.01441f
C3843 _0244_ _0455_ 0
C3844 VPWR _0668_/a_79_21# 0.23798f
C3845 net63 pp[5] 0.09731f
C3846 _1034_/a_592_47# _0213_ 0.00141f
C3847 _1034_/a_975_413# _0173_ 0
C3848 _1034_/a_891_413# _0208_ 0.00297f
C3849 _0971_/a_81_21# _0487_ 0.0619f
C3850 _0183_ net206 0.14316f
C3851 VPWR hold7/a_285_47# 0.29389f
C3852 _0176_ _0548_/a_245_297# 0
C3853 acc0.A\[4\] _0142_ 0
C3854 net23 clknet_1_1__leaf_clk 0.8206f
C3855 _0985_/a_27_47# _0446_ 0
C3856 _0343_ _0796_/a_297_297# 0
C3857 _0811_/a_81_21# _0296_ 0
C3858 hold31/a_285_47# acc0.A\[8\] 0.00956f
C3859 hold10/a_285_47# _0924_/a_27_47# 0.00508f
C3860 clknet_1_0__leaf__0458_ _1014_/a_27_47# 0
C3861 control0.count\[1\] _1069_/a_381_47# 0.00152f
C3862 _1070_/a_381_47# control0.count\[0\] 0
C3863 _0226_ _0248_ 0
C3864 _0080_ _0183_ 0.00338f
C3865 input1/a_27_47# input17/a_75_212# 0.01246f
C3866 B[13] B[10] 0.00508f
C3867 _1030_/a_193_47# _0336_ 0.00866f
C3868 net185 _1066_/a_466_413# 0
C3869 _0212_ _1066_/a_634_159# 0
C3870 _1056_/a_1059_315# _1058_/a_1059_315# 0.00209f
C3871 clkbuf_1_0__f__0458_/a_110_47# _0849_/a_215_47# 0
C3872 pp[17] net116 0
C3873 _0762_/a_215_47# _1005_/a_891_413# 0
C3874 _0369_ _1005_/a_193_47# 0
C3875 _1011_/a_381_47# net57 0
C3876 _0216_ _1011_/a_466_413# 0
C3877 _1000_/a_27_47# _0246_ 0
C3878 _0572_/a_27_297# _0572_/a_109_297# 0.17136f
C3879 _0601_/a_68_297# _0219_ 0.00546f
C3880 _0276_ hold91/a_49_47# 0
C3881 clkbuf_0__0462_/a_110_47# _0318_ 0.00182f
C3882 _1006_/a_381_47# _1006_/a_561_413# 0.00123f
C3883 _1006_/a_27_47# net92 0.22517f
C3884 _1006_/a_891_413# _1006_/a_975_413# 0.00851f
C3885 _0180_ _0146_ 0.08265f
C3886 _0199_ _0198_ 0
C3887 _0656_/a_59_75# acc0.A\[9\] 0.08314f
C3888 net21 VPWR 2.4232f
C3889 _0993_/a_466_413# net246 0
C3890 _0146_ net218 0
C3891 _0164_ _0487_ 0
C3892 _0461_ net87 0.00702f
C3893 clknet_1_0__leaf__0460_ _0754_/a_512_297# 0
C3894 _0695_/a_472_297# _0219_ 0.00115f
C3895 _0984_/a_634_159# _0984_/a_975_413# 0
C3896 _0984_/a_466_413# _0984_/a_561_413# 0.00772f
C3897 net210 acc0.A\[25\] 0
C3898 _0808_/a_266_47# _0417_ 0.04715f
C3899 _0438_ _0988_/a_193_47# 0
C3900 acc0.A\[9\] _0986_/a_1059_315# 0
C3901 net104 clknet_1_0__leaf__0461_ 0.12588f
C3902 _0550_/a_149_47# _0207_ 0.00154f
C3903 clkbuf_1_0__f__0457_/a_110_47# _0765_/a_79_21# 0
C3904 hold97/a_285_47# _0365_ 0
C3905 clknet_0__0464_ _0147_ 0.01381f
C3906 comp0.B\[5\] hold84/a_285_47# 0
C3907 _1039_/a_975_413# VPWR 0.0049f
C3908 _0730_/a_79_21# VPWR 0.43998f
C3909 _0986_/a_381_47# _0986_/a_561_413# 0.00123f
C3910 _0986_/a_891_413# _0986_/a_975_413# 0.00851f
C3911 net168 _1054_/a_27_47# 0.10133f
C3912 net148 net73 0.08469f
C3913 clknet_0__0458_ _0269_ 0.05645f
C3914 _1017_/a_1017_47# _0181_ 0.002f
C3915 _1023_/a_466_413# net109 0
C3916 _1023_/a_634_159# net177 0.01184f
C3917 _0118_ _0713_/a_27_47# 0.00121f
C3918 _1037_/a_634_159# _0175_ 0
C3919 _0371_ acc0.A\[24\] 0
C3920 hold25/a_285_47# _0176_ 0.03931f
C3921 _0796_/a_79_21# net5 0
C3922 _0753_/a_79_21# _0227_ 0
C3923 clknet_1_0__leaf__0458_ hold18/a_391_47# 0.0109f
C3924 _0337_ _0723_/a_27_413# 0
C3925 _0662_/a_384_47# VPWR 0
C3926 pp[9] acc0.A\[11\] 0.01025f
C3927 _1051_/a_466_413# _0142_ 0
C3928 net16 _0190_ 0.13094f
C3929 hold58/a_49_47# clknet_1_1__leaf__0463_ 0.01639f
C3930 control0.state\[0\] _0946_/a_184_297# 0
C3931 net34 _0946_/a_30_53# 0.29439f
C3932 _0080_ acc0.A\[15\] 0
C3933 VPWR hold4/a_391_47# 0.16309f
C3934 _1045_/a_975_413# net20 0.00107f
C3935 _0834_/a_109_297# _0186_ 0
C3936 _1037_/a_466_413# control0.sh 0.00101f
C3937 net215 acc0.A\[23\] 0.00397f
C3938 hold55/a_49_47# _0181_ 0.00267f
C3939 _0718_/a_285_47# hold62/a_285_47# 0
C3940 _0763_/a_109_47# _0384_ 0.01083f
C3941 _0644_/a_47_47# _0302_ 0.00185f
C3942 _0682_/a_68_297# _0359_ 0.00108f
C3943 _1036_/a_1017_47# comp0.B\[4\] 0
C3944 _0414_ _0346_ 0
C3945 _0466_ _1064_/a_1017_47# 0
C3946 net163 _1031_/a_27_47# 0.10134f
C3947 net133 _0531_/a_109_47# 0
C3948 _0129_ _1031_/a_634_159# 0
C3949 _0368_ _0324_ 0.05142f
C3950 _0616_/a_78_199# _0616_/a_215_47# 0.09071f
C3951 net208 hold61/a_391_47# 0.1341f
C3952 _0340_ _0195_ 0.02635f
C3953 _0404_ _0091_ 0.00279f
C3954 net64 hold31/a_285_47# 0.08884f
C3955 _1059_/a_634_159# net229 0.00279f
C3956 hold31/a_391_47# _0621_/a_35_297# 0
C3957 hold22/a_49_47# _0252_ 0
C3958 hold22/a_391_47# acc0.A\[7\] 0.06996f
C3959 _0417_ _0345_ 0.00476f
C3960 _1012_/a_466_413# _0218_ 0
C3961 hold42/a_49_47# _0156_ 0
C3962 _0196_ clknet_1_1__leaf__0464_ 0
C3963 _0234_ net51 0.18085f
C3964 _0476_ _0210_ 0.03504f
C3965 _1038_/a_193_47# _1037_/a_891_413# 0
C3966 _1038_/a_466_413# _1037_/a_466_413# 0
C3967 _0257_ _0835_/a_292_297# 0
C3968 control0.state\[2\] _0477_ 0.00571f
C3969 _0981_/a_373_47# _0466_ 0.00151f
C3970 clknet_1_0__leaf__0458_ _0195_ 0.00696f
C3971 _0998_/a_634_159# _0796_/a_79_21# 0
C3972 net101 _1020_/a_891_413# 0
C3973 _0997_/a_561_413# _0407_ 0
C3974 _0997_/a_634_159# _0095_ 0
C3975 _0574_/a_27_297# net110 0
C3976 hold99/a_49_47# net246 0.00134f
C3977 _0347_ _0738_/a_68_297# 0.01851f
C3978 net240 _0163_ 0
C3979 _0852_/a_117_297# _0264_ 0.00369f
C3980 hold24/a_49_47# _0176_ 0
C3981 _0236_ control0.add 0
C3982 _0743_/a_245_297# net237 0.00143f
C3983 _0770_/a_297_47# clknet_1_0__leaf__0457_ 0
C3984 _1065_/a_27_47# _1065_/a_634_159# 0.13601f
C3985 _1054_/a_592_47# net11 0
C3986 _0217_ _0760_/a_47_47# 0.01717f
C3987 net232 _1066_/a_193_47# 0.26549f
C3988 hold30/a_49_47# _0120_ 0
C3989 hold30/a_391_47# _0183_ 0.0611f
C3990 _0787_/a_80_21# _0281_ 0.07232f
C3991 _0571_/a_27_297# _0125_ 0.10885f
C3992 _0571_/a_373_47# acc0.A\[27\] 0.00266f
C3993 _0216_ _0199_ 0
C3994 _1036_/a_27_47# _1035_/a_27_47# 0.00268f
C3995 _0259_ _0293_ 0.08548f
C3996 _0584_/a_27_297# clknet_1_0__leaf__0461_ 0.07817f
C3997 clkbuf_1_1__f__0463_/a_110_47# _0956_/a_32_297# 0.01334f
C3998 hold85/a_391_47# net1 0
C3999 net200 _0682_/a_68_297# 0
C4000 VPWR _0261_ 0.8439f
C4001 _0714_/a_240_47# net162 0
C4002 net48 hold4/a_391_47# 0.00142f
C4003 _1033_/a_1059_315# _0565_/a_51_297# 0.00144f
C4004 _0743_/a_240_47# _0219_ 0.03122f
C4005 _0954_/a_32_297# _1042_/a_27_47# 0
C4006 _0637_/a_139_47# acc0.A\[15\] 0
C4007 _0195_ _1013_/a_381_47# 0.00486f
C4008 net169 _0252_ 0
C4009 net27 _1066_/a_1059_315# 0
C4010 VPWR _0957_/a_114_297# 0.00508f
C4011 clknet_0__0463_ net119 0
C4012 output55/a_27_47# output59/a_27_47# 0
C4013 clknet_1_0__leaf__0464_ net135 0.69469f
C4014 B[3] net26 0.00328f
C4015 input5/a_75_212# acc0.A\[13\] 0.00108f
C4016 VPWR _0582_/a_109_47# 0
C4017 net144 net38 0
C4018 _0362_ clknet_0__0460_ 0
C4019 net70 net77 0.00307f
C4020 _0195_ acc0.A\[16\] 0.05081f
C4021 hold38/a_391_47# net119 0
C4022 VPWR _1007_/a_634_159# 0.21281f
C4023 _0399_ _0989_/a_193_47# 0
C4024 _0710_/a_109_297# _0339_ 0.01005f
C4025 _0172_ _1040_/a_1059_315# 0
C4026 _1058_/a_1059_315# VPWR 0.39592f
C4027 _0179_ _1051_/a_193_47# 0.02574f
C4028 _0966_/a_27_47# net167 0
C4029 _0377_ net241 0.15217f
C4030 _0982_/a_1017_47# _0181_ 0
C4031 _0399_ _0992_/a_193_47# 0
C4032 _0262_ _0630_/a_109_297# 0.01483f
C4033 _0493_/a_27_47# _0173_ 0.10379f
C4034 _0992_/a_1017_47# _0283_ 0
C4035 _0307_ net219 0
C4036 _0448_ _0350_ 0.04177f
C4037 _0669_/a_183_297# _0345_ 0
C4038 _1064_/a_634_159# _1064_/a_592_47# 0
C4039 hold78/a_49_47# _0345_ 0
C4040 _0728_/a_145_75# _0345_ 0.00116f
C4041 clknet_1_0__leaf__0458_ _0852_/a_35_297# 0.00494f
C4042 _0441_ _0256_ 0.00486f
C4043 _0440_ _0271_ 0
C4044 hold34/a_285_47# _0512_/a_109_297# 0
C4045 _1015_/a_1059_315# net23 0.03063f
C4046 _0218_ net98 0
C4047 _0402_ acc0.A\[11\] 0
C4048 clkbuf_0_clk/a_110_47# _0166_ 0.00291f
C4049 clknet_1_1__leaf__0465_ _0988_/a_193_47# 0
C4050 _1000_/a_193_47# net219 0
C4051 _0197_ _0446_ 0
C4052 clknet_1_1__leaf_clk _1063_/a_466_413# 0
C4053 _0827_/a_109_297# _0434_ 0.01099f
C4054 _0707_/a_208_47# _0334_ 0
C4055 _1047_/a_381_47# _0171_ 0
C4056 net33 _1065_/a_193_47# 0
C4057 _0255_ _0434_ 0.00691f
C4058 _0440_ _0987_/a_891_413# 0.00102f
C4059 _0346_ _0300_ 0
C4060 net172 net171 0.00315f
C4061 _0672_/a_510_47# _0301_ 0.00225f
C4062 _0644_/a_47_47# net6 0
C4063 _0472_ _0171_ 0
C4064 _0786_/a_472_297# VPWR 0.00623f
C4065 _0280_ _0716_/a_27_47# 0.00311f
C4066 hold78/a_391_47# _0712_/a_79_21# 0
C4067 hold78/a_285_47# _0712_/a_297_297# 0.00151f
C4068 _0770_/a_297_47# _1001_/a_1059_315# 0
C4069 _1004_/a_193_47# net93 0.00159f
C4070 comp0.B\[14\] net198 0
C4071 input6/a_75_212# _0218_ 0
C4072 clkbuf_1_0__f__0459_/a_110_47# _1060_/a_634_159# 0.01307f
C4073 output57/a_27_47# pp[29] 0.15767f
C4074 _0386_ _0310_ 0
C4075 net137 _0524_/a_373_47# 0
C4076 _0427_ _0399_ 0
C4077 _1002_/a_466_413# _0369_ 0
C4078 _0752_/a_384_47# _0227_ 0
C4079 _0343_ _1017_/a_891_413# 0.00299f
C4080 _1056_/a_634_159# _1056_/a_975_413# 0
C4081 VPWR _0509_/a_27_47# 0.30031f
C4082 _0343_ net146 0
C4083 net125 _0175_ 0
C4084 control0.state\[0\] _0967_/a_297_297# 0.00629f
C4085 net34 _0967_/a_109_93# 0
C4086 control0.state\[1\] _0967_/a_215_297# 0.00591f
C4087 _0399_ hold60/a_285_47# 0.11533f
C4088 net34 _0487_ 0.22028f
C4089 control0.state\[0\] _0162_ 0.09928f
C4090 _0985_/a_27_47# net61 0
C4091 _0512_/a_27_297# _0510_/a_27_297# 0
C4092 _1013_/a_27_47# _0339_ 0
C4093 net43 _0347_ 0.01146f
C4094 _0596_/a_59_75# _0222_ 0
C4095 net39 net80 0.11364f
C4096 clknet_1_0__leaf__0458_ _0081_ 0.00425f
C4097 _0664_/a_382_297# _0281_ 0
C4098 _0284_ _0806_/a_113_297# 0
C4099 _0312_ net52 0.04076f
C4100 _1017_/a_1059_315# acc0.A\[17\] 0.08321f
C4101 net154 acc0.A\[6\] 0
C4102 net172 net24 0
C4103 _0857_/a_27_47# _0215_ 0.01593f
C4104 output67/a_27_47# clknet_1_1__leaf__0465_ 0
C4105 _1008_/a_466_413# _0345_ 0
C4106 _0360_ _0321_ 0.5721f
C4107 _0118_ _0579_/a_109_297# 0.00169f
C4108 _0129_ _0345_ 0
C4109 hold16/a_285_47# _0219_ 0
C4110 _0963_/a_35_297# _1070_/a_891_413# 0
C4111 _0854_/a_79_21# _0454_ 0.05483f
C4112 clkbuf_0__0460_/a_110_47# _0360_ 0
C4113 _0350_ _0444_ 0
C4114 hold56/a_285_47# clkbuf_1_1__f__0463_/a_110_47# 0
C4115 clkbuf_1_1__f_clk/a_110_47# _1063_/a_1059_315# 0
C4116 _0226_ _0235_ 0.07301f
C4117 _0322_ _0323_ 0
C4118 _0999_/a_27_47# _0347_ 0.00628f
C4119 net198 _0543_/a_68_297# 0
C4120 _0413_ _0997_/a_27_47# 0
C4121 hold63/a_285_47# net112 0.01848f
C4122 _0498_/a_51_297# _0498_/a_245_297# 0.01218f
C4123 _0088_ clknet_1_1__leaf__0458_ 0
C4124 hold36/a_49_47# _0143_ 0.04371f
C4125 _0830_/a_79_21# _0437_ 0.07744f
C4126 hold6/a_391_47# net153 0.13101f
C4127 _0245_ _0242_ 0.01857f
C4128 _0246_ acc0.A\[19\] 0
C4129 _0118_ _0399_ 0
C4130 _0227_ _0250_ 0
C4131 _0787_/a_303_47# VPWR 0.00405f
C4132 _0323_ _0327_ 0.00805f
C4133 _0199_ net247 0.02346f
C4134 net1 _0958_/a_109_47# 0.00186f
C4135 _0343_ pp[3] 0.00308f
C4136 _0179_ _0514_/a_373_47# 0
C4137 clknet_1_0__leaf__0465_ _1052_/a_381_47# 0.00102f
C4138 _0195_ _0532_/a_299_297# 0.07727f
C4139 _1037_/a_975_413# VPWR 0.00485f
C4140 _0557_/a_51_297# _0557_/a_149_47# 0.02487f
C4141 _0439_ net47 0
C4142 _0577_/a_27_297# _1005_/a_27_47# 0
C4143 _0465_ acc0.A\[6\] 0.00109f
C4144 net65 _0827_/a_27_47# 0
C4145 _0255_ acc0.A\[7\] 0.00862f
C4146 VPWR net47 2.49452f
C4147 acc0.A\[16\] _0081_ 0
C4148 _0516_/a_27_297# net142 0.01004f
C4149 _0402_ hold81/a_391_47# 0
C4150 _0367_ _0350_ 0
C4151 hold23/a_285_47# _0179_ 0
C4152 _0489_ _0976_/a_535_374# 0
C4153 net45 _0294_ 0.03777f
C4154 pp[15] _0995_/a_1017_47# 0
C4155 _0183_ _0773_/a_35_297# 0
C4156 hold12/a_49_47# clknet_1_0__leaf__0460_ 0.00908f
C4157 _1048_/a_466_413# _0196_ 0
C4158 _0368_ _0347_ 0
C4159 net26 hold84/a_49_47# 0
C4160 _0222_ _0216_ 0
C4161 hold43/a_285_47# hold44/a_391_47# 0.00144f
C4162 _0512_/a_27_297# _0181_ 0.12023f
C4163 clknet_1_1__leaf_clk _1062_/a_561_413# 0.00178f
C4164 _1018_/a_466_413# _0581_/a_109_297# 0
C4165 _0689_/a_68_297# _0365_ 0
C4166 _0082_ net229 0
C4167 _1060_/a_1017_47# _0185_ 0
C4168 _1008_/a_27_47# _1008_/a_193_47# 0.96639f
C4169 _0976_/a_76_199# _0167_ 0
C4170 _0488_ _1069_/a_466_413# 0
C4171 _0976_/a_505_21# clknet_1_0__leaf_clk 0.05571f
C4172 _0466_ _1069_/a_634_159# 0
C4173 _0352_ _0319_ 0
C4174 hold16/a_49_47# _0129_ 0.30045f
C4175 net1 _0160_ 0
C4176 pp[27] _0707_/a_544_297# 0.00162f
C4177 _1020_/a_634_159# _1020_/a_381_47# 0
C4178 net157 clknet_1_0__leaf__0457_ 0
C4179 hold18/a_49_47# hold18/a_391_47# 0.00188f
C4180 clknet_1_0__leaf__0458_ _1048_/a_193_47# 0
C4181 _0405_ acc0.A\[15\] 0
C4182 _0400_ net42 0.0265f
C4183 _1035_/a_27_47# comp0.B\[3\] 0
C4184 clkbuf_1_0__f__0464_/a_110_47# _1049_/a_634_159# 0.00527f
C4185 _0598_/a_79_21# _0234_ 0
C4186 _0229_ _0752_/a_27_413# 0
C4187 _0820_/a_510_47# net214 0.00164f
C4188 _0747_/a_215_47# clkbuf_1_0__f__0460_/a_110_47# 0.00206f
C4189 _0342_ acc0.A\[30\] 0.00582f
C4190 _0483_ control0.count\[0\] 0.00121f
C4191 _0404_ _0346_ 0.00142f
C4192 _0983_/a_381_47# net47 0.01679f
C4193 _0343_ _0273_ 0.34494f
C4194 _1016_/a_891_413# net43 0
C4195 net64 output47/a_27_47# 0
C4196 _0684_/a_145_75# clknet_1_1__leaf__0460_ 0
C4197 net205 _0176_ 0
C4198 B[13] net20 0.00165f
C4199 _1058_/a_561_413# clknet_1_1__leaf__0465_ 0
C4200 _0217_ _0350_ 0.38553f
C4201 output66/a_27_47# A[9] 0
C4202 _0473_ _0175_ 0
C4203 clknet_1_1__leaf_clk _0213_ 0.00244f
C4204 pp[27] pp[29] 0
C4205 _0747_/a_215_47# _0250_ 0.04878f
C4206 _0199_ _1048_/a_466_413# 0
C4207 _0998_/a_193_47# _1017_/a_891_413# 0
C4208 _0998_/a_381_47# _1017_/a_27_47# 0
C4209 _1013_/a_193_47# net99 0.00453f
C4210 net9 _0186_ 0.0693f
C4211 _0411_ _0297_ 0.00765f
C4212 clkbuf_1_0__f__0459_/a_110_47# _0115_ 0
C4213 _1001_/a_975_413# net46 0
C4214 _0313_ _0741_/a_109_297# 0
C4215 _0683_/a_113_47# _0315_ 0.01004f
C4216 _1041_/a_27_47# net30 0
C4217 _0388_ _0768_/a_109_297# 0
C4218 _0349_ hold95/a_285_47# 0.05679f
C4219 _1003_/a_381_47# _0466_ 0
C4220 comp0.B\[15\] acc0.A\[15\] 0.02152f
C4221 output56/a_27_47# _0195_ 0.01527f
C4222 net227 hold80/a_49_47# 0
C4223 _0399_ net142 0
C4224 acc0.A\[30\] _0334_ 0
C4225 _0645_/a_47_47# net41 0.40239f
C4226 _0243_ clknet_1_0__leaf__0461_ 0.19726f
C4227 _0826_/a_219_297# _0826_/a_27_53# 0.10125f
C4228 _0176_ _0540_/a_240_47# 0
C4229 clknet_1_0__leaf__0462_ _0752_/a_27_413# 0
C4230 pp[17] _0220_ 0.18168f
C4231 _0992_/a_193_47# _0295_ 0
C4232 _0982_/a_27_47# _0855_/a_81_21# 0.00185f
C4233 _0144_ _1049_/a_193_47# 0
C4234 _0536_/a_51_297# _0147_ 0
C4235 _1036_/a_891_413# net24 0
C4236 clkload1/a_268_47# clkload1/Y 0.00587f
C4237 _0274_ _0824_/a_59_75# 0.00958f
C4238 _1058_/a_27_47# _1057_/a_634_159# 0
C4239 _1058_/a_193_47# _1057_/a_193_47# 0.02521f
C4240 _1058_/a_634_159# _1057_/a_27_47# 0
C4241 _0307_ _0352_ 0.02587f
C4242 _0412_ _0411_ 0.11897f
C4243 _0311_ _0238_ 0.11981f
C4244 _0369_ net37 0
C4245 _0464_ _1061_/a_1059_315# 0.03246f
C4246 _0534_/a_384_47# clknet_1_1__leaf__0457_ 0.00108f
C4247 acc0.A\[7\] A[7] 0.0012f
C4248 _0294_ _0990_/a_1059_315# 0
C4249 control0.count\[1\] control0.count\[0\] 0.98666f
C4250 net35 hold17/a_391_47# 0
C4251 net104 _0218_ 0.00141f
C4252 _1000_/a_1059_315# _0347_ 0
C4253 _1000_/a_193_47# _0352_ 0.05112f
C4254 VPWR _1063_/a_1059_315# 0.4069f
C4255 net101 _0346_ 0
C4256 _0611_/a_68_297# _0611_/a_150_297# 0.00477f
C4257 net86 _0245_ 0.01903f
C4258 _0572_/a_109_297# _0124_ 0.00467f
C4259 _0572_/a_373_47# _0216_ 0
C4260 VPWR _0959_/a_80_21# 0.25417f
C4261 _0216_ _1006_/a_592_47# 0
C4262 _0616_/a_78_199# _0771_/a_215_297# 0.00188f
C4263 hold47/a_391_47# net135 0.00116f
C4264 VPWR net159 0.28268f
C4265 output46/a_27_47# net51 0
C4266 net46 output51/a_27_47# 0.00311f
C4267 _0453_ _0261_ 0
C4268 clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ 1.67439f
C4269 net190 hold9/a_285_47# 0.04421f
C4270 _0839_/a_109_297# _0444_ 0.01262f
C4271 _0275_ _0268_ 0
C4272 _1052_/a_1059_315# acc0.A\[8\] 0
C4273 _0984_/a_193_47# net229 0
C4274 hold55/a_391_47# net118 0
C4275 VPWR _1060_/a_1059_315# 0.41387f
C4276 _1019_/a_1059_315# acc0.A\[19\] 0.08367f
C4277 _0419_ _0091_ 0.03894f
C4278 pp[28] _0707_/a_201_297# 0.00956f
C4279 _0385_ _0369_ 0
C4280 hold84/a_49_47# hold84/a_285_47# 0.22264f
C4281 clknet_0__0457_ _0385_ 0.00213f
C4282 _0609_/a_109_297# VPWR 0.00427f
C4283 net2 acc0.A\[10\] 0.02681f
C4284 VPWR _0988_/a_592_47# 0
C4285 _1044_/a_27_47# _0542_/a_240_47# 0
C4286 _0499_/a_145_75# _0171_ 0.00256f
C4287 _1054_/a_891_413# _0186_ 0.00374f
C4288 pp[10] VPWR 0.82667f
C4289 _0791_/a_199_47# _0219_ 0.00154f
C4290 _0786_/a_472_297# _0283_ 0.00612f
C4291 net61 _0197_ 0
C4292 hold75/a_391_47# net58 0.08254f
C4293 _0342_ _0779_/a_79_21# 0
C4294 net157 _1047_/a_891_413# 0.00983f
C4295 _0195_ _0247_ 0
C4296 clknet_0_clk _0974_/a_79_199# 0.00344f
C4297 clknet_1_0__leaf__0463_ A[1] 0.01731f
C4298 _0311_ _0767_/a_145_75# 0
C4299 net109 net177 0.00256f
C4300 _1023_/a_1017_47# acc0.A\[23\] 0
C4301 hold89/a_49_47# control0.state\[2\] 0.36394f
C4302 _0247_ net92 0
C4303 net149 _0171_ 0
C4304 hold45/a_391_47# _0511_/a_81_21# 0
C4305 hold45/a_285_47# _0511_/a_299_297# 0
C4306 net82 _0996_/a_193_47# 0.01325f
C4307 _0619_/a_68_297# _0989_/a_193_47# 0
C4308 clknet_1_0__leaf__0462_ clknet_1_1__leaf__0460_ 0.00122f
C4309 _1031_/a_193_47# clknet_1_1__leaf__0462_ 0
C4310 _0732_/a_303_47# _0324_ 0
C4311 pp[27] _1010_/a_193_47# 0
C4312 net59 _0351_ 0
C4313 hold59/a_285_47# _0853_/a_68_297# 0
C4314 _0149_ _0142_ 0
C4315 _0322_ _0686_/a_27_53# 0.00282f
C4316 _0183_ hold71/a_285_47# 0
C4317 _0216_ acc0.A\[27\] 0.21723f
C4318 _0476_ _0467_ 0.02755f
C4319 clknet_1_0__leaf__0465_ _0440_ 0.07208f
C4320 _0457_ _1015_/a_381_47# 0.01017f
C4321 net183 _0172_ 0.07741f
C4322 _0322_ _1008_/a_891_413# 0
C4323 _0329_ _1008_/a_1059_315# 0
C4324 _0331_ _0318_ 0
C4325 _0402_ _0281_ 0.8478f
C4326 _0135_ control0.sh 0.0436f
C4327 _0327_ _0686_/a_27_53# 0.00238f
C4328 _1037_/a_891_413# net29 0
C4329 _1037_/a_381_47# B[6] 0
C4330 comp0.B\[6\] control0.reset 0
C4331 clknet_1_0__leaf__0459_ net47 0
C4332 _0326_ _0618_/a_79_21# 0
C4333 _0248_ _0350_ 0.10765f
C4334 net45 _1017_/a_561_413# 0
C4335 net78 _0179_ 0
C4336 _0179_ clknet_0__0465_ 0
C4337 VPWR _1062_/a_975_413# 0.00417f
C4338 net145 net229 0.21371f
C4339 _1018_/a_193_47# _0347_ 0.00359f
C4340 _0849_/a_215_47# acc0.A\[15\] 0.00395f
C4341 _0324_ clknet_0__0460_ 0
C4342 _1039_/a_891_413# _0137_ 0.04696f
C4343 _1021_/a_381_47# VPWR 0.07784f
C4344 net189 _0156_ 0.00146f
C4345 pp[29] _0216_ 0
C4346 _1038_/a_466_413# _0135_ 0
C4347 net172 _1037_/a_466_413# 0
C4348 _0178_ net201 0
C4349 acc0.A\[1\] _0580_/a_109_47# 0
C4350 _0762_/a_79_21# _0383_ 0.09503f
C4351 _0762_/a_215_47# _0369_ 0.08609f
C4352 _0481_ _0961_/a_199_47# 0
C4353 _0343_ hold88/a_285_47# 0.01086f
C4354 _0279_ _0647_/a_129_47# 0
C4355 _0753_/a_79_21# _0352_ 0
C4356 _0106_ _0738_/a_68_297# 0.00466f
C4357 _0476_ comp0.B\[0\] 0.00675f
C4358 _0984_/a_1059_315# clkbuf_1_0__f__0458_/a_110_47# 0.02221f
C4359 _1011_/a_27_47# _0332_ 0.01789f
C4360 net36 _1061_/a_27_47# 0
C4361 _0195_ _0455_ 0
C4362 pp[10] input4/a_75_212# 0.00432f
C4363 hold14/a_391_47# _0175_ 0.00238f
C4364 _0579_/a_27_297# acc0.A\[20\] 0
C4365 _1065_/a_891_413# _1065_/a_975_413# 0.00851f
C4366 _1065_/a_381_47# _1065_/a_561_413# 0.00123f
C4367 hold5/a_285_47# _0544_/a_240_47# 0
C4368 VPWR _0173_ 1.98475f
C4369 _0677_/a_129_47# _0347_ 0
C4370 _0183_ _0382_ 0.00284f
C4371 _0592_/a_68_297# _1022_/a_891_413# 0
C4372 clknet_0_clk _1062_/a_193_47# 0
C4373 _0999_/a_1059_315# net41 0
C4374 _0967_/a_215_297# _1066_/a_634_159# 0
C4375 hold28/a_285_47# VPWR 0.27188f
C4376 hold69/a_285_47# _0460_ 0.00284f
C4377 _0508_/a_81_21# _0185_ 0.16682f
C4378 hold66/a_285_47# _1005_/a_634_159# 0
C4379 _0817_/a_266_47# _0991_/a_891_413# 0
C4380 _0467_ hold89/a_285_47# 0
C4381 _0746_/a_299_297# net52 0.00112f
C4382 _0520_/a_109_47# net13 0
C4383 _1036_/a_634_159# B[15] 0
C4384 _1068_/a_466_413# _0487_ 0
C4385 _0723_/a_27_413# _0333_ 0
C4386 _0216_ _0110_ 0
C4387 _0707_/a_75_199# _0335_ 0.12168f
C4388 net24 _0474_ 0.02184f
C4389 comp0.B\[12\] _1042_/a_1059_315# 0
C4390 comp0.B\[11\] _1042_/a_891_413# 0.05471f
C4391 _0266_ _0265_ 0.3457f
C4392 _1014_/a_1059_315# _1014_/a_891_413# 0.31086f
C4393 _1014_/a_193_47# _1014_/a_975_413# 0
C4394 _1014_/a_466_413# _1014_/a_381_47# 0.03733f
C4395 _0453_ net47 0.0855f
C4396 _1071_/a_27_47# _1071_/a_466_413# 0.27314f
C4397 _1071_/a_193_47# _1071_/a_634_159# 0.12497f
C4398 acc0.A\[15\] hold71/a_285_47# 0.06889f
C4399 VPWR _1047_/a_1017_47# 0
C4400 _0996_/a_634_159# _0796_/a_79_21# 0.00153f
C4401 output59/a_27_47# acc0.A\[30\] 0
C4402 pp[30] _0704_/a_150_297# 0
C4403 _0343_ _0086_ 0
C4404 net36 hold60/a_391_47# 0
C4405 _1015_/a_27_47# _0208_ 0.11616f
C4406 _1015_/a_466_413# _0173_ 0
C4407 clknet_1_0__leaf__0460_ acc0.A\[23\] 0.10397f
C4408 pp[9] A[12] 0.2503f
C4409 _0816_/a_68_297# _0347_ 0.02422f
C4410 _0985_/a_1059_315# _0458_ 0.01972f
C4411 VPWR net93 0.55055f
C4412 _0343_ _0226_ 0
C4413 _0458_ _1049_/a_193_47# 0
C4414 _0217_ _0244_ 0.0071f
C4415 VPWR input17/a_75_212# 0.2664f
C4416 _0179_ net184 0
C4417 _0564_/a_68_297# _0161_ 0
C4418 clkbuf_0__0461_/a_110_47# _0115_ 0.00133f
C4419 _0617_/a_68_297# _0460_ 0.0125f
C4420 _0572_/a_27_297# _1026_/a_27_47# 0
C4421 clknet_0__0458_ clkbuf_0__0458_/a_110_47# 1.67884f
C4422 VPWR _0536_/a_512_297# 0.00729f
C4423 clknet_1_0__leaf__0463_ clkbuf_0__0463_/a_110_47# 0.00391f
C4424 VPWR _0796_/a_510_47# 0
C4425 comp0.B\[12\] net10 0
C4426 pp[28] _1010_/a_27_47# 0
C4427 _1039_/a_891_413# comp0.B\[6\] 0
C4428 hold13/a_285_47# _0175_ 0
C4429 _0717_/a_209_47# _0334_ 0.00209f
C4430 _0252_ _0830_/a_79_21# 0
C4431 net65 _0830_/a_510_47# 0.00528f
C4432 acc0.A\[7\] _0830_/a_215_47# 0
C4433 _0305_ _1059_/a_193_47# 0.01852f
C4434 _0499_/a_59_75# control0.sh 0.21271f
C4435 clkbuf_1_0__f__0459_/a_110_47# _1017_/a_891_413# 0
C4436 net45 _0581_/a_109_297# 0.00249f
C4437 hold63/a_285_47# net111 0.00611f
C4438 VPWR _0848_/a_109_297# 0.00389f
C4439 clknet_1_1__leaf_clk _0161_ 0.06473f
C4440 _0442_ _0085_ 0
C4441 VPWR _0547_/a_150_297# 0.00144f
C4442 _0454_ _0852_/a_117_297# 0
C4443 net2 _0510_/a_109_297# 0.01008f
C4444 net168 _0523_/a_299_297# 0
C4445 _0455_ _0852_/a_35_297# 0
C4446 _0341_ pp[31] 0.00542f
C4447 _1026_/a_891_413# acc0.A\[25\] 0.00204f
C4448 net36 _1039_/a_27_47# 0.44712f
C4449 _0462_ clknet_1_0__leaf__0457_ 0.04221f
C4450 net88 _1067_/a_27_47# 0
C4451 hold78/a_285_47# _0344_ 0
C4452 _1012_/a_634_159# _0347_ 0.00834f
C4453 output54/a_27_47# hold9/a_285_47# 0
C4454 _0290_ _0658_/a_113_47# 0.00992f
C4455 clkbuf_1_0__f__0459_/a_110_47# net146 0
C4456 hold67/a_391_47# net66 0.04085f
C4457 hold67/a_285_47# acc0.A\[8\] 0
C4458 net160 _0176_ 0.3853f
C4459 _0100_ _0369_ 0.13052f
C4460 VPWR _0294_ 2.30611f
C4461 hold13/a_391_47# control0.sh 0
C4462 _0183_ _1059_/a_891_413# 0
C4463 _0343_ _1016_/a_193_47# 0.00998f
C4464 clknet_1_0__leaf__0462_ _0233_ 0
C4465 clknet_1_0__leaf__0462_ _0575_/a_109_297# 0.00465f
C4466 hold75/a_49_47# _0263_ 0.01455f
C4467 _0504_/a_27_47# net149 0.00112f
C4468 _0831_/a_117_297# acc0.A\[6\] 0.00361f
C4469 _0512_/a_27_297# _0187_ 0
C4470 _0216_ _1010_/a_193_47# 0
C4471 clknet_0__0463_ _0463_ 0.52854f
C4472 _0981_/a_109_297# _0490_ 0.01066f
C4473 _0981_/a_27_297# net167 0.16195f
C4474 hold15/a_285_47# _0341_ 0.0011f
C4475 hold15/a_49_47# _0340_ 0
C4476 _0092_ _0647_/a_47_47# 0
C4477 clknet_1_0__leaf__0459_ _1060_/a_1059_315# 0.0019f
C4478 _1052_/a_193_47# _0180_ 0.02901f
C4479 _0275_ _0991_/a_466_413# 0
C4480 _1016_/a_27_47# acc0.A\[17\] 0
C4481 _0254_ acc0.A\[6\] 0.19272f
C4482 net247 _0449_ 0
C4483 _0222_ _1022_/a_592_47# 0
C4484 _0456_ net149 0.01599f
C4485 _0963_/a_285_297# _0168_ 0
C4486 _0455_ _0081_ 0
C4487 _0500_/a_27_47# _0182_ 0.00269f
C4488 _1037_/a_1059_315# _1036_/a_1059_315# 0
C4489 _1037_/a_466_413# _1036_/a_891_413# 0
C4490 _0602_/a_113_47# clknet_1_0__leaf__0460_ 0
C4491 _0179_ hold71/a_285_47# 0
C4492 _0571_/a_109_297# _1026_/a_1059_315# 0
C4493 _0571_/a_27_297# _1026_/a_891_413# 0
C4494 hold42/a_49_47# output37/a_27_47# 0.02146f
C4495 _0553_/a_512_297# net29 0
C4496 _0223_ _0366_ 0.00118f
C4497 hold23/a_391_47# _0530_/a_299_297# 0
C4498 _0279_ clkbuf_1_1__f__0459_/a_110_47# 0
C4499 _0346_ _0419_ 0.04729f
C4500 _0869_/a_27_47# acc0.A\[18\] 0
C4501 _0459_ _0612_/a_59_75# 0.01245f
C4502 _0999_/a_975_413# _0352_ 0
C4503 _1013_/a_891_413# pp[31] 0
C4504 _0498_/a_149_47# net247 0.00877f
C4505 net22 _0546_/a_512_297# 0.0021f
C4506 _0445_ _0986_/a_193_47# 0.00306f
C4507 _0595_/a_109_297# VPWR 0.00604f
C4508 hold29/a_391_47# net51 0
C4509 net182 net47 0
C4510 _0399_ _0988_/a_27_47# 0
C4511 _1038_/a_193_47# _0136_ 0
C4512 net172 _0553_/a_51_297# 0
C4513 comp0.B\[2\] _1033_/a_381_47# 0.02112f
C4514 net150 _1005_/a_891_413# 0
C4515 _0217_ _1005_/a_1059_315# 0
C4516 clkload1/a_110_47# _0257_ 0
C4517 _0126_ _1028_/a_466_413# 0
C4518 _0570_/a_109_297# net114 0
C4519 net190 _1028_/a_381_47# 0.02284f
C4520 _0949_/a_145_75# net231 0
C4521 hold46/a_391_47# VPWR 0.20188f
C4522 pp[28] pp[30] 0
C4523 _0316_ clknet_0__0460_ 0.08946f
C4524 _0180_ net12 0.27665f
C4525 _1032_/a_27_47# _0565_/a_51_297# 0
C4526 _0955_/a_32_297# _0561_/a_149_47# 0
C4527 net55 net98 0
C4528 VPWR input5/a_75_212# 0.26455f
C4529 pp[9] _1057_/a_193_47# 0
C4530 hold67/a_391_47# _0350_ 0.05655f
C4531 _0190_ net142 0.00546f
C4532 _1022_/a_27_47# _1022_/a_193_47# 0.9743f
C4533 acc0.A\[31\] _1013_/a_193_47# 0
C4534 _0576_/a_109_297# acc0.A\[23\] 0.01958f
C4535 _0441_ clknet_0__0465_ 0
C4536 _1003_/a_891_413# clknet_1_0__leaf__0460_ 0.00424f
C4537 _1021_/a_193_47# _0462_ 0
C4538 _0462_ hold90/a_391_47# 0.00433f
C4539 _1059_/a_891_413# acc0.A\[15\] 0.00603f
C4540 _0717_/a_209_297# pp[27] 0.00471f
C4541 VPWR _0775_/a_297_297# 0.01166f
C4542 net118 _0352_ 0
C4543 clknet_0__0460_ _0347_ 0
C4544 clkbuf_1_0__f__0460_/a_110_47# _0352_ 0.04263f
C4545 hold20/a_49_47# VPWR 0.31058f
C4546 _0663_/a_297_47# _0179_ 0
C4547 control0.sh _0160_ 0.00272f
C4548 _1018_/a_1059_315# _0116_ 0.00938f
C4549 _1018_/a_561_413# net206 0
C4550 _0579_/a_109_297# _1001_/a_27_47# 0
C4551 _0339_ _0704_/a_150_297# 0
C4552 _1008_/a_466_413# _1008_/a_592_47# 0.00553f
C4553 _1008_/a_634_159# _1008_/a_1017_47# 0
C4554 _1055_/a_634_159# _1055_/a_466_413# 0.23992f
C4555 _1055_/a_193_47# _1055_/a_1059_315# 0.03405f
C4556 _1055_/a_27_47# _1055_/a_891_413# 0.03224f
C4557 _0488_ _0167_ 0
C4558 _0466_ clknet_1_0__leaf_clk 1.25568f
C4559 _0349_ _1011_/a_193_47# 0
C4560 pp[16] _0995_/a_466_413# 0
C4561 _1020_/a_891_413# _0118_ 0.04718f
C4562 net53 _1025_/a_381_47# 0.00113f
C4563 pp[25] _1025_/a_1059_315# 0
C4564 _0250_ _0352_ 0.14633f
C4565 pp[18] _0218_ 0
C4566 _0559_/a_245_297# _0173_ 0.00175f
C4567 _0215_ _0208_ 0.002f
C4568 _0175_ _0132_ 0
C4569 _1003_/a_193_47# _1003_/a_634_159# 0.11072f
C4570 _1003_/a_27_47# _1003_/a_466_413# 0.27314f
C4571 net2 _0188_ 0
C4572 _0999_/a_634_159# _0408_ 0
C4573 net166 _0583_/a_109_297# 0.00117f
C4574 _1055_/a_634_159# net181 0
C4575 _0750_/a_109_47# net48 0
C4576 _0243_ _0218_ 0.26776f
C4577 net232 VPWR 0.53287f
C4578 _0292_ _0508_/a_299_297# 0
C4579 clknet_0__0458_ _0986_/a_975_413# 0
C4580 _0244_ _0248_ 0
C4581 net114 hold50/a_285_47# 0.04611f
C4582 hold58/a_49_47# hold58/a_285_47# 0.22264f
C4583 _0176_ _0542_/a_512_297# 0
C4584 net84 _1017_/a_1059_315# 0.00169f
C4585 net46 _0391_ 0.02261f
C4586 _0275_ _0401_ 0.57368f
C4587 _1032_/a_381_47# comp0.B\[0\] 0
C4588 VPWR _0690_/a_68_297# 0.13808f
C4589 _0997_/a_634_159# _0219_ 0.00633f
C4590 _0997_/a_381_47# _0345_ 0.00537f
C4591 _0266_ _0267_ 0.08534f
C4592 _0833_/a_297_297# _0439_ 0
C4593 net63 _0433_ 0.42765f
C4594 _1004_/a_891_413# _0758_/a_79_21# 0.00145f
C4595 _0992_/a_1017_47# _0345_ 0
C4596 VPWR _0833_/a_297_297# 0.00738f
C4597 pp[12] VPWR 0.39088f
C4598 hold75/a_285_47# net47 0
C4599 net197 _0739_/a_510_47# 0
C4600 net203 _1034_/a_193_47# 0
C4601 _0307_ hold72/a_285_47# 0.00105f
C4602 _0837_/a_585_47# acc0.A\[5\] 0
C4603 _1054_/a_193_47# _1053_/a_193_47# 0.00194f
C4604 _0221_ hold61/a_391_47# 0
C4605 net236 clknet_1_0__leaf_clk 0.03055f
C4606 net102 net221 0.09972f
C4607 _0982_/a_381_47# net234 0
C4608 comp0.B\[4\] B[1] 0.00321f
C4609 _0176_ acc0.A\[15\] 0.08869f
C4610 _0299_ _0668_/a_297_47# 0.01567f
C4611 _0951_/a_109_93# _0468_ 0
C4612 _0218_ _0407_ 0
C4613 _0179_ _1059_/a_891_413# 0
C4614 _0409_ hold91/a_49_47# 0.004f
C4615 _0343_ net41 0.14733f
C4616 _0985_/a_27_47# _0269_ 0
C4617 _1059_/a_193_47# _0181_ 0
C4618 _0924_/a_27_47# net133 0
C4619 _0387_ _0780_/a_35_297# 0.10617f
C4620 _0748_/a_299_297# _0462_ 0
C4621 _0367_ _0737_/a_285_297# 0
C4622 _0315_ _0737_/a_285_47# 0
C4623 hold2/a_391_47# _0465_ 0.01012f
C4624 _1016_/a_381_47# clknet_1_1__leaf__0461_ 0.01471f
C4625 clknet_1_0__leaf_clk _1064_/a_193_47# 0.01548f
C4626 _0330_ hold95/a_391_47# 0
C4627 net211 _0869_/a_27_47# 0.00235f
C4628 _0322_ _0320_ 0.00291f
C4629 _0310_ _0240_ 0.14227f
C4630 VPWR _1017_/a_561_413# 0.00213f
C4631 _1015_/a_193_47# _0178_ 0
C4632 _0717_/a_80_21# pp[28] 0.01113f
C4633 clknet_1_1__leaf__0464_ _0540_/a_51_297# 0
C4634 _0310_ _0369_ 0.02865f
C4635 _0365_ hold50/a_285_47# 0.07824f
C4636 clknet_1_0__leaf__0459_ _0294_ 0.16991f
C4637 net226 _0479_ 0
C4638 _1037_/a_891_413# comp0.B\[6\] 0.00261f
C4639 _1037_/a_381_47# comp0.B\[5\] 0
C4640 VPWR net153 0.43821f
C4641 _0846_/a_51_297# _0844_/a_79_21# 0
C4642 clknet_1_1__leaf__0460_ _0356_ 0.00127f
C4643 _0111_ _0999_/a_1059_315# 0
C4644 _0640_/a_215_297# _0826_/a_219_297# 0
C4645 pp[28] _0339_ 0.20538f
C4646 _0399_ _0459_ 0.00905f
C4647 _1017_/a_891_413# clkbuf_0__0461_/a_110_47# 0
C4648 _0675_/a_68_297# clknet_0__0461_ 0.02968f
C4649 VPWR _1033_/a_1059_315# 0.40565f
C4650 clknet_1_0__leaf__0464_ _0172_ 0.00359f
C4651 _1038_/a_1059_315# comp0.B\[8\] 0
C4652 clknet_1_1__leaf__0460_ _0574_/a_373_47# 0
C4653 _1044_/a_891_413# net19 0
C4654 clknet_1_0__leaf__0458_ _0183_ 0.04393f
C4655 _0343_ hold62/a_285_47# 0.01903f
C4656 _0429_ _0619_/a_150_297# 0
C4657 _0770_/a_297_47# _0246_ 0
C4658 _0600_/a_103_199# _0618_/a_79_21# 0.00119f
C4659 _0989_/a_27_47# _0434_ 0
C4660 hold86/a_285_47# VPWR 0.25912f
C4661 VPWR _1050_/a_975_413# 0.00468f
C4662 _0329_ clknet_1_1__leaf__0462_ 0.11076f
C4663 _0511_/a_384_47# _0156_ 0
C4664 _0179_ _0519_/a_81_21# 0.04984f
C4665 _0274_ _0432_ 0.08292f
C4666 _0275_ _0443_ 0.02689f
C4667 hold33/a_285_47# net31 0
C4668 _1010_/a_634_159# _1010_/a_381_47# 0
C4669 clknet_1_0__leaf__0462_ _1004_/a_891_413# 0.00664f
C4670 _0628_/a_109_297# _0260_ 0.01216f
C4671 _1056_/a_27_47# _0514_/a_27_297# 0
C4672 _0465_ _0826_/a_219_297# 0
C4673 _0991_/a_891_413# _0181_ 0.00242f
C4674 _1040_/a_27_47# _1040_/a_891_413# 0.02974f
C4675 _1040_/a_193_47# _1040_/a_1059_315# 0.03405f
C4676 _1040_/a_634_159# _1040_/a_466_413# 0.23992f
C4677 _0670_/a_297_297# _0409_ 0
C4678 hold79/a_49_47# _0976_/a_76_199# 0.00854f
C4679 _0305_ _0607_/a_109_47# 0.00253f
C4680 _0472_ _0494_/a_27_47# 0.02128f
C4681 _0146_ _1048_/a_891_413# 0.05721f
C4682 _0697_/a_217_297# _0328_ 0.00651f
C4683 _0432_ _0837_/a_266_47# 0
C4684 _0714_/a_51_297# clknet_1_1__leaf__0459_ 0
C4685 _0195_ _1027_/a_193_47# 0
C4686 net243 _0216_ 0.07778f
C4687 _0662_/a_384_47# _0345_ 0
C4688 _1002_/a_1059_315# _0183_ 0
C4689 _1002_/a_381_47# _0217_ 0.00184f
C4690 hold24/a_49_47# net28 0
C4691 _0385_ _0764_/a_384_47# 0
C4692 B[13] B[9] 0.18789f
C4693 _0372_ _1006_/a_193_47# 0
C4694 _0183_ acc0.A\[16\] 0.21965f
C4695 _0221_ clknet_1_1__leaf__0462_ 0
C4696 clknet_0__0459_ _0280_ 0
C4697 _1020_/a_592_47# _0461_ 0
C4698 _0118_ _0891_/a_27_47# 0.01245f
C4699 acc0.A\[14\] _0996_/a_27_47# 0.00846f
C4700 _0846_/a_51_297# _0846_/a_240_47# 0.03076f
C4701 net45 _1016_/a_466_413# 0
C4702 _1067_/a_634_159# _1067_/a_466_413# 0.23992f
C4703 _1067_/a_193_47# _1067_/a_1059_315# 0.03405f
C4704 _1067_/a_27_47# _1067_/a_891_413# 0.03224f
C4705 net9 _0987_/a_634_159# 0.00211f
C4706 _0968_/a_109_297# _0468_ 0
C4707 net172 _0135_ 0
C4708 _1019_/a_27_47# _1015_/a_193_47# 0
C4709 _1019_/a_193_47# _1015_/a_27_47# 0
C4710 hold31/a_285_47# _0369_ 0
C4711 net180 comp0.B\[10\] 0.02653f
C4712 _1071_/a_27_47# _0480_ 0
C4713 _0231_ _0102_ 0
C4714 _0346_ _0992_/a_193_47# 0
C4715 _0399_ _0265_ 0
C4716 _1000_/a_193_47# _0392_ 0
C4717 _1072_/a_193_47# _1071_/a_1059_315# 0
C4718 _0647_/a_285_47# _0347_ 0
C4719 VPWR _0581_/a_109_297# 0.17739f
C4720 clknet_1_0__leaf__0458_ acc0.A\[15\] 0.61534f
C4721 _0314_ _0368_ 0
C4722 _1009_/a_193_47# _1009_/a_592_47# 0.00128f
C4723 _1009_/a_466_413# _1009_/a_561_413# 0.00772f
C4724 _1009_/a_634_159# _1009_/a_975_413# 0
C4725 _0620_/a_113_47# acc0.A\[7\] 0
C4726 _0482_ _0961_/a_113_297# 0
C4727 _0217_ _0592_/a_68_297# 0
C4728 _0330_ acc0.A\[28\] 0.02031f
C4729 net65 _0989_/a_193_47# 0.03687f
C4730 acc0.A\[7\] _0989_/a_27_47# 0
C4731 acc0.A\[7\] hold1/a_49_47# 0
C4732 _0989_/a_27_47# _0989_/a_1059_315# 0.04875f
C4733 _0989_/a_193_47# _0989_/a_466_413# 0.07482f
C4734 input18/a_75_212# B[10] 0.19732f
C4735 _0645_/a_285_47# _1059_/a_1059_315# 0
C4736 comp0.B\[13\] hold36/a_49_47# 0
C4737 control0.state\[0\] _0950_/a_75_212# 0
C4738 output58/a_27_47# _0438_ 0
C4739 net228 _0806_/a_199_47# 0
C4740 comp0.B\[15\] _0565_/a_240_47# 0.01132f
C4741 _0956_/a_114_297# net201 0.00304f
C4742 hold65/a_391_47# acc0.A\[8\] 0
C4743 _0800_/a_512_297# _0218_ 0
C4744 hold18/a_391_47# _0448_ 0
C4745 _0982_/a_561_413# VPWR 0.00297f
C4746 _0476_ _1066_/a_381_47# 0.00695f
C4747 hold66/a_285_47# net91 0
C4748 hold66/a_49_47# _0103_ 0
C4749 _0992_/a_27_47# _0992_/a_1059_315# 0.04875f
C4750 _0992_/a_193_47# _0992_/a_466_413# 0.08301f
C4751 _1036_/a_592_47# net121 0.00149f
C4752 comp0.B\[4\] _1035_/a_891_413# 0.00138f
C4753 net24 _0563_/a_51_297# 0.13504f
C4754 _0498_/a_240_47# _0138_ 0
C4755 _0476_ net1 0.21523f
C4756 _0606_/a_215_297# VPWR 0.15079f
C4757 _0166_ _0487_ 0.02633f
C4758 VPWR _1053_/a_466_413# 0.25244f
C4759 _0607_/a_109_297# net43 0.01173f
C4760 _0427_ _0346_ 0.00302f
C4761 _0125_ _1027_/a_634_159# 0.01128f
C4762 _0718_/a_377_297# pp[27] 0
C4763 acc0.A\[27\] _1027_/a_891_413# 0.01117f
C4764 _0335_ _0338_ 0.17241f
C4765 comp0.B\[1\] net201 0.17533f
C4766 _0280_ _0655_/a_109_93# 0.07433f
C4767 _1032_/a_891_413# net118 0
C4768 _0329_ net242 0
C4769 _0354_ _1029_/a_27_47# 0
C4770 _0959_/a_80_21# comp0.B\[3\] 0
C4771 _1014_/a_466_413# acc0.A\[0\] 0.00156f
C4772 _1014_/a_561_413# net100 0
C4773 _1071_/a_1059_315# _1071_/a_1017_47# 0
C4774 _0996_/a_891_413# _0410_ 0
C4775 _0996_/a_466_413# _0094_ 0.00131f
C4776 _0996_/a_381_47# net238 0.00507f
C4777 clknet_1_1__leaf__0464_ _0524_/a_27_297# 0.01175f
C4778 _0768_/a_27_47# _0240_ 0.01989f
C4779 _0835_/a_292_297# _0218_ 0
C4780 _1000_/a_891_413# clkbuf_1_0__f__0461_/a_110_47# 0.00652f
C4781 _1000_/a_634_159# clknet_0__0461_ 0.00263f
C4782 _0113_ _0173_ 0.00174f
C4783 _0270_ acc0.A\[3\] 0
C4784 _0212_ _1036_/a_193_47# 0
C4785 hold96/a_391_47# net243 0.13105f
C4786 _0261_ _0345_ 0.02314f
C4787 _0346_ hold60/a_285_47# 0.03247f
C4788 _0260_ net247 0.00167f
C4789 clkload4/a_268_47# _0219_ 0
C4790 _0768_/a_27_47# _0369_ 0
C4791 net45 _0714_/a_240_47# 0.00168f
C4792 _0179_ net130 0
C4793 hold54/a_285_47# _0565_/a_51_297# 0.0133f
C4794 _0255_ _0186_ 0.00485f
C4795 net136 net9 0.00959f
C4796 net187 hold40/a_49_47# 0
C4797 acc0.A\[16\] acc0.A\[15\] 0
C4798 _0251_ _0437_ 0.14182f
C4799 _0659_/a_68_297# _0990_/a_27_47# 0.00143f
C4800 hold39/a_285_47# net186 0.00733f
C4801 output49/a_27_47# VPWR 0.31509f
C4802 _0946_/a_184_297# VPWR 0
C4803 net64 _0517_/a_384_47# 0
C4804 _0216_ _1026_/a_634_159# 0.00953f
C4805 _0195_ _1026_/a_1059_315# 0.02869f
C4806 _0124_ _1026_/a_27_47# 0.07487f
C4807 B[15] B[3] 0.01396f
C4808 VPWR _0144_ 0.28784f
C4809 _0464_ _0472_ 0
C4810 _0625_/a_59_75# acc0.A\[6\] 0
C4811 _0553_/a_512_297# comp0.B\[6\] 0.00281f
C4812 clknet_0__0458_ net248 0
C4813 _0817_/a_266_297# acc0.A\[9\] 0.00114f
C4814 _0549_/a_68_297# net171 0.17745f
C4815 _0437_ _0989_/a_592_47# 0
C4816 acc0.A\[24\] _1006_/a_1059_315# 0
C4817 _0284_ _0399_ 0
C4818 _0190_ _0988_/a_27_47# 0
C4819 clknet_0__0459_ net103 0
C4820 net245 pp[14] 0.02479f
C4821 acc0.A\[10\] hold70/a_285_47# 0.00364f
C4822 _0343_ net66 0
C4823 _0118_ _0346_ 0
C4824 clkload1/a_110_47# clknet_1_1__leaf__0458_ 0
C4825 clkbuf_1_0__f__0459_/a_110_47# _1016_/a_193_47# 0.00236f
C4826 _1020_/a_1059_315# acc0.A\[20\] 0.0943f
C4827 _0217_ _1014_/a_27_47# 0.07748f
C4828 _0295_ _0420_ 0
C4829 net25 _0175_ 0.02228f
C4830 net202 _0181_ 0.03536f
C4831 _0243_ _0099_ 0
C4832 _1042_/a_27_47# net19 0
C4833 _1042_/a_466_413# _0203_ 0
C4834 _1012_/a_1017_47# _0352_ 0
C4835 _0239_ _0240_ 0.10963f
C4836 _0369_ _0184_ 0
C4837 net36 _0953_/a_32_297# 0
C4838 _0555_/a_149_47# _0175_ 0
C4839 clknet_1_1__leaf__0463_ _0181_ 0
C4840 _0239_ _0369_ 0
C4841 clknet_1_0__leaf__0458_ _0179_ 0.45999f
C4842 hold58/a_49_47# _0554_/a_68_297# 0
C4843 clknet_0_clk net17 0.02163f
C4844 _0131_ _0564_/a_68_297# 0
C4845 _0786_/a_472_297# _0345_ 0
C4846 _0780_/a_285_297# _0392_ 0
C4847 _0984_/a_1059_315# acc0.A\[15\] 0.00759f
C4848 clknet_1_0__leaf__0459_ _1017_/a_561_413# 0
C4849 _0343_ _0991_/a_27_47# 0.02578f
C4850 hold87/a_391_47# net165 0
C4851 _0120_ _0222_ 0.03153f
C4852 VPWR _1028_/a_634_159# 0.18021f
C4853 _1069_/a_634_159# _1069_/a_1059_315# 0
C4854 _1069_/a_27_47# _1069_/a_381_47# 0.06222f
C4855 _1069_/a_193_47# _1069_/a_891_413# 0.19286f
C4856 hold4/a_49_47# net109 0.01001f
C4857 _0230_ net46 0.01986f
C4858 net167 _0170_ 0.01669f
C4859 _0343_ _0773_/a_285_297# 0.00989f
C4860 _0151_ VPWR 0.87797f
C4861 _0275_ _0089_ 0
C4862 net128 net20 0.00158f
C4863 _1059_/a_466_413# _0507_/a_109_297# 0
C4864 output43/a_27_47# hold78/a_285_47# 0
C4865 net106 net118 0.1233f
C4866 _0714_/a_240_47# _0587_/a_27_47# 0
C4867 _1037_/a_634_159# comp0.B\[4\] 0
C4868 _1041_/a_27_47# _1040_/a_27_47# 0.01278f
C4869 _1031_/a_27_47# _0220_ 0.05572f
C4870 _0955_/a_32_297# _0160_ 0
C4871 _0536_/a_245_297# _0172_ 0
C4872 net69 _0446_ 0
C4873 _0136_ net29 0.05137f
C4874 _0253_ _0827_/a_27_47# 0.00112f
C4875 net8 _0181_ 0
C4876 output48/a_27_47# net49 0.00747f
C4877 net48 output49/a_27_47# 0.00313f
C4878 net58 _1055_/a_193_47# 0
C4879 _1059_/a_193_47# hold82/a_391_47# 0
C4880 _1059_/a_634_159# hold82/a_285_47# 0.00139f
C4881 output66/a_27_47# _0515_/a_299_297# 0
C4882 clknet_1_1__leaf__0460_ _0387_ 0.00244f
C4883 hold37/a_391_47# VPWR 0.18033f
C4884 _0400_ net5 0
C4885 _1030_/a_27_47# net209 0.09822f
C4886 _0985_/a_381_47# _0350_ 0
C4887 net50 net51 0.00201f
C4888 net7 _0159_ 0.02768f
C4889 _0486_ _0468_ 0.24486f
C4890 net22 _0139_ 0.07716f
C4891 _0733_/a_79_199# acc0.A\[25\] 0.00127f
C4892 hold87/a_391_47# acc0.A\[19\] 0
C4893 hold87/a_49_47# _0242_ 0
C4894 _0176_ _0544_/a_51_297# 0
C4895 _0718_/a_47_47# pp[28] 0.03706f
C4896 _1002_/a_27_47# _0181_ 0.02205f
C4897 hold89/a_285_47# _0961_/a_113_297# 0
C4898 comp0.B\[2\] comp0.B\[1\] 0.14223f
C4899 _0257_ _0434_ 0
C4900 net239 _0219_ 0
C4901 _0183_ net91 0.00162f
C4902 acc0.A\[22\] _0103_ 0
C4903 clknet_0__0463_ clkbuf_1_0__f__0463_/a_110_47# 0.31962f
C4904 _0607_/a_109_47# _0181_ 0
C4905 net190 acc0.A\[28\] 0.5698f
C4906 _0538_/a_51_297# _0538_/a_240_47# 0.03076f
C4907 _0343_ _0350_ 0.37623f
C4908 hold75/a_49_47# _0848_/a_27_47# 0
C4909 _1037_/a_891_413# net26 0.00186f
C4910 clknet_1_1__leaf__0462_ _1008_/a_975_413# 0
C4911 _0715_/a_27_47# _0428_ 0
C4912 _0474_ _0561_/a_149_47# 0.00276f
C4913 comp0.B\[3\] _0173_ 0
C4914 _0216_ _0366_ 0
C4915 hold43/a_49_47# clknet_1_1__leaf__0462_ 0
C4916 hold47/a_391_47# _0172_ 0
C4917 _0343_ _0111_ 0.05672f
C4918 _0183_ hold18/a_49_47# 0.03081f
C4919 _1022_/a_634_159# _1022_/a_1017_47# 0
C4920 _1022_/a_466_413# _1022_/a_592_47# 0.00553f
C4921 _1065_/a_27_47# _1062_/a_193_47# 0
C4922 net47 _0345_ 0.31771f
C4923 net87 net223 0
C4924 _0677_/a_47_47# clknet_0__0461_ 0
C4925 _0994_/a_634_159# _0994_/a_466_413# 0.23992f
C4926 _0994_/a_193_47# _0994_/a_1059_315# 0.03405f
C4927 _0994_/a_27_47# _0994_/a_891_413# 0.03224f
C4928 clknet_1_0__leaf__0463_ _0139_ 0
C4929 _0153_ _0189_ 0
C4930 acc0.A\[26\] _0737_/a_35_297# 0
C4931 _1020_/a_193_47# clknet_1_0__leaf__0457_ 0.04019f
C4932 _0275_ _0986_/a_891_413# 0.04718f
C4933 _0284_ _0808_/a_266_297# 0
C4934 _0285_ _0808_/a_368_297# 0.00571f
C4935 net211 _1001_/a_381_47# 0.01148f
C4936 _0475_ comp0.B\[6\] 0.03852f
C4937 net62 _0840_/a_68_297# 0.12262f
C4938 _0179_ _0525_/a_299_297# 0.0529f
C4939 pp[7] pp[5] 0.19978f
C4940 _1055_/a_634_159# net179 0.02916f
C4941 _1055_/a_466_413# net141 0
C4942 _1023_/a_193_47# output51/a_27_47# 0
C4943 VPWR hold3/a_49_47# 0.31281f
C4944 _0718_/a_377_297# _0216_ 0
C4945 _0422_ hold81/a_49_47# 0
C4946 hold5/a_285_47# _1043_/a_1059_315# 0
C4947 net53 acc0.A\[25\] 0.66536f
C4948 _0399_ _0267_ 0.02266f
C4949 _0995_/a_193_47# _0218_ 0.00643f
C4950 _0984_/a_1059_315# _0179_ 0
C4951 _1003_/a_1059_315# _1003_/a_1017_47# 0
C4952 _1003_/a_193_47# net89 0.00679f
C4953 _1003_/a_27_47# _0101_ 0.09837f
C4954 _0343_ _0621_/a_35_297# 0.02771f
C4955 net36 _1047_/a_634_159# 0.03777f
C4956 _1036_/a_466_413# net27 0
C4957 _0984_/a_27_47# _0181_ 0.00441f
C4958 _0693_/a_150_297# _0324_ 0.00105f
C4959 net171 _1040_/a_891_413# 0
C4960 _0217_ _0195_ 0.09516f
C4961 hold26/a_285_47# comp0.B\[10\] 0
C4962 hold2/a_49_47# net47 0
C4963 _0967_/a_297_297# VPWR 0.00866f
C4964 VPWR _0162_ 0.92254f
C4965 hold33/a_285_47# _0548_/a_240_47# 0
C4966 net185 comp0.B\[5\] 0.12869f
C4967 _0176_ _0141_ 0.07244f
C4968 hold46/a_285_47# _0172_ 0
C4969 VPWR _0371_ 0.59008f
C4970 _0211_ B[5] 0
C4971 _0183_ _0856_/a_297_297# 0.00166f
C4972 clkload0/X clknet_1_0__leaf_clk 0.02668f
C4973 _0257_ _0989_/a_1059_315# 0
C4974 _0844_/a_297_47# _0447_ 0.00798f
C4975 _1004_/a_561_413# _0352_ 0
C4976 _1004_/a_381_47# _0102_ 0.13116f
C4977 _0456_ net206 0
C4978 net33 _1062_/a_27_47# 0.00459f
C4979 _0733_/a_222_93# _0737_/a_35_297# 0
C4980 _0534_/a_81_21# net175 0
C4981 hold56/a_391_47# comp0.B\[2\] 0.00482f
C4982 net162 _0704_/a_68_297# 0.00107f
C4983 hold15/a_285_47# acc0.A\[30\] 0
C4984 net23 _1065_/a_891_413# 0.0274f
C4985 hold91/a_285_47# acc0.A\[15\] 0
C4986 hold18/a_49_47# acc0.A\[15\] 0.30157f
C4987 clknet_1_1__leaf__0459_ _0405_ 0.00641f
C4988 net140 _1053_/a_27_47# 0.03595f
C4989 net229 net6 0
C4990 _0626_/a_150_297# _0465_ 0
C4991 _0080_ _0456_ 0
C4992 clkbuf_1_0__f_clk/a_110_47# _0484_ 0
C4993 _0793_/a_51_297# net41 0.00562f
C4994 _0992_/a_27_47# _0809_/a_81_21# 0
C4995 VPWR _0987_/a_975_413# 0.00523f
C4996 clkbuf_1_0__f__0459_/a_110_47# net41 0
C4997 _0183_ _0247_ 0.07888f
C4998 hold30/a_285_47# _0225_ 0.01818f
C4999 _1024_/a_193_47# _1024_/a_381_47# 0.0982f
C5000 _1024_/a_634_159# _1024_/a_891_413# 0.03684f
C5001 _1024_/a_27_47# _1024_/a_561_413# 0.0027f
C5002 hold23/a_391_47# net175 0
C5003 net86 hold72/a_49_47# 0
C5004 net150 _0369_ 0.45955f
C5005 _0458_ VPWR 0.9108f
C5006 _0816_/a_68_297# _0425_ 0
C5007 net48 hold3/a_49_47# 0.02519f
C5008 _0349_ _0707_/a_75_199# 0
C5009 hold41/a_391_47# net67 0.02466f
C5010 clkbuf_1_0__f__0457_/a_110_47# _0183_ 0.00104f
C5011 hold56/a_49_47# clkbuf_1_1__f_clk/a_110_47# 0
C5012 _1011_/a_466_413# _0333_ 0
C5013 _0797_/a_27_413# net6 0
C5014 _0985_/a_634_159# _0180_ 0
C5015 net33 _0561_/a_51_297# 0
C5016 _1000_/a_975_413# _0244_ 0
C5017 VPWR _1029_/a_975_413# 0.00515f
C5018 net61 _0829_/a_109_297# 0
C5019 net46 _0236_ 0
C5020 comp0.B\[2\] _1032_/a_634_159# 0
C5021 clk _1064_/a_634_159# 0.00448f
C5022 hold96/a_49_47# _0217_ 0.05073f
C5023 _1048_/a_634_159# _1048_/a_592_47# 0
C5024 _0712_/a_79_21# _0220_ 0.01953f
C5025 _1034_/a_891_413# clknet_1_1__leaf__0463_ 0.01594f
C5026 net165 _0264_ 0.12327f
C5027 acc0.A\[14\] _0794_/a_27_47# 0
C5028 hold34/a_49_47# acc0.A\[9\] 0.30062f
C5029 _0831_/a_35_297# _0826_/a_27_53# 0
C5030 _0225_ _0102_ 0
C5031 clknet_0__0461_ _0242_ 0.3312f
C5032 net235 pp[4] 0
C5033 VPWR _1016_/a_466_413# 0.23576f
C5034 acc0.A\[16\] _0780_/a_35_297# 0
C5035 _1035_/a_27_47# net24 0
C5036 _0846_/a_149_47# _0448_ 0.0215f
C5037 net173 _0138_ 0
C5038 _0512_/a_27_297# clknet_1_1__leaf__0465_ 0
C5039 _0433_ _0824_/a_59_75# 0
C5040 _0376_ _0350_ 0
C5041 _0429_ _0434_ 0.00601f
C5042 _0856_/a_297_297# acc0.A\[15\] 0
C5043 net204 VPWR 0.29691f
C5044 _0254_ _0826_/a_219_297# 0
C5045 _0460_ net241 0
C5046 _0133_ net33 0
C5047 net68 net157 0
C5048 hold11/a_285_47# net158 0.01139f
C5049 _0305_ clkbuf_0__0460_/a_110_47# 0
C5050 net172 _0206_ 0
C5051 _1016_/a_193_47# clkbuf_0__0461_/a_110_47# 0
C5052 _1060_/a_27_47# _0219_ 0
C5053 _0670_/a_215_47# acc0.A\[15\] 0.05952f
C5054 _0096_ _0218_ 0.05513f
C5055 hold23/a_49_47# acc0.A\[3\] 0.30589f
C5056 _0217_ _0081_ 0
C5057 _0183_ _0455_ 0
C5058 _0264_ acc0.A\[19\] 0
C5059 hold27/a_49_47# VPWR 0.29749f
C5060 hold33/a_285_47# net7 0.03968f
C5061 _0569_/a_27_297# _1028_/a_1059_315# 0
C5062 _0273_ acc0.A\[6\] 0.22627f
C5063 net78 clknet_1_1__leaf__0459_ 0.17284f
C5064 net32 _0544_/a_240_47# 0.00544f
C5065 _0205_ _0204_ 0
C5066 _0546_/a_240_47# net18 0
C5067 _0192_ net140 0
C5068 _0357_ _0219_ 0.01295f
C5069 net45 _0408_ 0.00118f
C5070 _0948_/a_109_297# _0471_ 0.0039f
C5071 _0349_ _0351_ 0.08977f
C5072 comp0.B\[1\] _1015_/a_193_47# 0
C5073 _1010_/a_381_47# net96 0
C5074 _0179_ hold18/a_49_47# 0
C5075 _1032_/a_193_47# _0584_/a_27_297# 0
C5076 _1056_/a_27_47# _0189_ 0.0028f
C5077 hold6/a_49_47# net152 0.01635f
C5078 comp0.B\[15\] _0171_ 0.14832f
C5079 _0130_ _1015_/a_381_47# 0
C5080 _1040_/a_634_159# net174 0.02969f
C5081 _0216_ _0689_/a_68_297# 0
C5082 _0797_/a_207_413# _0797_/a_297_47# 0.00476f
C5083 _1053_/a_193_47# acc0.A\[6\] 0
C5084 clknet_1_0__leaf__0465_ _1054_/a_634_159# 0
C5085 hold28/a_391_47# net71 0
C5086 _0748_/a_299_297# _0312_ 0
C5087 _0357_ _0728_/a_59_75# 0.1131f
C5088 _0979_/a_27_297# _0169_ 0.10893f
C5089 _0979_/a_373_47# net164 0.0019f
C5090 _0617_/a_68_297# _0373_ 0
C5091 _1031_/a_193_47# _0218_ 0
C5092 net232 comp0.B\[3\] 0
C5093 _1072_/a_193_47# _1072_/a_381_47# 0.10164f
C5094 _1072_/a_634_159# _1072_/a_891_413# 0.03684f
C5095 _1072_/a_27_47# _1072_/a_561_413# 0.00163f
C5096 _0830_/a_215_47# _0186_ 0
C5097 _0216_ _1027_/a_1017_47# 0.00125f
C5098 _0841_/a_215_47# _0841_/a_510_47# 0.00529f
C5099 net168 _0437_ 0.00455f
C5100 _0278_ _0414_ 0
C5101 _0183_ _0505_/a_109_297# 0.01134f
C5102 _0172_ net127 0.00292f
C5103 net30 net153 0
C5104 clkbuf_1_0__f__0458_/a_110_47# _0448_ 0
C5105 _0714_/a_240_47# VPWR 0.00139f
C5106 _0313_ _0732_/a_209_47# 0.00132f
C5107 _0248_ net92 0.0319f
C5108 _1020_/a_27_47# _0586_/a_27_47# 0
C5109 net237 hold90/a_49_47# 0
C5110 hold68/a_285_47# _0758_/a_79_21# 0
C5111 _0221_ hold80/a_49_47# 0
C5112 net45 net166 0.00154f
C5113 acc0.A\[7\] net11 0
C5114 net9 net73 0
C5115 control0.count\[2\] _0484_ 0
C5116 _0136_ _0137_ 0.0019f
C5117 net44 hold95/a_391_47# 0
C5118 _0251_ _0252_ 0.35992f
C5119 _0429_ acc0.A\[7\] 0.10818f
C5120 _0244_ _1018_/a_891_413# 0
C5121 clknet_1_0__leaf__0460_ clknet_1_0__leaf__0461_ 0.16169f
C5122 _1001_/a_592_47# _0345_ 0.00135f
C5123 _0369_ control0.add 0.11077f
C5124 comp0.B\[4\] _0561_/a_512_297# 0
C5125 _0429_ _0989_/a_1059_315# 0
C5126 _0251_ _0989_/a_381_47# 0.00261f
C5127 _0413_ _0410_ 0
C5128 clknet_0__0457_ control0.add 0.00934f
C5129 _0608_/a_109_297# _0097_ 0
C5130 _0179_ _0288_ 0.0091f
C5131 _0713_/a_27_47# _1019_/a_27_47# 0.00192f
C5132 _1003_/a_27_47# net35 0.00774f
C5133 _0462_ _0246_ 0.00453f
C5134 _0819_/a_81_21# net47 0.00497f
C5135 _0217_ net90 0
C5136 clknet_1_1__leaf__0460_ _1006_/a_27_47# 0
C5137 _0985_/a_193_47# net10 0
C5138 _0343_ _0244_ 0.04502f
C5139 clknet_0_clk _0165_ 0
C5140 _1004_/a_634_159# _0380_ 0
C5141 _0252_ _0989_/a_592_47# 0
C5142 _0989_/a_891_413# _0989_/a_1017_47# 0.00617f
C5143 _0997_/a_193_47# _0997_/a_381_47# 0.09503f
C5144 _0997_/a_634_159# _0997_/a_891_413# 0.03684f
C5145 _0997_/a_27_47# _0997_/a_561_413# 0.00163f
C5146 _0314_ clknet_0__0460_ 0
C5147 hold56/a_49_47# VPWR 0.32936f
C5148 _0455_ acc0.A\[15\] 0
C5149 _0544_/a_149_47# _1042_/a_891_413# 0
C5150 _0544_/a_240_47# _1042_/a_1059_315# 0
C5151 _0093_ _0218_ 0.02706f
C5152 net78 _0292_ 0
C5153 _0181_ _0986_/a_561_413# 0
C5154 _0348_ _0335_ 0.03367f
C5155 _0121_ net46 0.038f
C5156 net162 _0216_ 0.17928f
C5157 _0292_ clknet_0__0465_ 0.0595f
C5158 acc0.A\[27\] _0319_ 0
C5159 _0439_ clkbuf_1_1__f__0458_/a_110_47# 0.00241f
C5160 _0476_ control0.sh 0.09175f
C5161 _0992_/a_891_413# _0992_/a_1017_47# 0.00617f
C5162 VPWR _1051_/a_891_413# 0.19541f
C5163 _0569_/a_27_297# _0347_ 0
C5164 _0327_ clkbuf_1_0__f__0462_/a_110_47# 0
C5165 _0255_ net62 0
C5166 VPWR clkbuf_1_1__f__0458_/a_110_47# 1.35349f
C5167 _0309_ _0240_ 0.08066f
C5168 hold6/a_285_47# _1042_/a_634_159# 0
C5169 VPWR _1045_/a_561_413# 0.00296f
C5170 _0465_ control0.reset 0.00533f
C5171 _0309_ _0369_ 0
C5172 _1052_/a_1059_315# _0369_ 0
C5173 _0355_ _1029_/a_1017_47# 0
C5174 _0109_ _1029_/a_381_47# 0
C5175 hold13/a_391_47# _0474_ 0.00146f
C5176 hold63/a_285_47# VPWR 0.29303f
C5177 net230 acc0.A\[6\] 0
C5178 clknet_1_1__leaf__0464_ _0194_ 0.00291f
C5179 _1045_/a_193_47# net129 0
C5180 _0407_ _0792_/a_80_21# 0.05315f
C5181 net86 clknet_0__0461_ 0.02393f
C5182 _1027_/a_27_47# _1027_/a_1059_315# 0.04875f
C5183 _1027_/a_193_47# _1027_/a_466_413# 0.07855f
C5184 _0743_/a_512_297# _0105_ 0
C5185 net58 _0252_ 0
C5186 _1055_/a_27_47# net47 0.00209f
C5187 _0253_ _0830_/a_510_47# 0
C5188 hold46/a_391_47# hold26/a_391_47# 0
C5189 acc0.A\[15\] _0505_/a_109_297# 0.00366f
C5190 hold59/a_285_47# net149 0
C5191 _0996_/a_193_47# net41 0.00691f
C5192 _0465_ _1061_/a_891_413# 0.00701f
C5193 VPWR _1032_/a_27_47# 0.64116f
C5194 _1061_/a_634_159# _1061_/a_592_47# 0
C5195 _0753_/a_79_21# _0222_ 0.03453f
C5196 A[13] _0277_ 0
C5197 _0305_ _1009_/a_27_47# 0.00122f
C5198 _0955_/a_114_297# net25 0
C5199 _0368_ _0360_ 0.29478f
C5200 acc0.A\[8\] _0990_/a_891_413# 0
C5201 _0291_ _0990_/a_1059_315# 0
C5202 net66 _0990_/a_381_47# 0
C5203 net160 net28 0
C5204 net203 _0171_ 0
C5205 _0143_ _0527_/a_27_297# 0
C5206 clkbuf_1_0__f__0457_/a_110_47# hold40/a_285_47# 0.02f
C5207 hold101/a_49_47# _0440_ 0.0017f
C5208 _0216_ net112 0.10464f
C5209 _1007_/a_592_47# _0219_ 0
C5210 _0136_ comp0.B\[6\] 0.11043f
C5211 net126 _1038_/a_381_47# 0
C5212 _0266_ _0347_ 0
C5213 _0107_ _0362_ 0
C5214 _0319_ _0364_ 0.06856f
C5215 clkbuf_0__0459_/a_110_47# net5 0.00164f
C5216 _0216_ acc0.A\[24\] 0.02302f
C5217 _1035_/a_634_159# _1035_/a_1059_315# 0
C5218 _1035_/a_27_47# _1035_/a_381_47# 0.06222f
C5219 _1035_/a_193_47# _1035_/a_891_413# 0.19489f
C5220 net207 _0526_/a_27_47# 0
C5221 _0734_/a_285_47# _0219_ 0.01028f
C5222 _0483_ _0482_ 0.10484f
C5223 _0279_ _0277_ 0.01551f
C5224 VPWR pp[14] 0.44923f
C5225 _0278_ _0300_ 0
C5226 clknet_1_1__leaf__0458_ _0434_ 0.06442f
C5227 _0697_/a_80_21# _0690_/a_68_297# 0.00113f
C5228 _1053_/a_27_47# input14/a_75_212# 0
C5229 clknet_1_0__leaf__0462_ hold68/a_285_47# 0.01225f
C5230 net36 _0174_ 0.03359f
C5231 net56 _0690_/a_68_297# 0
C5232 _0489_ _1069_/a_381_47# 0.00133f
C5233 _0218_ _0395_ 0.06429f
C5234 _0661_/a_205_297# _0425_ 0
C5235 _0289_ _0815_/a_113_297# 0
C5236 _0217_ _0573_/a_27_47# 0.33689f
C5237 input33/a_75_212# B[4] 0.00215f
C5238 _1013_/a_634_159# clknet_1_1__leaf__0461_ 0
C5239 VPWR _0767_/a_59_75# 0.2365f
C5240 net140 A[5] 0.01531f
C5241 _1010_/a_27_47# _0701_/a_80_21# 0
C5242 hold11/a_391_47# net134 0
C5243 _1054_/a_27_47# acc0.A\[8\] 0
C5244 hold20/a_391_47# _0466_ 0
C5245 acc0.A\[15\] _0506_/a_299_297# 0.00308f
C5246 acc0.A\[29\] _1029_/a_634_159# 0.00273f
C5247 _0294_ _0345_ 0.11584f
C5248 _0294_ _0814_/a_27_47# 0.00205f
C5249 clknet_1_0__leaf__0459_ _1016_/a_466_413# 0
C5250 _0399_ _0178_ 0
C5251 _1069_/a_466_413# _0167_ 0.00559f
C5252 _1069_/a_1059_315# clknet_1_0__leaf_clk 0
C5253 _1069_/a_27_47# control0.count\[0\] 0.01326f
C5254 VPWR net114 0.37926f
C5255 net44 net209 0.06143f
C5256 hold88/a_285_47# acc0.A\[6\] 0
C5257 _0384_ hold73/a_391_47# 0
C5258 hold74/a_49_47# _0781_/a_150_297# 0
C5259 _1059_/a_592_47# acc0.A\[13\] 0
C5260 pp[8] _1055_/a_1059_315# 0
C5261 _0233_ _0600_/a_253_47# 0.00268f
C5262 _0181_ _0498_/a_245_297# 0
C5263 _0474_ _0160_ 0
C5264 net213 _0383_ 0.09043f
C5265 hold10/a_285_47# net125 0
C5266 net145 hold82/a_285_47# 0
C5267 _0157_ hold82/a_49_47# 0
C5268 _0525_/a_81_21# hold83/a_285_47# 0
C5269 _0482_ control0.count\[1\] 0.0115f
C5270 _0488_ _0970_/a_114_47# 0
C5271 _0953_/a_32_297# _1061_/a_27_47# 0.00121f
C5272 hold19/a_391_47# _0219_ 0
C5273 _0846_/a_245_297# acc0.A\[15\] 0
C5274 _0243_ _0238_ 0
C5275 _1001_/a_27_47# _0346_ 0.01123f
C5276 net104 clkbuf_1_0__f__0461_/a_110_47# 0
C5277 _0415_ _0399_ 0.00967f
C5278 _0461_ _0869_/a_27_47# 0.0088f
C5279 _0568_/a_27_297# hold62/a_285_47# 0.00104f
C5280 _0959_/a_300_47# net33 0
C5281 net167 net35 0.00507f
C5282 net87 clkbuf_0__0457_/a_110_47# 0
C5283 _0311_ _0679_/a_68_297# 0.10805f
C5284 _0183_ _1022_/a_891_413# 0
C5285 acc0.A\[22\] _1022_/a_381_47# 0
C5286 _0120_ _1022_/a_466_413# 0
C5287 _0577_/a_27_297# net151 0.00905f
C5288 comp0.B\[2\] _0496_/a_27_47# 0.0073f
C5289 acc0.A\[7\] clknet_1_1__leaf__0458_ 0.05504f
C5290 clknet_1_1__leaf__0458_ _0989_/a_1059_315# 0
C5291 clknet_0__0457_ clknet_1_1__leaf__0457_ 0.00758f
C5292 _0538_/a_512_297# _0143_ 0
C5293 _0233_ _0751_/a_29_53# 0
C5294 _0086_ acc0.A\[6\] 0.00314f
C5295 VPWR _0760_/a_129_47# 0
C5296 clknet_1_0__leaf__0463_ _0498_/a_240_47# 0.00228f
C5297 _0411_ _0668_/a_79_21# 0
C5298 _0524_/a_27_297# net148 0.10471f
C5299 hold20/a_391_47# net236 0
C5300 net53 net210 0.03943f
C5301 _0343_ _0986_/a_634_159# 0
C5302 clknet_1_0__leaf__0459_ _1019_/a_592_47# 0
C5303 _0298_ A[13] 0
C5304 hold64/a_391_47# _0580_/a_109_297# 0
C5305 _0579_/a_109_297# _1019_/a_27_47# 0
C5306 net45 net117 0
C5307 _0575_/a_27_297# acc0.A\[25\] 0
C5308 net36 _0208_ 0
C5309 _0550_/a_51_297# B[7] 0.00143f
C5310 _0259_ _0427_ 0.58664f
C5311 _0284_ _0091_ 0.2366f
C5312 net141 net179 0.01115f
C5313 VPWR _0365_ 0.76167f
C5314 _0972_/a_93_21# _0972_/a_584_47# 0.00278f
C5315 clkbuf_0__0463_/a_110_47# control0.sh 0.01043f
C5316 _0290_ _0990_/a_1059_315# 0
C5317 _0401_ _0990_/a_466_413# 0
C5318 _0966_/a_27_47# _0484_ 0.10131f
C5319 _0416_ _0277_ 0.00238f
C5320 _0752_/a_384_47# _0222_ 0.01016f
C5321 _0179_ _0506_/a_299_297# 0.10916f
C5322 hold37/a_285_47# _0172_ 0
C5323 net161 net27 0
C5324 comp0.B\[11\] net20 0.11621f
C5325 _0279_ _0298_ 0.10455f
C5326 _0278_ _0404_ 0
C5327 _0993_/a_193_47# _0993_/a_381_47# 0.10164f
C5328 _0993_/a_634_159# _0993_/a_891_413# 0.03684f
C5329 _0993_/a_27_47# _0993_/a_561_413# 0.0027f
C5330 _1058_/a_381_47# net192 0
C5331 _1058_/a_1059_315# _0156_ 0
C5332 clkload1/a_110_47# _0218_ 0
C5333 _0180_ net201 0
C5334 hold48/a_49_47# comp0.B\[12\] 0.33522f
C5335 net63 _0399_ 0.00139f
C5336 hold45/a_391_47# net144 0.05937f
C5337 _1039_/a_634_159# _1039_/a_592_47# 0
C5338 net185 hold84/a_49_47# 0
C5339 _0182_ _0531_/a_109_47# 0.00324f
C5340 _0180_ _0531_/a_109_297# 0.01807f
C5341 hold67/a_285_47# _0369_ 0.04285f
C5342 net46 _0380_ 0.01029f
C5343 _0785_/a_299_297# clknet_0__0465_ 0.03492f
C5344 hold32/a_285_47# acc0.A\[9\] 0.00157f
C5345 net175 hold71/a_391_47# 0
C5346 _1039_/a_27_47# _0953_/a_32_297# 0
C5347 _1038_/a_27_47# _0463_ 0
C5348 _0551_/a_27_47# _0175_ 0
C5349 _0483_ hold89/a_285_47# 0.00135f
C5350 _0663_/a_207_413# _0289_ 0.00567f
C5351 _0663_/a_27_413# _0287_ 0.03203f
C5352 _0346_ _0420_ 0.12082f
C5353 _0736_/a_311_297# _0371_ 0
C5354 _0172_ _1046_/a_975_413# 0
C5355 hold52/a_49_47# _0105_ 0
C5356 clknet_0__0462_ _0686_/a_219_297# 0.03971f
C5357 net55 net224 0.24023f
C5358 _0222_ clkbuf_1_0__f__0460_/a_110_47# 0.01163f
C5359 net26 net27 0.23494f
C5360 _0402_ _0511_/a_81_21# 0
C5361 _1026_/a_193_47# _1026_/a_592_47# 0.00135f
C5362 _1026_/a_466_413# _1026_/a_561_413# 0.00772f
C5363 _1026_/a_634_159# _1026_/a_975_413# 0
C5364 hold74/a_391_47# _0369_ 0.00148f
C5365 clknet_0__0462_ _1008_/a_1059_315# 0
C5366 _0991_/a_27_47# _0842_/a_59_75# 0
C5367 _0346_ _0459_ 0
C5368 _0330_ net97 0
C5369 acc0.A\[4\] acc0.A\[6\] 0
C5370 _0222_ _0250_ 0.00257f
C5371 _0629_/a_145_75# _0263_ 0.00281f
C5372 pp[9] net181 0.02174f
C5373 net17 _1065_/a_27_47# 0
C5374 _0181_ _1009_/a_27_47# 0.04875f
C5375 _0695_/a_80_21# _0359_ 0.01376f
C5376 VPWR _0408_ 0.36204f
C5377 _1024_/a_891_413# net110 0
C5378 _1024_/a_1059_315# _0122_ 0
C5379 _1024_/a_193_47# acc0.A\[24\] 0
C5380 acc0.A\[21\] _0228_ 0.11261f
C5381 clkbuf_0_clk/a_110_47# _0471_ 0.02646f
C5382 _0349_ _0338_ 0
C5383 B[9] net128 0.01762f
C5384 _1014_/a_891_413# _0181_ 0
C5385 _0278_ _0646_/a_285_47# 0.05006f
C5386 clknet_1_1__leaf__0464_ net195 0
C5387 _0715_/a_27_47# net72 0
C5388 _0375_ _0223_ 0.00873f
C5389 _0083_ _0182_ 0.01165f
C5390 net93 net52 0.20054f
C5391 net61 _0827_/a_27_47# 0.00136f
C5392 hold99/a_49_47# output38/a_27_47# 0.02626f
C5393 _1057_/a_466_413# net143 0
C5394 pp[16] _0997_/a_634_159# 0
C5395 net45 _0388_ 0
C5396 hold89/a_285_47# control0.count\[1\] 0
C5397 hold21/a_285_47# _1054_/a_1059_315# 0
C5398 VPWR _0291_ 0.43499f
C5399 _0180_ _1049_/a_1017_47# 0
C5400 _0202_ net20 0.0252f
C5401 _0949_/a_59_75# _0166_ 0
C5402 net168 _0252_ 0.01058f
C5403 _0186_ _0989_/a_27_47# 0
C5404 hold1/a_49_47# _0186_ 0
C5405 _0470_ net26 0.00148f
C5406 _0957_/a_114_297# net24 0.00396f
C5407 _0195_ _0999_/a_1059_315# 0
C5408 _0533_/a_109_297# control0.sh 0
C5409 _0350_ _0842_/a_59_75# 0
C5410 _0562_/a_68_297# _0493_/a_27_47# 0.0013f
C5411 _0790_/a_35_297# _0790_/a_117_297# 0.00641f
C5412 VPWR net166 0.33889f
C5413 _1068_/a_975_413# _0468_ 0
C5414 net120 hold39/a_285_47# 0
C5415 _0538_/a_51_297# _0473_ 0.10608f
C5416 _1041_/a_634_159# _1041_/a_1059_315# 0
C5417 _1041_/a_27_47# _1041_/a_381_47# 0.05761f
C5418 _1041_/a_193_47# _1041_/a_891_413# 0.19207f
C5419 _0343_ _1013_/a_975_413# 0
C5420 VPWR _0991_/a_634_159# 0.19008f
C5421 clknet_1_0__leaf__0460_ _0105_ 0
C5422 _0362_ _0322_ 0
C5423 _1059_/a_1059_315# _0289_ 0
C5424 net22 _0954_/a_32_297# 0
C5425 _0294_ net52 0
C5426 _0362_ _0327_ 0
C5427 _0603_/a_68_297# _0383_ 0
C5428 _0176_ _1043_/a_27_47# 0.01235f
C5429 hold76/a_285_47# _1001_/a_1059_315# 0.0054f
C5430 input12/a_75_212# A[7] 0.0031f
C5431 A[5] input14/a_75_212# 0.00249f
C5432 net31 hold6/a_285_47# 0
C5433 _0346_ _0265_ 0.01824f
C5434 hold54/a_285_47# VPWR 0.27409f
C5435 acc0.A\[12\] _0650_/a_68_297# 0.0109f
C5436 _0569_/a_109_47# net114 0
C5437 _0490_ net159 0
C5438 acc0.A\[29\] _0723_/a_27_413# 0.0517f
C5439 _1051_/a_466_413# acc0.A\[6\] 0
C5440 hold86/a_285_47# _0345_ 0.01294f
C5441 _0416_ _0296_ 0
C5442 _0616_/a_215_47# _0242_ 0
C5443 hold12/a_285_47# net17 0
C5444 _0399_ _0812_/a_79_21# 0.10311f
C5445 net44 clknet_0__0461_ 0.0123f
C5446 _0369_ _0610_/a_145_75# 0.00331f
C5447 clknet_1_0__leaf__0465_ net140 0.10016f
C5448 _1057_/a_381_47# _0512_/a_27_297# 0
C5449 hold44/a_391_47# _1029_/a_466_413# 0
C5450 hold44/a_49_47# _1029_/a_891_413# 0
C5451 pp[6] pp[4] 0.18239f
C5452 _0195_ _0530_/a_81_21# 0.08008f
C5453 hold54/a_49_47# _1015_/a_1059_315# 0.00266f
C5454 _0476_ _0955_/a_32_297# 0.0279f
C5455 _0343_ _0984_/a_381_47# 0.00654f
C5456 _0794_/a_326_47# net41 0
C5457 net81 net43 0
C5458 _0176_ _0171_ 0
C5459 _0782_/a_27_47# hold60/a_285_47# 0.00123f
C5460 hold38/a_49_47# net186 0.00836f
C5461 clkbuf_1_1__f_clk/a_110_47# _0950_/a_75_212# 0
C5462 _0081_ _0583_/a_373_47# 0
C5463 _0454_ net165 0
C5464 _0135_ _0549_/a_68_297# 0
C5465 _1013_/a_561_413# net60 0
C5466 _0661_/a_27_297# net67 0.0082f
C5467 _0661_/a_277_297# _0089_ 0
C5468 net31 _1041_/a_1017_47# 0.00171f
C5469 _0467_ hold39/a_391_47# 0
C5470 _0258_ net72 0
C5471 comp0.B\[4\] _0132_ 0.016f
C5472 _0432_ _0433_ 0.02931f
C5473 _0624_/a_59_75# acc0.A\[4\] 0.08318f
C5474 _0743_/a_512_297# _0359_ 0.00325f
C5475 _0182_ _0584_/a_27_297# 0
C5476 _1012_/a_193_47# _0351_ 0.00205f
C5477 _1063_/a_1059_315# hold93/a_49_47# 0.00135f
C5478 _0472_ _1040_/a_1059_315# 0
C5479 _0461_ _0457_ 0.17242f
C5480 _0225_ _1005_/a_193_47# 0
C5481 _0216_ net111 0
C5482 VPWR _0621_/a_285_297# 0.23911f
C5483 _0190_ _0833_/a_510_47# 0
C5484 _0643_/a_253_47# _0445_ 0
C5485 _1059_/a_193_47# clknet_1_1__leaf__0465_ 0
C5486 _0195_ _0570_/a_373_47# 0
C5487 _0107_ _0324_ 0
C5488 _0216_ _0570_/a_109_297# 0.0091f
C5489 _0118_ _0782_/a_27_47# 0
C5490 net22 net173 0.02796f
C5491 acc0.A\[3\] _0529_/a_109_297# 0
C5492 _0259_ _0818_/a_193_47# 0
C5493 hold99/a_49_47# hold99/a_285_47# 0.22264f
C5494 _0284_ _0346_ 0.22088f
C5495 _0439_ _0290_ 0
C5496 _0140_ _1042_/a_381_47# 0.1253f
C5497 VPWR _1044_/a_381_47# 0.07629f
C5498 _0569_/a_27_297# _0106_ 0
C5499 hold100/a_391_47# _0219_ 0.00219f
C5500 VPWR _0290_ 2.35531f
C5501 _0349_ _1010_/a_1017_47# 0.00172f
C5502 _0127_ _0347_ 0
C5503 acc0.A\[29\] _0352_ 0
C5504 clknet_0__0459_ _1059_/a_1059_315# 0.00369f
C5505 _0732_/a_303_47# _0360_ 0.00139f
C5506 hold39/a_391_47# comp0.B\[0\] 0
C5507 hold35/a_49_47# net2 0
C5508 _0631_/a_109_297# _0262_ 0.00175f
C5509 _0576_/a_27_297# net51 0
C5510 _0470_ hold84/a_285_47# 0.00965f
C5511 _0965_/a_47_47# _0468_ 0
C5512 _0399_ _0347_ 0.57368f
C5513 _0756_/a_377_297# _0378_ 0.00284f
C5514 _0095_ _0405_ 0
C5515 _1001_/a_381_47# _0461_ 0.00265f
C5516 _0285_ _0992_/a_1059_315# 0
C5517 _0983_/a_27_47# _0264_ 0
C5518 _1027_/a_891_413# _1027_/a_1017_47# 0.00617f
C5519 _1027_/a_193_47# net156 0.26008f
C5520 output44/a_27_47# _0340_ 0
C5521 _0606_/a_215_297# _0345_ 0.02926f
C5522 _0764_/a_384_47# control0.add 0
C5523 _0181_ _1067_/a_466_413# 0
C5524 clknet_1_0__leaf__0463_ net173 0.00186f
C5525 hold8/a_285_47# net113 0.01836f
C5526 _0547_/a_150_297# _1040_/a_27_47# 0
C5527 VPWR _0528_/a_81_21# 0.21013f
C5528 hold11/a_391_47# clknet_1_0__leaf__0463_ 0.00814f
C5529 net205 clknet_0__0463_ 0
C5530 net101 _1019_/a_634_159# 0
C5531 _0749_/a_299_297# _0749_/a_384_47# 0
C5532 clknet_1_0__leaf__0462_ _1023_/a_1059_315# 0.00412f
C5533 clknet_0__0460_ _0360_ 0
C5534 _0216_ hold50/a_285_47# 0
C5535 clknet_1_0__leaf__0464_ _1061_/a_1059_315# 0.02633f
C5536 net36 comp0.B\[9\] 0
C5537 _0448_ acc0.A\[15\] 0.00393f
C5538 clknet_0__0458_ _0275_ 0.00839f
C5539 _1052_/a_27_47# _1052_/a_193_47# 0.96066f
C5540 _1032_/a_27_47# _0113_ 0
C5541 net202 _1015_/a_27_47# 0
C5542 control0.reset _1063_/a_634_159# 0
C5543 _0991_/a_891_413# clknet_1_1__leaf__0465_ 0.00207f
C5544 acc0.A\[12\] net42 0.12964f
C5545 _1035_/a_466_413# _0133_ 0.03984f
C5546 _1035_/a_1059_315# net121 0
C5547 _1012_/a_27_47# _1010_/a_27_47# 0
C5548 hold10/a_285_47# _0497_/a_68_297# 0
C5549 _0243_ clkbuf_1_0__f__0461_/a_110_47# 0.00776f
C5550 pp[10] _0156_ 0
C5551 _0094_ _0219_ 0
C5552 _0108_ _0729_/a_68_297# 0
C5553 _1058_/a_193_47# _1058_/a_634_159# 0.11072f
C5554 _1058_/a_27_47# _1058_/a_466_413# 0.27314f
C5555 _0450_ _0843_/a_68_297# 0.00183f
C5556 _0446_ _0843_/a_150_297# 0.00168f
C5557 hold39/a_285_47# _1034_/a_466_413# 0.00148f
C5558 _0329_ _0690_/a_150_297# 0
C5559 hold10/a_49_47# _0499_/a_59_75# 0
C5560 _1000_/a_1017_47# _0247_ 0
C5561 hold69/a_49_47# _0350_ 0.03996f
C5562 _0312_ _0747_/a_510_47# 0
C5563 _1051_/a_1059_315# _0172_ 0.06688f
C5564 _0489_ control0.count\[0\] 0.43621f
C5565 VPWR _0969_/a_109_297# 0.0044f
C5566 net172 A[1] 0
C5567 _1057_/a_27_47# net66 0
C5568 _0172_ _1045_/a_381_47# 0.00553f
C5569 VPWR acc0.A\[1\] 1.08979f
C5570 _0558_/a_68_297# _1035_/a_466_413# 0
C5571 _1050_/a_27_47# _0527_/a_27_297# 0
C5572 clknet_1_1__leaf__0459_ _1013_/a_381_47# 0
C5573 _0680_/a_80_21# _0680_/a_472_297# 0.01636f
C5574 net63 _0619_/a_68_297# 0.00139f
C5575 _0310_ _0780_/a_117_297# 0.00529f
C5576 net117 VPWR 0.35209f
C5577 _0634_/a_113_47# net47 0
C5578 _0230_ _0601_/a_68_297# 0
C5579 _0725_/a_80_21# hold62/a_285_47# 0
C5580 VPWR _0205_ 0.22885f
C5581 net44 _0607_/a_373_47# 0.00164f
C5582 acc0.A\[29\] net115 0.01017f
C5583 _1011_/a_193_47# _0354_ 0.04034f
C5584 _1011_/a_27_47# _0355_ 0.01593f
C5585 _1056_/a_1017_47# _0189_ 0
C5586 clknet_1_0__leaf__0459_ net166 0.26458f
C5587 net46 _0590_/a_113_47# 0
C5588 _0109_ _0350_ 0
C5589 net32 _1043_/a_1059_315# 0
C5590 _0139_ _1043_/a_193_47# 0
C5591 VPWR _0950_/a_75_212# 0.20503f
C5592 _0257_ _0186_ 0.02913f
C5593 _1052_/a_27_47# net12 0.03746f
C5594 net55 hold77/a_391_47# 0.07202f
C5595 _0344_ _0218_ 0.03117f
C5596 _0642_/a_27_413# _0434_ 0
C5597 _1041_/a_975_413# net174 0
C5598 _0179_ _0524_/a_109_47# 0.00142f
C5599 _0174_ _1061_/a_27_47# 0.00195f
C5600 _0346_ _0267_ 0
C5601 net125 _1061_/a_592_47# 0.00107f
C5602 _0974_/a_79_199# clknet_1_0__leaf_clk 0.01f
C5603 _0217_ _0183_ 4.22013f
C5604 comp0.B\[10\] _1061_/a_634_159# 0
C5605 _1027_/a_193_47# acc0.A\[26\] 0.00392f
C5606 net156 _1026_/a_1059_315# 0.00226f
C5607 hold65/a_391_47# _0369_ 0.01419f
C5608 _0195_ _1018_/a_891_413# 0.03105f
C5609 _0346_ _0772_/a_79_21# 0
C5610 net58 _0988_/a_891_413# 0.00143f
C5611 hold77/a_285_47# _0347_ 0.00132f
C5612 _0467_ _1067_/a_381_47# 0
C5613 _0128_ hold62/a_285_47# 0.07478f
C5614 _0349_ _0396_ 0
C5615 hold97/a_285_47# _0319_ 0.01323f
C5616 hold49/a_391_47# _0539_/a_68_297# 0.01025f
C5617 hold15/a_391_47# net162 0.13057f
C5618 clkbuf_0__0462_/a_110_47# _0350_ 0
C5619 _1038_/a_634_159# _0176_ 0.02092f
C5620 _0343_ _0195_ 0.60114f
C5621 _0120_ net151 0.23682f
C5622 _0214_ _0213_ 0.00302f
C5623 _0563_/a_149_47# _0208_ 0
C5624 _0343_ net92 0
C5625 _0530_/a_81_21# _1048_/a_193_47# 0
C5626 output45/a_27_47# _0341_ 0.00643f
C5627 hold59/a_285_47# net206 0.0755f
C5628 hold58/a_391_47# _1034_/a_1059_315# 0.00615f
C5629 _0179_ _0448_ 0.01817f
C5630 init B[2] 0
C5631 net148 _0194_ 0.00663f
C5632 net9 _0196_ 0.23359f
C5633 _0304_ net228 0.03852f
C5634 net59 _1012_/a_634_159# 0
C5635 _0403_ _0993_/a_193_47# 0.00124f
C5636 hold75/a_49_47# _0268_ 0.01674f
C5637 comp0.B\[12\] _0203_ 0
C5638 _1037_/a_193_47# net121 0
C5639 _0399_ clkbuf_0__0465_/a_110_47# 0.04498f
C5640 _0995_/a_634_159# pp[14] 0.00647f
C5641 clknet_1_0__leaf__0465_ input14/a_75_212# 0.06418f
C5642 _0172_ B[7] 0.00297f
C5643 _0982_/a_1017_47# net36 0.00169f
C5644 _0520_/a_27_297# net14 0.17065f
C5645 net89 _0460_ 0
C5646 VPWR _1042_/a_193_47# 0.28147f
C5647 _0629_/a_59_75# _0267_ 0
C5648 net45 _1013_/a_1017_47# 0
C5649 output35/a_27_47# net35 0.1789f
C5650 net61 _0830_/a_510_47# 0
C5651 _1028_/a_27_47# _1008_/a_27_47# 0.00113f
C5652 hold91/a_391_47# net5 0.05034f
C5653 _0285_ _0421_ 0.00495f
C5654 _0401_ _0088_ 0
C5655 clknet_1_1__leaf__0464_ _0204_ 0
C5656 _0388_ VPWR 0.69147f
C5657 _0218_ _0434_ 0
C5658 _0642_/a_27_413# _0989_/a_1059_315# 0
C5659 _0255_ net73 0.0021f
C5660 pp[27] _1030_/a_1059_315# 0.0019f
C5661 _0988_/a_27_47# _0988_/a_634_159# 0.14145f
C5662 _0500_/a_27_47# clkbuf_1_1__f__0457_/a_110_47# 0
C5663 _0352_ _0754_/a_512_297# 0.00216f
C5664 _1039_/a_27_47# _0174_ 0
C5665 _1039_/a_1059_315# _0553_/a_240_47# 0
C5666 pp[18] _1013_/a_27_47# 0
C5667 _0199_ net9 0.00565f
C5668 clknet_0__0462_ clknet_1_1__leaf__0462_ 0.00537f
C5669 _0217_ acc0.A\[15\] 0
C5670 clknet_1_1__leaf__0460_ _1010_/a_466_413# 0
C5671 net240 clknet_1_0__leaf__0460_ 0.21269f
C5672 _0295_ _0347_ 0.05984f
C5673 net10 _1043_/a_1059_315# 0.02802f
C5674 hold20/a_49_47# _0490_ 0
C5675 hold21/a_391_47# hold22/a_49_47# 0.00222f
C5676 hold21/a_285_47# hold22/a_285_47# 0.00385f
C5677 net202 _0215_ 0
C5678 _0542_/a_51_297# _0542_/a_512_297# 0.0116f
C5679 _0967_/a_215_297# _1064_/a_1059_315# 0.00129f
C5680 acc0.A\[3\] net170 0.05935f
C5681 _0162_ _1064_/a_466_413# 0.00472f
C5682 _0485_ _1064_/a_381_47# 0
C5683 _0487_ _1064_/a_891_413# 0
C5684 pp[9] net179 0
C5685 hold52/a_391_47# _0123_ 0
C5686 hold52/a_49_47# net200 0
C5687 net171 _0173_ 0.01184f
C5688 clknet_1_1__leaf__0463_ _0215_ 0.34324f
C5689 net122 _0175_ 0
C5690 _1026_/a_1059_315# acc0.A\[26\] 0.08864f
C5691 hold94/a_49_47# net51 0.2917f
C5692 _0465_ _1047_/a_561_413# 0
C5693 _0480_ _0486_ 0
C5694 _0224_ _0592_/a_68_297# 0.11141f
C5695 _1072_/a_891_413# _0486_ 0
C5696 _0880_/a_27_47# _1062_/a_27_47# 0
C5697 _0322_ _0324_ 0.07107f
C5698 _0356_ _0725_/a_209_47# 0
C5699 VPWR _0562_/a_68_297# 0.16016f
C5700 _0817_/a_266_47# _0817_/a_585_47# 0.0013f
C5701 clknet_1_1__leaf__0460_ _1009_/a_1059_315# 0.02176f
C5702 _0242_ _0771_/a_215_297# 0.01118f
C5703 _0349_ _0348_ 0.00446f
C5704 _0981_/a_27_297# _0484_ 0.00406f
C5705 clknet_1_1__leaf__0458_ _0988_/a_466_413# 0
C5706 _0327_ _0324_ 0.35834f
C5707 _0290_ _0283_ 0
C5708 _0982_/a_27_47# hold60/a_285_47# 0
C5709 _0982_/a_193_47# hold60/a_49_47# 0
C5710 pp[26] _0571_/a_109_47# 0.00295f
C5711 net153 _1040_/a_27_47# 0
C5712 _0787_/a_80_21# _0787_/a_209_297# 0.06257f
C5713 net40 output40/a_27_47# 0.17325f
C5714 hold47/a_49_47# net154 0.01091f
C5715 net78 clkbuf_1_1__f__0465_/a_110_47# 0.01192f
C5716 _0461_ _0614_/a_29_53# 0
C5717 net11 _0186_ 0.34614f
C5718 clkbuf_1_1__f__0465_/a_110_47# clknet_0__0465_ 0.31304f
C5719 net24 _0173_ 0.00808f
C5720 hold76/a_391_47# _0241_ 0.02598f
C5721 _0229_ _0219_ 0.07182f
C5722 _0789_/a_315_47# _0405_ 0
C5723 _0343_ _0081_ 0.03067f
C5724 _0429_ _0186_ 0
C5725 comp0.B\[4\] net25 0.02978f
C5726 net43 _0790_/a_35_297# 0
C5727 net189 net143 0.00114f
C5728 _0174_ _1040_/a_975_413# 0
C5729 _0136_ _1040_/a_466_413# 0
C5730 _0458_ _0345_ 0
C5731 _1037_/a_634_159# _1037_/a_592_47# 0
C5732 _0504_/a_27_47# clknet_1_0__leaf__0458_ 0.03278f
C5733 _0997_/a_27_47# _0218_ 0.00102f
C5734 _0350_ acc0.A\[6\] 0
C5735 _0195_ _0998_/a_193_47# 0.04516f
C5736 acc0.A\[22\] _0379_ 0
C5737 _1008_/a_1059_315# _0687_/a_59_75# 0.00755f
C5738 comp0.B\[10\] _1040_/a_1017_47# 0
C5739 pp[30] _1030_/a_27_47# 0.03548f
C5740 net59 _1030_/a_634_159# 0
C5741 clknet_1_0__leaf__0458_ _0456_ 0
C5742 VPWR _1005_/a_381_47# 0.08423f
C5743 _0227_ acc0.A\[23\] 0
C5744 clknet_1_1__leaf__0459_ hold91/a_285_47# 0
C5745 _0790_/a_285_47# _0406_ 0.00223f
C5746 _0343_ _0505_/a_373_47# 0
C5747 VPWR net77 0.37752f
C5748 _0985_/a_27_47# _0447_ 0
C5749 _0157_ _0287_ 0
C5750 net234 _0854_/a_79_21# 0
C5751 clkbuf_1_1__f__0462_/a_110_47# _1010_/a_1059_315# 0
C5752 _0349_ _0332_ 0
C5753 _1054_/a_975_413# _0180_ 0
C5754 clknet_1_0__leaf__0462_ _0219_ 0.00547f
C5755 output39/a_27_47# _0994_/a_891_413# 0.01654f
C5756 _1001_/a_27_47# _1001_/a_634_159# 0.14145f
C5757 _0390_ _0388_ 0
C5758 _0621_/a_35_297# acc0.A\[6\] 0.10929f
C5759 _0100_ net1 0.02439f
C5760 pp[28] _1030_/a_466_413# 0
C5761 VPWR _0223_ 0.52893f
C5762 net160 clknet_0__0463_ 0
C5763 net7 hold6/a_285_47# 0
C5764 _0984_/a_27_47# clknet_1_1__leaf__0465_ 0
C5765 _0217_ hold40/a_285_47# 0.0159f
C5766 VPWR _0765_/a_215_47# 0.00587f
C5767 _0717_/a_209_297# _0333_ 0.03686f
C5768 _1039_/a_592_47# _0473_ 0
C5769 _0608_/a_27_47# _0677_/a_285_47# 0
C5770 hold9/a_391_47# _1008_/a_1059_315# 0
C5771 hold9/a_285_47# _1008_/a_891_413# 0.00219f
C5772 hold7/a_391_47# _0186_ 0
C5773 _0831_/a_35_297# _0831_/a_117_297# 0.00641f
C5774 _0235_ _0764_/a_299_297# 0
C5775 _0808_/a_81_21# net246 0
C5776 _0198_ _0531_/a_373_47# 0
C5777 _0146_ _0531_/a_27_297# 0.08652f
C5778 net45 net83 0.00317f
C5779 _1049_/a_1059_315# _1048_/a_27_47# 0.01216f
C5780 _1049_/a_193_47# _1048_/a_466_413# 0
C5781 _1049_/a_466_413# _1048_/a_193_47# 0.00121f
C5782 hold44/a_391_47# net191 0.13065f
C5783 hold8/a_49_47# hold8/a_391_47# 0.00188f
C5784 hold14/a_49_47# _1037_/a_27_47# 0
C5785 hold54/a_285_47# _0113_ 0.0012f
C5786 B[9] comp0.B\[11\] 0
C5787 _0254_ _0831_/a_35_297# 0
C5788 VPWR _1006_/a_1059_315# 0.41934f
C5789 _0271_ _0826_/a_27_53# 0.00118f
C5790 VPWR _0656_/a_59_75# 0.22813f
C5791 _1029_/a_381_47# _1008_/a_27_47# 0
C5792 _1029_/a_27_47# _1008_/a_381_47# 0
C5793 _0476_ _0474_ 0.25441f
C5794 clkload1/Y _0270_ 0
C5795 _0453_ acc0.A\[1\] 0.00271f
C5796 _0181_ _0580_/a_27_297# 0
C5797 _1055_/a_1059_315# A[10] 0
C5798 net45 _0781_/a_68_297# 0.00144f
C5799 _0307_ _0097_ 0
C5800 _0195_ _1030_/a_381_47# 0.00699f
C5801 net48 _1005_/a_381_47# 0.00207f
C5802 hold49/a_285_47# net21 0
C5803 VPWR _0986_/a_1059_315# 0.42473f
C5804 _1046_/a_193_47# _1061_/a_27_47# 0
C5805 _0293_ net67 0
C5806 _0714_/a_51_297# _0219_ 0.19542f
C5807 _0714_/a_240_47# _0345_ 0
C5808 _0550_/a_149_47# _0176_ 0.00579f
C5809 pp[9] _1058_/a_634_159# 0
C5810 net118 _1067_/a_891_413# 0
C5811 _0501_/a_27_47# control0.sh 0.00121f
C5812 _0185_ _0505_/a_27_297# 0.00108f
C5813 _0951_/a_209_311# _0951_/a_296_53# 0.0049f
C5814 _0179_ _0142_ 0.0107f
C5815 _1013_/a_193_47# _0567_/a_109_297# 0
C5816 _1013_/a_634_159# _0567_/a_27_297# 0
C5817 _0701_/a_209_297# _0332_ 0.00894f
C5818 input15/a_75_212# A[8] 0.21182f
C5819 _0161_ hold93/a_285_47# 0.00102f
C5820 _1004_/a_193_47# _0216_ 0.02893f
C5821 _0175_ _0560_/a_150_297# 0
C5822 net126 net36 0
C5823 net48 _0765_/a_215_47# 0
C5824 _1072_/a_27_47# _1068_/a_634_159# 0
C5825 _1072_/a_193_47# _1068_/a_193_47# 0
C5826 _1072_/a_634_159# _1068_/a_27_47# 0
C5827 _0388_ clknet_1_0__leaf__0459_ 0
C5828 _0180_ _0522_/a_109_47# 0.0019f
C5829 _0689_/a_68_297# _0319_ 0.17718f
C5830 output36/a_27_47# A[1] 0.01105f
C5831 net36 input8/a_75_212# 0
C5832 _0527_/a_27_297# _0987_/a_27_47# 0
C5833 hold46/a_49_47# _0201_ 0
C5834 comp0.B\[13\] _0538_/a_512_297# 0
C5835 _0957_/a_32_297# _0561_/a_240_47# 0
C5836 net95 _1009_/a_381_47# 0
C5837 _0252_ _0833_/a_79_21# 0
C5838 _0316_ _0322_ 0.21839f
C5839 net55 _0329_ 0
C5840 _0292_ _0288_ 0.33573f
C5841 _0287_ acc0.A\[9\] 0.00367f
C5842 _1003_/a_891_413# _0227_ 0
C5843 acc0.A\[14\] _0301_ 0
C5844 net47 clknet_1_0__leaf__0457_ 0
C5845 _0478_ _1072_/a_193_47# 0
C5846 net45 _0216_ 0.013f
C5847 _0316_ _0327_ 0.24058f
C5848 _1035_/a_466_413# _0208_ 0
C5849 _1035_/a_193_47# _0132_ 0
C5850 _0133_ _0561_/a_51_297# 0.03573f
C5851 _0272_ _0274_ 0.16686f
C5852 _1047_/a_27_47# _1047_/a_1059_315# 0.04875f
C5853 _1047_/a_193_47# _1047_/a_466_413# 0.07537f
C5854 _1030_/a_27_47# _0339_ 0.01741f
C5855 clknet_1_1__leaf__0458_ _0186_ 0.54549f
C5856 _0206_ _1040_/a_891_413# 0.0313f
C5857 comp0.B\[8\] _1040_/a_381_47# 0.01316f
C5858 hold97/a_391_47# _0317_ 0
C5859 hold1/a_391_47# _0987_/a_27_47# 0.00109f
C5860 _0957_/a_32_297# _0472_ 0.0642f
C5861 _0957_/a_220_297# _0473_ 0
C5862 net101 net105 0.01055f
C5863 _0371_ net52 0.21341f
C5864 net47 _0988_/a_1059_315# 0.01771f
C5865 control0.add hold40/a_391_47# 0
C5866 clknet_1_0__leaf__0460_ hold3/a_285_47# 0.00153f
C5867 _1041_/a_466_413# _0174_ 0.00115f
C5868 _0327_ _0347_ 0.03393f
C5869 _0664_/a_382_297# _0664_/a_297_47# 0
C5870 hold5/a_285_47# hold51/a_49_47# 0
C5871 net40 net81 0
C5872 output57/a_27_47# VPWR 0.29857f
C5873 net133 net147 0
C5874 _1041_/a_891_413# comp0.B\[10\] 0.00213f
C5875 net234 _1014_/a_193_47# 0.00259f
C5876 net55 _0221_ 0.06317f
C5877 net178 _0517_/a_81_21# 0.10863f
C5878 _1007_/a_466_413# _1007_/a_561_413# 0.00772f
C5879 _1007_/a_634_159# _1007_/a_975_413# 0
C5880 _1052_/a_466_413# _1052_/a_592_47# 0.00553f
C5881 _1052_/a_634_159# _1052_/a_1017_47# 0
C5882 hold22/a_49_47# _0519_/a_81_21# 0
C5883 _0253_ _0988_/a_27_47# 0
C5884 hold96/a_391_47# _1004_/a_193_47# 0
C5885 hold96/a_285_47# _1004_/a_634_159# 0.01555f
C5886 VPWR _0854_/a_297_297# 0.01145f
C5887 _0177_ _1061_/a_634_159# 0.00518f
C5888 _0432_ _0835_/a_78_199# 0.20028f
C5889 _0837_/a_368_297# _0837_/a_266_47# 0.00153f
C5890 _0501_/a_27_47# net157 0
C5891 _1058_/a_1059_315# _1058_/a_1017_47# 0
C5892 _1058_/a_193_47# net144 0.01326f
C5893 _0172_ _1044_/a_891_413# 0.04336f
C5894 _1020_/a_634_159# _0352_ 0.011f
C5895 hold69/a_285_47# _1006_/a_193_47# 0
C5896 hold69/a_391_47# _1006_/a_27_47# 0
C5897 _0179_ _1052_/a_891_413# 0.01564f
C5898 net197 _1027_/a_27_47# 0
C5899 _0178_ _0935_/a_27_47# 0
C5900 _1021_/a_27_47# clknet_1_0__leaf__0461_ 0.00691f
C5901 clknet_0__0463_ acc0.A\[15\] 0.00241f
C5902 VPWR B[8] 0.19402f
C5903 _0257_ net62 0.07942f
C5904 _0558_/a_68_297# _0133_ 0
C5905 _0705_/a_59_75# _0705_/a_145_75# 0.00658f
C5906 _1050_/a_891_413# net154 0.0034f
C5907 _0459_ net221 0.00601f
C5908 _1003_/a_193_47# _0487_ 0.00497f
C5909 _0971_/a_81_21# _0971_/a_384_47# 0.00138f
C5910 input22/a_75_212# net22 0.10977f
C5911 _0216_ _0726_/a_51_297# 0.01882f
C5912 _1011_/a_1017_47# net227 0
C5913 VPWR _1013_/a_1017_47# 0
C5914 _1033_/a_634_159# control0.reset 0.01746f
C5915 _1002_/a_975_413# VPWR 0.00494f
C5916 _1061_/a_27_47# comp0.B\[9\] 0
C5917 comp0.B\[11\] hold6/a_285_47# 0
C5918 clkbuf_0_clk/a_110_47# _1063_/a_193_47# 0.00177f
C5919 net61 _0989_/a_193_47# 0.00504f
C5920 _0243_ _0616_/a_78_199# 0
C5921 clkbuf_1_0__f__0462_/a_110_47# hold90/a_49_47# 0.01547f
C5922 hold75/a_49_47# net222 0
C5923 net114 _0345_ 0
C5924 _0617_/a_150_297# _1006_/a_27_47# 0
C5925 _0983_/a_27_47# _0454_ 0.05458f
C5926 _0617_/a_68_297# _1006_/a_193_47# 0
C5927 net169 _0519_/a_81_21# 0
C5928 _0201_ comp0.B\[14\] 0.18103f
C5929 clkload4/Y hold19/a_49_47# 0.00464f
C5930 _1059_/a_193_47# _0277_ 0
C5931 clknet_0_clk _0468_ 0.44473f
C5932 _1063_/a_27_47# _1063_/a_466_413# 0.26005f
C5933 _1063_/a_193_47# _1063_/a_634_159# 0.11072f
C5934 _0504_/a_27_47# hold18/a_49_47# 0
C5935 _1058_/a_891_413# _0186_ 0.00201f
C5936 _0645_/a_47_47# acc0.A\[15\] 0.01279f
C5937 _0645_/a_377_297# net42 0
C5938 _0197_ _0447_ 0
C5939 net99 clknet_1_1__leaf__0461_ 0.15167f
C5940 _0463_ comp0.B\[5\] 0.00134f
C5941 _1019_/a_27_47# _0346_ 0.03683f
C5942 comp0.B\[10\] net147 0.00431f
C5943 clkbuf_1_0__f__0459_/a_110_47# _0195_ 0
C5944 _1027_/a_1059_315# hold50/a_391_47# 0
C5945 _1027_/a_891_413# hold50/a_285_47# 0
C5946 _1037_/a_27_47# _0208_ 0
C5947 _0788_/a_68_297# _0403_ 0.17733f
C5948 clknet_1_0__leaf__0463_ input22/a_75_212# 0
C5949 acc0.A\[20\] _0772_/a_297_297# 0
C5950 _0195_ _0147_ 0.23546f
C5951 _0786_/a_80_21# _0402_ 0.1187f
C5952 net63 _0346_ 0.12995f
C5953 _0456_ hold18/a_49_47# 0.01554f
C5954 _0310_ clkbuf_1_1__f__0461_/a_110_47# 0
C5955 _1063_/a_1059_315# clknet_1_0__leaf__0457_ 0.00549f
C5956 net124 _0176_ 0
C5957 output43/a_27_47# _0218_ 0.00295f
C5958 net37 _0418_ 0
C5959 net199 _0216_ 0.1296f
C5960 hold34/a_391_47# acc0.A\[10\] 0
C5961 _1039_/a_634_159# _0177_ 0
C5962 _0536_/a_240_47# clkbuf_0__0464_/a_110_47# 0
C5963 net158 _1049_/a_193_47# 0
C5964 net63 net65 0.05154f
C5965 _0984_/a_975_413# VPWR 0.00502f
C5966 _0336_ hold92/a_391_47# 0
C5967 net63 _0989_/a_466_413# 0
C5968 input20/a_75_212# comp0.B\[10\] 0
C5969 _0994_/a_1017_47# _0218_ 0
C5970 clknet_0__0461_ net102 0
C5971 clknet_0__0459_ _0670_/a_297_297# 0
C5972 _0305_ net43 0.04335f
C5973 _0354_ _0707_/a_75_199# 0.0012f
C5974 _1011_/a_466_413# acc0.A\[29\] 0.00416f
C5975 _1004_/a_466_413# net90 0
C5976 hold57/a_285_47# _0209_ 0
C5977 _1004_/a_193_47# _1024_/a_193_47# 0
C5978 _1004_/a_27_47# _1024_/a_634_159# 0
C5979 _0183_ _0583_/a_373_47# 0.00135f
C5980 _0369_ _0990_/a_891_413# 0.0013f
C5981 _0732_/a_80_21# _0366_ 0.06867f
C5982 _0143_ _0174_ 0
C5983 _0306_ _0347_ 0.04995f
C5984 _1002_/a_975_413# net48 0
C5985 VPWR _0704_/a_68_297# 0.15562f
C5986 _0982_/a_592_47# _0346_ 0.00104f
C5987 _1060_/a_27_47# _1060_/a_466_413# 0.27314f
C5988 _1060_/a_193_47# _1060_/a_634_159# 0.11072f
C5989 _0510_/a_27_297# acc0.A\[10\] 0.14626f
C5990 hold43/a_391_47# _1028_/a_193_47# 0
C5991 net15 acc0.A\[7\] 0.07531f
C5992 net40 _0797_/a_207_413# 0.00314f
C5993 pp[27] VPWR 0.75007f
C5994 net45 _0608_/a_109_297# 0
C5995 pp[26] net155 0.15576f
C5996 net196 _1042_/a_891_413# 0.00557f
C5997 _1039_/a_27_47# comp0.B\[9\] 0
C5998 _0143_ _1050_/a_27_47# 0
C5999 _0850_/a_68_297# net47 0.12404f
C6000 hold47/a_49_47# clknet_0__0464_ 0
C6001 _1030_/a_592_47# acc0.A\[30\] 0
C6002 _0805_/a_27_47# acc0.A\[11\] 0
C6003 hold56/a_49_47# _1065_/a_1059_315# 0
C6004 hold56/a_391_47# _1065_/a_634_159# 0
C6005 clknet_1_1__leaf__0463_ _0955_/a_304_297# 0
C6006 _0365_ _0345_ 0.0477f
C6007 _0988_/a_891_413# _0988_/a_975_413# 0.00851f
C6008 _0988_/a_27_47# net74 0.2288f
C6009 _0988_/a_381_47# _0988_/a_561_413# 0.00123f
C6010 _0787_/a_209_297# _0402_ 0.03795f
C6011 _0118_ hold55/a_285_47# 0
C6012 _0553_/a_245_297# _0553_/a_240_47# 0
C6013 net22 clknet_1_1__leaf__0457_ 0
C6014 _0967_/a_109_93# _0471_ 0
C6015 _0671_/a_113_297# _0302_ 0.01738f
C6016 _0487_ _0471_ 0.06281f
C6017 _1053_/a_1059_315# acc0.A\[7\] 0.08503f
C6018 clk _1062_/a_634_159# 0
C6019 clkbuf_0_clk/a_110_47# _1062_/a_891_413# 0
C6020 _0174_ _0953_/a_32_297# 0
C6021 _0357_ _0108_ 0.00101f
C6022 _0820_/a_79_21# net76 0
C6023 _0331_ _0350_ 0.13413f
C6024 net125 comp0.B\[10\] 0
C6025 _0947_/a_109_297# control0.state\[2\] 0.00285f
C6026 _1041_/a_27_47# _0206_ 0
C6027 _1041_/a_193_47# comp0.B\[8\] 0
C6028 output37/a_27_47# pp[10] 0.35271f
C6029 VPWR _0198_ 0.36473f
C6030 _0982_/a_1059_315# _0465_ 0.00388f
C6031 _0753_/a_79_21# _0378_ 0.01441f
C6032 _0953_/a_220_297# comp0.B\[10\] 0.00325f
C6033 _0606_/a_109_53# hold94/a_285_47# 0
C6034 _0606_/a_215_297# hold94/a_391_47# 0
C6035 VPWR _1014_/a_634_159# 0.1838f
C6036 net58 hold100/a_391_47# 0.05189f
C6037 _0325_ clknet_1_0__leaf__0460_ 0.00187f
C6038 _0323_ _0326_ 0.11218f
C6039 _0542_/a_51_297# _0141_ 0.10639f
C6040 _0542_/a_240_47# net195 0.04783f
C6041 _0542_/a_149_47# net19 0.00138f
C6042 _0366_ _0250_ 0
C6043 _0176_ _0494_/a_27_47# 0
C6044 hold96/a_391_47# net199 0
C6045 clknet_1_0__leaf__0465_ _0826_/a_27_53# 0
C6046 _0982_/a_466_413# net58 0
C6047 _1001_/a_592_47# clknet_1_0__leaf__0457_ 0
C6048 _0163_ _0951_/a_109_93# 0
C6049 net82 _1060_/a_193_47# 0
C6050 clknet_0__0457_ net234 0
C6051 _0172_ _1042_/a_27_47# 0
C6052 clknet_1_0__leaf__0463_ clknet_1_1__leaf__0457_ 0.00662f
C6053 _0467_ net231 0
C6054 hold14/a_49_47# _0133_ 0
C6055 hold14/a_285_47# net121 0.01875f
C6056 _0216_ _0584_/a_109_297# 0.04264f
C6057 net121 input27/a_75_212# 0
C6058 _1021_/a_381_47# clknet_1_0__leaf__0457_ 0.00314f
C6059 _1021_/a_1059_315# _0460_ 0.00765f
C6060 _0170_ _0484_ 0
C6061 _0701_/a_209_297# _0701_/a_209_47# 0
C6062 _0701_/a_80_21# _0701_/a_303_47# 0.01146f
C6063 net133 _1047_/a_1059_315# 0
C6064 net46 _0240_ 0.00536f
C6065 B[15] net27 0
C6066 net23 B[4] 0.19776f
C6067 clknet_1_1__leaf__0462_ _0687_/a_59_75# 0.00143f
C6068 clkbuf_0__0462_/a_110_47# _0737_/a_285_297# 0
C6069 _1067_/a_27_47# clkbuf_1_1__f_clk/a_110_47# 0.01577f
C6070 _0181_ acc0.A\[10\] 0.12558f
C6071 clkbuf_1_1__f__0462_/a_110_47# clkbuf_1_1__f__0460_/a_110_47# 0.03464f
C6072 pp[17] net59 0
C6073 _0580_/a_373_47# acc0.A\[19\] 0
C6074 net46 _0369_ 0.43203f
C6075 net44 pp[30] 0.10318f
C6076 clkbuf_0__0464_/a_110_47# _1046_/a_27_47# 0.0304f
C6077 hold73/a_49_47# hold73/a_285_47# 0.22264f
C6078 clknet_0__0457_ net46 0
C6079 VPWR net83 0.38158f
C6080 hold79/a_49_47# _0167_ 0
C6081 hold79/a_285_47# clknet_1_0__leaf_clk 0.07903f
C6082 _1008_/a_1059_315# _0739_/a_215_47# 0
C6083 clknet_1_1__leaf__0460_ _0367_ 0.23192f
C6084 _0405_ _0219_ 0.14058f
C6085 _0408_ _0345_ 0.14653f
C6086 _0559_/a_51_297# _0557_/a_51_297# 0.07173f
C6087 _0557_/a_240_47# _0175_ 0
C6088 _0347_ _1008_/a_561_413# 0
C6089 _0228_ _0381_ 0.03034f
C6090 _0136_ net174 0
C6091 _1037_/a_975_413# _0135_ 0
C6092 net16 _0189_ 0
C6093 net175 _1048_/a_27_47# 0.00133f
C6094 _0356_ _0219_ 0.08152f
C6095 _0596_/a_59_75# VPWR 0.21477f
C6096 hold25/a_285_47# _1038_/a_27_47# 0
C6097 hold25/a_49_47# _1038_/a_193_47# 0.01238f
C6098 _0238_ clknet_1_0__leaf__0460_ 0.3137f
C6099 VPWR _0781_/a_68_297# 0.14707f
C6100 hold96/a_285_47# net46 0
C6101 net231 comp0.B\[0\] 0.09456f
C6102 _0465_ _0451_ 0.00284f
C6103 _0276_ _0794_/a_27_47# 0
C6104 _0396_ clknet_1_1__leaf__0461_ 0
C6105 _0538_/a_51_297# _1045_/a_193_47# 0.0021f
C6106 output66/a_27_47# input2/a_75_212# 0.00713f
C6107 _0291_ _0345_ 0
C6108 _0467_ hold38/a_285_47# 0
C6109 _0814_/a_27_47# _0291_ 0
C6110 clknet_1_0__leaf_clk net17 0
C6111 clknet_1_1__leaf__0460_ _0680_/a_80_21# 0.07896f
C6112 _0664_/a_297_47# _0402_ 0.02853f
C6113 _0728_/a_59_75# _0356_ 0.18568f
C6114 hold9/a_49_47# net113 0
C6115 hold9/a_391_47# clknet_1_1__leaf__0462_ 0.01319f
C6116 _0553_/a_51_297# _0173_ 0
C6117 _0698_/a_113_297# _0319_ 0.08447f
C6118 hold30/a_49_47# acc0.A\[23\] 0
C6119 input1/a_27_47# rst 0
C6120 A[0] input34/a_27_47# 0.00343f
C6121 _1001_/a_634_159# _0772_/a_79_21# 0
C6122 _1001_/a_381_47# _1001_/a_561_413# 0.00123f
C6123 _1001_/a_891_413# _1001_/a_975_413# 0.00851f
C6124 _0537_/a_150_297# clknet_1_1__leaf__0464_ 0
C6125 _0991_/a_634_159# _0345_ 0
C6126 net1 _0972_/a_93_21# 0
C6127 _0115_ _1060_/a_193_47# 0
C6128 _1035_/a_193_47# net25 0.00586f
C6129 _0399_ _0180_ 0
C6130 _1062_/a_634_159# _1062_/a_592_47# 0
C6131 _0487_ hold93/a_391_47# 0.00254f
C6132 clkbuf_1_1__f__0459_/a_110_47# _0795_/a_81_21# 0
C6133 _1011_/a_193_47# _0353_ 0
C6134 _0992_/a_1059_315# net228 0.0016f
C6135 _0473_ comp0.B\[10\] 0.01849f
C6136 hold38/a_285_47# comp0.B\[0\] 0.00103f
C6137 acc0.A\[9\] input16/a_75_212# 0.0556f
C6138 _1021_/a_27_47# _1021_/a_561_413# 0.0027f
C6139 _1021_/a_634_159# _1021_/a_891_413# 0.03684f
C6140 _1021_/a_193_47# _1021_/a_381_47# 0.09503f
C6141 _0239_ clkbuf_1_1__f__0461_/a_110_47# 0.00121f
C6142 _1033_/a_27_47# net23 0
C6143 _1003_/a_561_413# net49 0
C6144 hold41/a_49_47# net188 0
C6145 control0.add acc0.A\[19\] 0.25783f
C6146 net199 _1024_/a_193_47# 0
C6147 _0518_/a_109_47# clknet_1_1__leaf__0458_ 0.00332f
C6148 _1017_/a_27_47# _0459_ 0.00348f
C6149 _0147_ _1048_/a_193_47# 0
C6150 _1049_/a_634_159# net134 0.0014f
C6151 _0352_ acc0.A\[23\] 0.26069f
C6152 _0476_ _0563_/a_51_297# 0
C6153 _0645_/a_47_47# _0645_/a_129_47# 0.00369f
C6154 _0216_ VPWR 9.73713f
C6155 _0510_/a_27_297# _0510_/a_109_297# 0.17136f
C6156 _0996_/a_891_413# _0670_/a_79_21# 0
C6157 _0459_ _1060_/a_975_413# 0
C6158 hold64/a_285_47# net45 0
C6159 net152 _0545_/a_68_297# 0
C6160 _0530_/a_81_21# acc0.A\[15\] 0
C6161 _0432_ _0399_ 0
C6162 _0346_ _0347_ 0.66823f
C6163 VPWR _0548_/a_149_47# 0.00189f
C6164 VPWR clknet_1_1__leaf__0464_ 2.99018f
C6165 clkbuf_1_0__f__0465_/a_110_47# _0989_/a_634_159# 0
C6166 _0195_ clkbuf_0__0461_/a_110_47# 0
C6167 control0.state\[0\] control0.state\[2\] 0.34177f
C6168 _0234_ _0756_/a_285_47# 0
C6169 _0195_ _0568_/a_27_297# 0.14646f
C6170 net43 _0181_ 0
C6171 _0216_ _1015_/a_466_413# 0.00443f
C6172 _0996_/a_27_47# _0369_ 0
C6173 _0891_/a_27_47# comp0.B\[1\] 0
C6174 net225 _0219_ 0.08572f
C6175 pp[9] net144 0
C6176 _0817_/a_266_47# _0816_/a_68_297# 0
C6177 _0628_/a_109_297# VPWR 0.00649f
C6178 _0185_ _0184_ 0.03625f
C6179 _1034_/a_193_47# clknet_0__0463_ 0.00389f
C6180 _1034_/a_1059_315# clkbuf_1_1__f__0463_/a_110_47# 0.00113f
C6181 _0092_ _0994_/a_381_47# 0.11464f
C6182 _0130_ _0461_ 0
C6183 hold26/a_49_47# net152 0
C6184 hold38/a_285_47# _1034_/a_634_159# 0
C6185 _0104_ _0346_ 0.18415f
C6186 _0225_ _1022_/a_1059_315# 0
C6187 hold17/a_49_47# _1071_/a_27_47# 0.01463f
C6188 net46 _1024_/a_27_47# 0
C6189 _0561_/a_240_47# _0213_ 0
C6190 _0561_/a_149_47# _0173_ 0.02579f
C6191 _0561_/a_51_297# _0208_ 0.13411f
C6192 control0.add _0249_ 0
C6193 VPWR _1067_/a_27_47# 0.70804f
C6194 net82 _0796_/a_79_21# 0.01f
C6195 hold29/a_391_47# _1022_/a_27_47# 0
C6196 hold100/a_49_47# _0263_ 0.04455f
C6197 hold100/a_285_47# _0261_ 0.05516f
C6198 hold90/a_285_47# _0105_ 0
C6199 _0487_ control0.reset 0
C6200 net53 _0733_/a_79_199# 0.00928f
C6201 _0313_ _0743_/a_51_297# 0.0016f
C6202 _0515_/a_299_297# net2 0.07965f
C6203 _0241_ clknet_1_0__leaf__0461_ 0.03144f
C6204 _0982_/a_193_47# _0263_ 0
C6205 _0982_/a_634_159# _0261_ 0
C6206 pp[17] _0335_ 0
C6207 net44 _0339_ 0.04599f
C6208 net62 clknet_1_1__leaf__0458_ 0.10302f
C6209 _0640_/a_215_297# _0271_ 0.03025f
C6210 _0869_/a_27_47# net223 0.00103f
C6211 _1020_/a_634_159# net106 0
C6212 _0182_ net71 0.04173f
C6213 _0618_/a_79_21# _0618_/a_510_47# 0.00844f
C6214 _0618_/a_297_297# _0618_/a_215_47# 0
C6215 comp0.B\[13\] _0143_ 0
C6216 _0472_ _0213_ 0.15962f
C6217 hold39/a_285_47# _0175_ 0.01503f
C6218 _1036_/a_381_47# net122 0
C6219 _1036_/a_975_413# clknet_1_1__leaf__0463_ 0
C6220 _0346_ _0792_/a_209_297# 0
C6221 _1050_/a_891_413# clknet_0__0464_ 0
C6222 _0348_ _1030_/a_193_47# 0
C6223 _0510_/a_109_297# _0181_ 0.01895f
C6224 _0644_/a_47_47# _0304_ 0
C6225 _0461_ _1019_/a_381_47# 0.00325f
C6226 hold96/a_391_47# VPWR 0.17828f
C6227 _0290_ _0345_ 0.04725f
C6228 _0290_ _0814_/a_27_47# 0.08066f
C6229 _0423_ _0814_/a_109_47# 0
C6230 VPWR _0852_/a_285_297# 0.24869f
C6231 _1001_/a_466_413# _0218_ 0
C6232 _0133_ _0208_ 0.29649f
C6233 _1041_/a_381_47# net153 0.12992f
C6234 _1041_/a_466_413# comp0.B\[9\] 0
C6235 _0350_ _1008_/a_27_47# 0.00298f
C6236 _1047_/a_891_413# _1047_/a_1017_47# 0.00617f
C6237 _1047_/a_193_47# _0145_ 0.43174f
C6238 _0322_ _0106_ 0
C6239 _0083_ clknet_0__0458_ 0
C6240 clknet_1_1__leaf__0460_ _0742_/a_299_297# 0
C6241 input12/a_75_212# net11 0.11082f
C6242 hold12/a_49_47# _0237_ 0
C6243 hold12/a_285_47# _0381_ 0
C6244 _0401_ _0304_ 0
C6245 _0425_ _0295_ 0
C6246 clknet_0__0465_ _0826_/a_301_297# 0
C6247 _0131_ _0214_ 0.0239f
C6248 _0271_ _0465_ 0.01375f
C6249 _0212_ _0561_/a_240_47# 0
C6250 _0849_/a_215_47# _0219_ 0.0503f
C6251 control0.state\[1\] _0467_ 0.02456f
C6252 _0973_/a_109_297# clknet_1_0__leaf__0461_ 0
C6253 _0479_ _1072_/a_27_47# 0
C6254 pp[28] net227 0.00332f
C6255 net188 _0513_/a_299_297# 0.06355f
C6256 hold41/a_49_47# _0155_ 0
C6257 _0183_ _1018_/a_891_413# 0
C6258 _0855_/a_81_21# acc0.A\[0\] 0.00146f
C6259 _0953_/a_32_297# _1046_/a_193_47# 0
C6260 hold85/a_285_47# _0959_/a_217_297# 0
C6261 _1004_/a_193_47# _0756_/a_377_297# 0
C6262 _0390_ _0216_ 0
C6263 _0536_/a_149_47# _0473_ 0.00631f
C6264 _0536_/a_245_297# _0472_ 0
C6265 acc0.A\[31\] clknet_1_1__leaf__0461_ 0
C6266 _0525_/a_81_21# net13 0.01198f
C6267 _0177_ net147 0
C6268 net62 _0263_ 0
C6269 _0233_ _0217_ 0
C6270 _0343_ _0183_ 0.12439f
C6271 _0805_/a_27_47# _0281_ 0.20826f
C6272 _0450_ _0263_ 0.31223f
C6273 _0305_ _0677_/a_129_47# 0.00233f
C6274 B[11] net195 0
C6275 _0387_ _0776_/a_27_47# 0.04339f
C6276 _0217_ _0575_/a_109_297# 0.01063f
C6277 VPWR net247 1.70364f
C6278 hold42/a_49_47# net37 0.0163f
C6279 _0350_ _0611_/a_68_297# 0
C6280 _0642_/a_27_413# _0186_ 0
C6281 _1057_/a_466_413# net37 0
C6282 _0421_ net228 0.00142f
C6283 _0732_/a_80_21# acc0.A\[24\] 0.00994f
C6284 clknet_1_0__leaf__0459_ _0781_/a_68_297# 0.07147f
C6285 _0734_/a_47_47# _0362_ 0.15546f
C6286 _0269_ _0843_/a_150_297# 0
C6287 _0514_/a_27_297# net142 0
C6288 net150 net1 0.69915f
C6289 control0.state\[1\] comp0.B\[0\] 0.07494f
C6290 _0266_ _1014_/a_1059_315# 0
C6291 _0796_/a_79_21# _0796_/a_297_297# 0.01735f
C6292 _0591_/a_109_297# _0219_ 0
C6293 hold15/a_391_47# _1030_/a_1059_315# 0
C6294 acc0.A\[1\] _0345_ 0.07878f
C6295 _0195_ _0109_ 0
C6296 _0960_/a_27_47# _0960_/a_181_47# 0.00401f
C6297 _0305_ _0816_/a_68_297# 0
C6298 net119 control0.reset 0.03743f
C6299 hold24/a_391_47# VPWR 0.18115f
C6300 _0387_ _0219_ 0.00177f
C6301 _0608_/a_109_297# VPWR 0.00368f
C6302 hold42/a_391_47# net67 0.00704f
C6303 _0819_/a_299_297# acc0.A\[8\] 0
C6304 clkbuf_0__0465_/a_110_47# _0346_ 0.00196f
C6305 _0427_ _0659_/a_68_297# 0
C6306 _0982_/a_193_47# clknet_1_0__leaf__0461_ 0.00357f
C6307 net117 _0345_ 0.00788f
C6308 _1057_/a_891_413# net67 0.00341f
C6309 hold25/a_391_47# _0550_/a_51_297# 0
C6310 _0399_ hold70/a_285_47# 0
C6311 _0385_ _0462_ 0.02761f
C6312 _0983_/a_1017_47# _0455_ 0
C6313 VPWR _0825_/a_68_297# 0.15069f
C6314 net39 clknet_1_1__leaf__0459_ 0.59051f
C6315 clkbuf_0__0463_/a_110_47# _0563_/a_51_297# 0
C6316 acc0.A\[12\] acc0.A\[11\] 0.00243f
C6317 clkbuf_1_0__f__0460_/a_110_47# acc0.A\[24\] 0
C6318 _1063_/a_27_47# _0161_ 0.17171f
C6319 _1063_/a_1059_315# _1063_/a_1017_47# 0
C6320 VPWR _0844_/a_382_297# 0.00464f
C6321 net204 net171 0
C6322 _0968_/a_109_297# _1068_/a_27_47# 0
C6323 hold74/a_391_47# _0507_/a_27_297# 0
C6324 acc0.A\[20\] _1019_/a_193_47# 0
C6325 _0135_ _0173_ 0
C6326 acc0.A\[8\] _0437_ 0.02524f
C6327 hold100/a_285_47# net47 0
C6328 acc0.A\[1\] hold2/a_49_47# 0.05536f
C6329 _0250_ acc0.A\[24\] 0
C6330 VPWR _1024_/a_193_47# 0.30629f
C6331 _0188_ _0181_ 0.00888f
C6332 _0462_ _1006_/a_1017_47# 0
C6333 _0174_ _0535_/a_68_297# 0
C6334 _0121_ _0576_/a_373_47# 0
C6335 _1071_/a_193_47# _0976_/a_505_21# 0
C6336 _0982_/a_27_47# _0265_ 0
C6337 hold76/a_391_47# _0352_ 0
C6338 clknet_1_0__leaf__0464_ _1050_/a_1059_315# 0
C6339 net180 net31 0.00198f
C6340 _1049_/a_466_413# acc0.A\[15\] 0
C6341 _0748_/a_299_297# _0294_ 0.05955f
C6342 _0349_ _1012_/a_634_159# 0.00165f
C6343 VPWR _1048_/a_466_413# 0.25387f
C6344 net125 _0177_ 0.1621f
C6345 net232 _1062_/a_466_413# 0
C6346 _0343_ acc0.A\[15\] 0.2168f
C6347 _0855_/a_299_297# _0580_/a_27_297# 0
C6348 _0216_ clknet_1_0__leaf__0459_ 0.02914f
C6349 _1028_/a_561_413# clknet_1_1__leaf__0462_ 0
C6350 net204 net24 0
C6351 _1055_/a_634_159# net66 0
C6352 _1055_/a_193_47# acc0.A\[8\] 0
C6353 hold57/a_391_47# _0175_ 0
C6354 _0218_ _0186_ 0.01975f
C6355 _0273_ _0831_/a_35_297# 0.00119f
C6356 _0642_/a_215_297# _0253_ 0.02332f
C6357 hold47/a_49_47# hold47/a_285_47# 0.22264f
C6358 _0809_/a_81_21# net228 0.0108f
C6359 _0382_ _0219_ 0.0677f
C6360 clk _0958_/a_27_47# 0.00237f
C6361 _0355_ _0335_ 0
C6362 hold101/a_391_47# _0835_/a_215_47# 0
C6363 _0570_/a_373_47# acc0.A\[26\] 0
C6364 VPWR _1010_/a_561_413# 0.0031f
C6365 _1000_/a_27_47# _1000_/a_561_413# 0.0027f
C6366 _1000_/a_634_159# _1000_/a_891_413# 0.03684f
C6367 _1000_/a_193_47# _1000_/a_381_47# 0.09503f
C6368 _1033_/a_1059_315# clknet_1_0__leaf__0457_ 0
C6369 _1060_/a_27_47# _0158_ 0.07923f
C6370 _1060_/a_193_47# net146 0.00585f
C6371 _1060_/a_1059_315# _1060_/a_1017_47# 0
C6372 _1051_/a_634_159# net154 0.01634f
C6373 _0361_ _0319_ 0.00723f
C6374 _0513_/a_299_297# _0155_ 0.00152f
C6375 hold19/a_285_47# _0294_ 0
C6376 net114 _1008_/a_592_47# 0
C6377 _0187_ acc0.A\[10\] 0.12193f
C6378 _0168_ _0979_/a_109_297# 0
C6379 VPWR _0979_/a_373_47# 0
C6380 input32/a_75_212# B[9] 0.19816f
C6381 _1072_/a_193_47# VPWR 0.28648f
C6382 VPWR _0841_/a_79_21# 0.40984f
C6383 _1053_/a_975_413# net11 0
C6384 _0258_ clkbuf_1_0__f__0465_/a_110_47# 0.03203f
C6385 clknet_1_1__leaf__0458_ _0987_/a_634_159# 0
C6386 clkbuf_1_0__f__0458_/a_110_47# _0842_/a_59_75# 0.01108f
C6387 _0953_/a_32_297# comp0.B\[9\] 0.04627f
C6388 _0233_ _0742_/a_299_297# 0
C6389 _0320_ _0739_/a_297_297# 0
C6390 _0568_/a_373_47# acc0.A\[30\] 0
C6391 _0553_/a_149_47# _0136_ 0.02882f
C6392 _0399_ _0986_/a_381_47# 0.00364f
C6393 net105 hold60/a_285_47# 0.00335f
C6394 net207 hold60/a_49_47# 0
C6395 VPWR _1009_/a_975_413# 0.00487f
C6396 _0698_/a_199_47# _0317_ 0.01052f
C6397 acc0.A\[12\] hold81/a_391_47# 0.00206f
C6398 hold14/a_49_47# _0208_ 0.0018f
C6399 _0446_ _0265_ 0.00974f
C6400 net211 net187 0
C6401 net1 control0.add 0.01763f
C6402 _0457_ _1033_/a_634_159# 0
C6403 _0963_/a_35_297# _0963_/a_285_47# 0.00723f
C6404 _0346_ _0824_/a_59_75# 0.0533f
C6405 clknet_1_0__leaf__0458_ hold59/a_285_47# 0
C6406 _0401_ _0811_/a_384_47# 0
C6407 _0216_ _0453_ 0
C6408 _0655_/a_369_297# _0302_ 0
C6409 _0161_ _1062_/a_1059_315# 0.01421f
C6410 _0583_/a_109_47# net165 0
C6411 clknet_1_0__leaf__0462_ hold4/a_285_47# 0.01816f
C6412 _1071_/a_1017_47# VPWR 0
C6413 VPWR net100 0.71749f
C6414 _1056_/a_466_413# net178 0
C6415 _0998_/a_891_413# _0097_ 0
C6416 _0959_/a_80_21# _0160_ 0.15085f
C6417 _0476_ _1035_/a_27_47# 0
C6418 _0330_ _0701_/a_303_47# 0
C6419 _0216_ _0567_/a_373_47# 0
C6420 _0985_/a_381_47# _0179_ 0.0163f
C6421 _1055_/a_634_159# _0350_ 0
C6422 _0735_/a_109_297# _1010_/a_27_47# 0
C6423 net186 VPWR 0.30476f
C6424 net42 net5 0.01553f
C6425 clknet_1_1__leaf__0462_ _0739_/a_215_47# 0.00316f
C6426 net113 _0739_/a_79_21# 0
C6427 _0305_ clknet_0__0460_ 0
C6428 _0270_ _0261_ 0
C6429 acc0.A\[27\] acc0.A\[29\] 0
C6430 _0179_ _1049_/a_466_413# 0.0472f
C6431 clknet_1_1__leaf__0463_ _1065_/a_193_47# 0.0025f
C6432 clknet_1_1__leaf__0462_ _0352_ 0.00518f
C6433 _0707_/a_544_297# acc0.A\[29\] 0
C6434 _1059_/a_891_413# _0219_ 0.00211f
C6435 _0684_/a_145_75# _0328_ 0
C6436 _0778_/a_68_297# _0347_ 0
C6437 _0343_ _0179_ 0.02145f
C6438 _0459_ _0245_ 0
C6439 net64 _0437_ 0
C6440 net36 net8 0.42512f
C6441 _0499_/a_59_75# _0173_ 0
C6442 net157 net173 0
C6443 _0858_/a_27_47# _0261_ 0
C6444 hold25/a_49_47# net29 0
C6445 _0222_ _0754_/a_512_297# 0
C6446 clknet_0__0464_ _1046_/a_381_47# 0.02178f
C6447 _0997_/a_466_413# net41 0.03247f
C6448 _0997_/a_193_47# pp[14] 0
C6449 hold11/a_391_47# net157 0.04913f
C6450 _1071_/a_381_47# clkbuf_1_0__f_clk/a_110_47# 0.00145f
C6451 _1071_/a_466_413# clknet_0_clk 0.00397f
C6452 hold79/a_391_47# clk 0.0011f
C6453 net54 _1027_/a_381_47# 0.00674f
C6454 hold13/a_391_47# _0173_ 0.00197f
C6455 net185 net27 0.02032f
C6456 _0585_/a_109_47# _0208_ 0
C6457 _0473_ _0177_ 0
C6458 _0309_ clkbuf_1_1__f__0461_/a_110_47# 0
C6459 _0337_ _1030_/a_1059_315# 0
C6460 hold64/a_285_47# VPWR 0.2691f
C6461 net64 _1055_/a_193_47# 0
C6462 _0178_ _1047_/a_466_413# 0.00111f
C6463 _0538_/a_51_297# _1044_/a_27_47# 0
C6464 acc0.A\[27\] _0699_/a_68_297# 0
C6465 _1065_/a_27_47# _0468_ 0
C6466 _0577_/a_27_297# VPWR 0.25229f
C6467 _1055_/a_193_47# _0621_/a_117_297# 0
C6468 comp0.B\[11\] _1043_/a_381_47# 0
C6469 pp[29] acc0.A\[29\] 0.0244f
C6470 clkbuf_1_1__f__0465_/a_110_47# _0288_ 0
C6471 control0.state\[2\] _1066_/a_193_47# 0
C6472 net46 _0756_/a_47_47# 0.01003f
C6473 acc0.A\[14\] _1060_/a_27_47# 0.0057f
C6474 clknet_0__0459_ _0184_ 0
C6475 hold101/a_285_47# _0624_/a_59_75# 0
C6476 control0.state\[2\] _1068_/a_193_47# 0
C6477 _0486_ _1068_/a_27_47# 0.49098f
C6478 net21 _1045_/a_634_159# 0.01587f
C6479 _0201_ _1045_/a_891_413# 0.00494f
C6480 net183 _1045_/a_466_413# 0
C6481 clknet_1_0__leaf__0465_ net154 0.06899f
C6482 VPWR _1022_/a_592_47# 0
C6483 _0174_ _0208_ 0.0606f
C6484 _0852_/a_285_297# _0453_ 0.05532f
C6485 _0610_/a_145_75# acc0.A\[19\] 0
C6486 _0537_/a_68_297# _0202_ 0.0038f
C6487 _0978_/a_27_297# _0976_/a_76_199# 0
C6488 acc0.A\[17\] _0676_/a_113_47# 0
C6489 net214 _0401_ 0
C6490 _0999_/a_466_413# _0999_/a_561_413# 0.00772f
C6491 _0999_/a_634_159# _0999_/a_975_413# 0
C6492 _0854_/a_510_47# _0399_ 0.00153f
C6493 net17 _1063_/a_381_47# 0.01915f
C6494 _0295_ hold70/a_285_47# 0
C6495 _1001_/a_27_47# _1019_/a_634_159# 0.00638f
C6496 _1001_/a_193_47# _1019_/a_193_47# 0.00253f
C6497 _1017_/a_1059_315# _0115_ 0
C6498 _0772_/a_79_21# _0772_/a_215_47# 0.04584f
C6499 _0972_/a_584_47# clknet_1_1__leaf_clk 0
C6500 _1001_/a_381_47# net223 0
C6501 _1001_/a_891_413# _0391_ 0
C6502 _1001_/a_466_413# _0099_ 0.0035f
C6503 VPWR _0993_/a_193_47# 0.33357f
C6504 _1016_/a_27_47# _0582_/a_27_297# 0
C6505 clknet_1_1__leaf__0463_ net33 0
C6506 _1021_/a_27_47# net240 0
C6507 _0478_ control0.state\[2\] 0
C6508 net77 _0345_ 0
C6509 _1004_/a_1059_315# acc0.A\[22\] 0
C6510 _1004_/a_891_413# _0217_ 0
C6511 net1 net231 0
C6512 clknet_1_0__leaf__0462_ _1007_/a_193_47# 0.03933f
C6513 net43 clknet_1_1__leaf__0461_ 0.40639f
C6514 _1033_/a_634_159# _0475_ 0
C6515 net121 B[2] 0
C6516 _0534_/a_81_21# _0465_ 0.01354f
C6517 _0244_ _0611_/a_68_297# 0
C6518 net185 _0470_ 0
C6519 _0217_ _0171_ 0
C6520 pp[28] net208 0
C6521 _1020_/a_1059_315# net202 0
C6522 net115 clknet_1_1__leaf__0462_ 0.19606f
C6523 net57 _0725_/a_209_297# 0.00317f
C6524 _0223_ _0345_ 0
C6525 _0600_/a_253_47# _0219_ 0.00312f
C6526 _0232_ _0754_/a_240_47# 0
C6527 _1043_/a_27_47# _0542_/a_51_297# 0
C6528 _0642_/a_215_297# output61/a_27_47# 0
C6529 _0858_/a_27_47# _0509_/a_27_47# 0.00964f
C6530 B[7] _0207_ 0
C6531 _1021_/a_1059_315# _0119_ 0
C6532 _0961_/a_113_297# _0975_/a_59_75# 0
C6533 net135 net134 0.02205f
C6534 net242 _0352_ 0
C6535 _0999_/a_27_47# clknet_1_1__leaf__0461_ 0
C6536 _0732_/a_209_47# _0368_ 0.00297f
C6537 _0577_/a_27_297# net48 0.01196f
C6538 _0324_ hold90/a_49_47# 0.00935f
C6539 _0359_ hold90/a_285_47# 0.06011f
C6540 _0510_/a_109_297# _0187_ 0.00169f
C6541 _0510_/a_373_47# net4 0.00135f
C6542 clkbuf_1_1__f__0462_/a_110_47# net244 0
C6543 _1017_/a_193_47# _0218_ 0
C6544 _0733_/a_448_47# _0361_ 0
C6545 hold23/a_391_47# acc0.A\[2\] 0.00113f
C6546 _0200_ comp0.B\[10\] 0
C6547 _0481_ clk 0.01031f
C6548 acc0.A\[12\] _0303_ 0.33398f
C6549 hold86/a_285_47# _0850_/a_68_297# 0
C6550 _1043_/a_466_413# net20 0
C6551 net62 _0988_/a_1017_47# 0
C6552 _0160_ _0173_ 0
C6553 _0456_ _0448_ 0
C6554 _0782_/a_27_47# _0178_ 0
C6555 _1011_/a_891_413# _0219_ 0
C6556 net158 VPWR 0.35072f
C6557 net48 _1022_/a_592_47# 0
C6558 net126 _1041_/a_466_413# 0
C6559 _1006_/a_27_47# _0219_ 0
C6560 _0656_/a_59_75# _0345_ 0.00405f
C6561 net235 net47 0
C6562 hold12/a_285_47# _0468_ 0
C6563 output39/a_27_47# input5/a_75_212# 0.00124f
C6564 _0751_/a_111_297# net241 0
C6565 _0751_/a_29_53# _0219_ 0.01306f
C6566 _0216_ _0113_ 0.00275f
C6567 _0195_ _0128_ 0.01729f
C6568 _0241_ _0218_ 0.1698f
C6569 net150 _0225_ 0
C6570 clknet_1_0__leaf__0462_ _0328_ 0
C6571 _0183_ _0224_ 0
C6572 _0467_ _1068_/a_634_159# 0
C6573 _0614_/a_29_53# _0614_/a_111_297# 0.005f
C6574 _0461_ _0773_/a_117_297# 0
C6575 comp0.B\[10\] comp0.B\[8\] 0.5817f
C6576 _0985_/a_193_47# _0985_/a_634_159# 0.11897f
C6577 _0985_/a_27_47# _0985_/a_466_413# 0.27314f
C6578 net1 clknet_1_1__leaf__0457_ 0
C6579 comp0.B\[13\] _0535_/a_68_297# 0
C6580 hold85/a_391_47# net232 0.16486f
C6581 _0780_/a_35_297# _0397_ 0.17697f
C6582 _1018_/a_27_47# _1018_/a_193_47# 0.96163f
C6583 _0086_ _0831_/a_35_297# 0
C6584 _0833_/a_510_47# _0253_ 0
C6585 _0243_ hold64/a_391_47# 0
C6586 _0902_/a_27_47# _0369_ 0
C6587 control0.count\[2\] _1071_/a_381_47# 0.02077f
C6588 _0985_/a_27_47# _1049_/a_27_47# 0.00133f
C6589 _0535_/a_68_297# _1046_/a_193_47# 0
C6590 net50 _1022_/a_27_47# 0
C6591 _0642_/a_215_297# _0642_/a_382_47# 0.01048f
C6592 hold47/a_391_47# _1050_/a_1059_315# 0
C6593 hold47/a_285_47# _1050_/a_891_413# 0.01406f
C6594 acc0.A\[12\] _0281_ 0.29158f
C6595 _0275_ _0990_/a_27_47# 0.00134f
C6596 _0831_/a_117_297# _0271_ 0
C6597 _1050_/a_592_47# _0186_ 0.00106f
C6598 _0353_ _0707_/a_75_199# 0.02084f
C6599 _1010_/a_193_47# acc0.A\[29\] 0
C6600 _0267_ _0446_ 0.30937f
C6601 _0080_ _0262_ 0
C6602 net45 _0674_/a_113_47# 0
C6603 _0282_ _0650_/a_150_297# 0
C6604 _0582_/a_373_47# net219 0.0012f
C6605 _1019_/a_634_159# _0459_ 0
C6606 _0753_/a_297_297# _0753_/a_561_47# 0
C6607 _0254_ _0271_ 0.003f
C6608 hold55/a_391_47# clknet_1_0__leaf__0461_ 0.00148f
C6609 net11 net73 0.18587f
C6610 _0530_/a_81_21# _0530_/a_384_47# 0.00138f
C6611 comp0.B\[4\] net122 0.0015f
C6612 _0330_ hold50/a_49_47# 0
C6613 _0363_ acc0.A\[27\] 0
C6614 VPWR _0756_/a_377_297# 0.00667f
C6615 _0172_ _0548_/a_512_297# 0
C6616 _0734_/a_47_47# _0324_ 0
C6617 hold27/a_391_47# clkbuf_0__0464_/a_110_47# 0
C6618 net85 _0307_ 0.0023f
C6619 VPWR _1027_/a_891_413# 0.21261f
C6620 _0369_ _0673_/a_103_199# 0.00413f
C6621 _0586_/a_27_47# _0391_ 0
C6622 pp[7] _0619_/a_68_297# 0
C6623 net45 _0406_ 0
C6624 net56 _0704_/a_68_297# 0
C6625 _1003_/a_891_413# _0237_ 0.01489f
C6626 _0997_/a_193_47# _0408_ 0
C6627 _0805_/a_181_47# _0286_ 0
C6628 comp0.B\[13\] _0174_ 0.20059f
C6629 pp[27] net56 0.00704f
C6630 _0181_ clknet_0__0460_ 0
C6631 output39/a_27_47# pp[12] 0.16308f
C6632 _1056_/a_193_47# acc0.A\[10\] 0.01034f
C6633 net51 pp[23] 0.10517f
C6634 net109 _1005_/a_1059_315# 0
C6635 _1042_/a_466_413# hold51/a_285_47# 0
C6636 _1042_/a_634_159# hold51/a_391_47# 0
C6637 _0174_ _1046_/a_193_47# 0.01058f
C6638 net193 comp0.B\[10\] 0
C6639 _0677_/a_47_47# _0677_/a_285_47# 0.01755f
C6640 _0487_ _1063_/a_193_47# 0
C6641 _0546_/a_240_47# _1040_/a_466_413# 0
C6642 clkbuf_1_0__f__0459_/a_110_47# _0183_ 0.13028f
C6643 _0340_ _0219_ 0.03716f
C6644 _1019_/a_466_413# clknet_1_0__leaf__0461_ 0
C6645 _0584_/a_27_297# clkbuf_1_1__f__0457_/a_110_47# 0
C6646 _1004_/a_1059_315# _0379_ 0.03986f
C6647 clkbuf_0__0460_/a_110_47# _0743_/a_51_297# 0
C6648 _0252_ acc0.A\[8\] 1.07806f
C6649 _0188_ _0187_ 0
C6650 acc0.A\[8\] _0989_/a_381_47# 0.01974f
C6651 output67/a_27_47# _0512_/a_27_297# 0.00165f
C6652 _0346_ _0991_/a_1059_315# 0
C6653 clknet_1_0__leaf__0458_ _0219_ 0.03634f
C6654 net15 _0186_ 0.02665f
C6655 _0994_/a_634_159# net80 0
C6656 _0982_/a_193_47# _0218_ 0
C6657 hold78/a_49_47# _0341_ 0.05865f
C6658 _0487_ _0460_ 0.00587f
C6659 hold88/a_391_47# _0988_/a_891_413# 0.00206f
C6660 _0544_/a_51_297# net198 0.14583f
C6661 _0647_/a_47_47# _0403_ 0
C6662 hold64/a_285_47# clknet_1_0__leaf__0459_ 0
C6663 hold15/a_391_47# VPWR 0.19826f
C6664 _0272_ _0433_ 0
C6665 hold7/a_391_47# net73 0.00123f
C6666 hold7/a_285_47# _0085_ 0.01594f
C6667 net10 hold51/a_49_47# 0.01806f
C6668 net189 net37 0.00273f
C6669 _0730_/a_297_297# _0352_ 0
C6670 net68 _0509_/a_27_47# 0
C6671 _1058_/a_1059_315# net143 0.00915f
C6672 _0637_/a_56_297# _0263_ 0.06586f
C6673 _0637_/a_311_297# _0261_ 0
C6674 VPWR net148 0.76368f
C6675 _0189_ net142 0.00226f
C6676 _0650_/a_68_297# _0281_ 0
C6677 _1034_/a_634_159# _1034_/a_592_47# 0
C6678 _0536_/a_149_47# _0200_ 0.00154f
C6679 hold6/a_49_47# _0544_/a_240_47# 0
C6680 net219 clknet_1_0__leaf__0461_ 0
C6681 _0796_/a_215_47# _0094_ 0
C6682 VPWR rst 0.28956f
C6683 net162 _1030_/a_1017_47# 0
C6684 _0497_/a_68_297# _0177_ 0.10549f
C6685 _0310_ _0462_ 0
C6686 _0559_/a_149_47# net205 0.00831f
C6687 net168 _1053_/a_1017_47# 0
C6688 _0430_ _0434_ 1.0897f
C6689 _0251_ clknet_0__0465_ 0
C6690 hold25/a_391_47# _0172_ 0.00228f
C6691 hold25/a_49_47# _0137_ 0
C6692 net124 net28 0
C6693 _0729_/a_150_297# _0350_ 0
C6694 _0627_/a_215_53# VPWR 0.14046f
C6695 _0640_/a_109_53# clknet_0__0465_ 0.00379f
C6696 _0217_ _0456_ 0.05475f
C6697 _0259_ _0347_ 0
C6698 _0770_/a_297_47# control0.add 0.00714f
C6699 _1013_/a_381_47# _0219_ 0.00395f
C6700 hold36/a_285_47# comp0.B\[12\] 0
C6701 _0787_/a_80_21# _0807_/a_68_297# 0.01348f
C6702 control0.state\[0\] _1066_/a_561_413# 0
C6703 _0570_/a_27_297# net190 0.12602f
C6704 _0570_/a_109_47# net197 0
C6705 _1002_/a_1059_315# _0219_ 0
C6706 _0226_ _0460_ 0.04552f
C6707 _0963_/a_35_297# net226 0
C6708 _0086_ _0988_/a_381_47# 0.11277f
C6709 _0746_/a_81_21# _1006_/a_27_47# 0
C6710 acc0.A\[16\] _0219_ 0.4637f
C6711 control0.count\[3\] _0169_ 0
C6712 control0.state\[1\] _1068_/a_381_47# 0
C6713 control0.state\[1\] net1 0.03413f
C6714 _0129_ _0341_ 0
C6715 _0359_ clknet_0__0462_ 0.02351f
C6716 VPWR _1026_/a_975_413# 0.00482f
C6717 _0535_/a_68_297# comp0.B\[9\] 0
C6718 net63 _0253_ 0
C6719 _0848_/a_27_47# _0450_ 0.04679f
C6720 acc0.A\[22\] pp[19] 0
C6721 hold78/a_285_47# _1013_/a_1059_315# 0.00334f
C6722 _0344_ _1013_/a_27_47# 0
C6723 VPWR _0817_/a_266_297# 0.00295f
C6724 _0547_/a_150_297# _0206_ 0.00137f
C6725 _0218_ net62 0.27403f
C6726 _0793_/a_245_297# net42 0.00112f
C6727 net59 _1031_/a_27_47# 0
C6728 hold27/a_285_47# net147 0.03627f
C6729 _0218_ _0450_ 0.02728f
C6730 clkbuf_1_0__f__0459_/a_110_47# acc0.A\[15\] 0.01277f
C6731 _1058_/a_193_47# A[11] 0
C6732 net180 net7 0.13304f
C6733 _0517_/a_81_21# _0153_ 0.14476f
C6734 _0223_ net52 0
C6735 _1071_/a_634_159# _0488_ 0
C6736 _1071_/a_193_47# _0466_ 0.04024f
C6737 hold8/a_285_47# _0739_/a_79_21# 0
C6738 _0993_/a_27_47# _0286_ 0
C6739 _0993_/a_193_47# _0283_ 0
C6740 _0147_ acc0.A\[15\] 0
C6741 net81 _0995_/a_27_47# 0.22514f
C6742 acc0.A\[21\] net51 0.00406f
C6743 hold77/a_49_47# _1009_/a_27_47# 0
C6744 _1050_/a_27_47# _0987_/a_27_47# 0
C6745 net232 _0160_ 0.00947f
C6746 _1017_/a_1059_315# _1017_/a_891_413# 0.31086f
C6747 _1017_/a_193_47# _1017_/a_975_413# 0
C6748 _1017_/a_466_413# _1017_/a_381_47# 0.03733f
C6749 _0487_ _1062_/a_891_413# 0.05932f
C6750 _0348_ _0354_ 0
C6751 _0357_ _0727_/a_277_47# 0.00149f
C6752 net58 clknet_0__0465_ 0.09114f
C6753 net45 _0307_ 0.04504f
C6754 _0243_ _0766_/a_109_297# 0
C6755 _0343_ _0752_/a_27_413# 0
C6756 _0753_/a_381_47# _0234_ 0
C6757 _0753_/a_79_21# _0375_ 0.04295f
C6758 _1052_/a_466_413# net9 0.02234f
C6759 _0644_/a_377_297# _0346_ 0
C6760 net103 _1060_/a_1059_315# 0
C6761 clk _0477_ 0
C6762 _0473_ _1046_/a_1017_47# 0.00121f
C6763 _0472_ _1046_/a_975_413# 0
C6764 _0984_/a_1059_315# _0219_ 0.04742f
C6765 _1016_/a_193_47# _1060_/a_193_47# 0
C6766 _0463_ control0.reset 0
C6767 _0181_ net201 0
C6768 net178 _0088_ 0
C6769 net190 hold50/a_49_47# 0
C6770 net197 hold50/a_391_47# 0.12945f
C6771 _1006_/a_1059_315# net52 0.14466f
C6772 _1000_/a_193_47# net45 0.0413f
C6773 _0507_/a_109_297# acc0.A\[13\] 0.0015f
C6774 _1000_/a_891_413# net86 0
C6775 _1000_/a_1059_315# _0098_ 0
C6776 net64 _0252_ 0.335f
C6777 net137 net154 0
C6778 _0958_/a_197_47# _0161_ 0
C6779 _1051_/a_1017_47# net11 0
C6780 _0129_ _1013_/a_891_413# 0
C6781 hold54/a_285_47# net24 0
C6782 net163 _1013_/a_466_413# 0
C6783 _0363_ _1010_/a_193_47# 0.00125f
C6784 _0346_ _0425_ 0.16881f
C6785 _0303_ net42 0.198f
C6786 _0174_ comp0.B\[9\] 0.69371f
C6787 _0361_ _0250_ 0.00115f
C6788 _0804_/a_215_47# _0804_/a_510_47# 0.00529f
C6789 _0959_/a_217_297# _0477_ 0.00262f
C6790 _0452_ _0580_/a_27_297# 0
C6791 hold82/a_49_47# acc0.A\[13\] 0.29654f
C6792 clknet_1_1__leaf__0458_ net73 0.10085f
C6793 net204 _0553_/a_51_297# 0
C6794 clknet_0__0463_ _0171_ 0.02107f
C6795 _0704_/a_68_297# _0345_ 0.00372f
C6796 _0536_/a_240_47# _1046_/a_634_159# 0
C6797 _1033_/a_27_47# _1033_/a_466_413# 0.26036f
C6798 _1033_/a_193_47# _1033_/a_634_159# 0.12729f
C6799 pp[27] _0345_ 0.15466f
C6800 net55 _0734_/a_377_297# 0
C6801 _1012_/a_27_47# _1012_/a_466_413# 0.27314f
C6802 _1012_/a_193_47# _1012_/a_634_159# 0.12729f
C6803 _0292_ _0424_ 0.00439f
C6804 _0973_/a_373_47# _0161_ 0
C6805 hold23/a_49_47# _0509_/a_27_47# 0.00191f
C6806 _0195_ _0331_ 0.02984f
C6807 _0216_ net56 0.03756f
C6808 net221 _0347_ 0.03794f
C6809 _0197_ _1049_/a_27_47# 0
C6810 _0347_ _1007_/a_381_47# 0
C6811 _0352_ _1007_/a_466_413# 0
C6812 acc0.A\[12\] A[12] 0
C6813 _1056_/a_193_47# _0510_/a_109_297# 0
C6814 net9 _0194_ 0
C6815 _0216_ _1031_/a_634_159# 0
C6816 _0195_ _1031_/a_1059_315# 0
C6817 _0457_ net119 0.00371f
C6818 _0363_ _1009_/a_634_159# 0
C6819 _0274_ _0438_ 0
C6820 hold27/a_285_47# net125 0
C6821 _0343_ hold98/a_49_47# 0.00345f
C6822 clknet_1_0__leaf__0465_ clknet_0__0464_ 0.09052f
C6823 _0480_ clknet_0_clk 0
C6824 _1072_/a_891_413# clknet_0_clk 0.00525f
C6825 _1050_/a_634_159# _1050_/a_592_47# 0
C6826 _0257_ _0529_/a_27_297# 0
C6827 _0518_/a_27_297# _0987_/a_27_47# 0
C6828 _0720_/a_68_297# net209 0
C6829 _0343_ clkload3/a_110_47# 0
C6830 _0990_/a_634_159# _0181_ 0.00562f
C6831 _0717_/a_209_297# acc0.A\[29\] 0
C6832 pp[1] VPWR 0.58646f
C6833 _0443_ _0434_ 0
C6834 clkbuf_1_0__f__0459_/a_110_47# _0179_ 0
C6835 _1041_/a_634_159# _0546_/a_51_297# 0
C6836 _1024_/a_466_413# net50 0.00479f
C6837 clknet_1_0__leaf__0464_ _1051_/a_193_47# 0
C6838 clknet_1_1__leaf__0460_ _0397_ 0
C6839 net67 _0419_ 0
C6840 _0457_ clkbuf_0__0457_/a_110_47# 0.3114f
C6841 _0179_ _0147_ 0.73176f
C6842 hold29/a_391_47# _0122_ 0
C6843 VPWR _0837_/a_81_21# 0.60369f
C6844 _0465_ _0849_/a_510_47# 0
C6845 _1036_/a_1059_315# net28 0
C6846 hold24/a_49_47# comp0.B\[5\] 0
C6847 _0241_ _0099_ 0
C6848 _0180_ _0527_/a_109_297# 0.01373f
C6849 _0343_ clknet_1_1__leaf__0460_ 0.03804f
C6850 net61 _0267_ 0
C6851 clknet_1_0__leaf__0460_ _0616_/a_78_199# 0
C6852 _0337_ VPWR 0.57772f
C6853 _0662_/a_299_297# clknet_0__0465_ 0
C6854 _0259_ clkbuf_0__0465_/a_110_47# 0.00247f
C6855 _0615_/a_109_297# _0242_ 0.00152f
C6856 _0294_ _0246_ 0.23519f
C6857 _0598_/a_297_47# net51 0.0014f
C6858 _1054_/a_466_413# _1052_/a_891_413# 0
C6859 _0302_ _0300_ 0
C6860 clknet_1_1__leaf__0460_ net95 0.183f
C6861 _0409_ _0794_/a_27_47# 0.03303f
C6862 _0795_/a_81_21# _0277_ 0
C6863 _0982_/a_381_47# net149 0
C6864 _0176_ _1040_/a_1059_315# 0.03731f
C6865 _1014_/a_193_47# hold2/a_285_47# 0
C6866 _1014_/a_634_159# hold2/a_49_47# 0
C6867 _1014_/a_27_47# hold2/a_391_47# 0
C6868 net65 _0180_ 0.00339f
C6869 _0179_ _1054_/a_193_47# 0.09388f
C6870 _0178_ _0145_ 0.02622f
C6871 net141 _0621_/a_35_297# 0
C6872 net21 _1044_/a_193_47# 0.01868f
C6873 _0201_ _1044_/a_1059_315# 0
C6874 _0120_ VPWR 0.23315f
C6875 net83 _0345_ 0.04122f
C6876 _0788_/a_68_297# VPWR 0.19022f
C6877 _1056_/a_381_47# _0179_ 0.02776f
C6878 _1020_/a_1017_47# net187 0
C6879 _0833_/a_215_47# net62 0.00128f
C6880 _1001_/a_381_47# clkbuf_0__0457_/a_110_47# 0
C6881 _0995_/a_27_47# _0797_/a_207_413# 0
C6882 _0995_/a_193_47# _0797_/a_27_413# 0
C6883 net21 net131 0
C6884 net183 net184 0
C6885 net84 net42 0.00103f
C6886 net205 _1036_/a_634_159# 0
C6887 clknet_1_0__leaf__0461_ _0352_ 0
C6888 _0973_/a_109_297# net240 0.02967f
C6889 _0555_/a_240_47# _0173_ 0.01676f
C6890 _0555_/a_245_297# _0208_ 0.00151f
C6891 _1024_/a_193_47# _1023_/a_27_47# 0
C6892 _1024_/a_27_47# _1023_/a_193_47# 0
C6893 comp0.B\[13\] _1046_/a_193_47# 0
C6894 comp0.B\[2\] _0181_ 0
C6895 _0592_/a_68_297# net109 0
C6896 pp[1] output62/a_27_47# 0.04597f
C6897 _0180_ _0935_/a_27_47# 0
C6898 _0533_/a_373_47# _0465_ 0
C6899 _0781_/a_68_297# _0345_ 0
C6900 _0432_ _0346_ 0.17553f
C6901 acc0.A\[15\] _0842_/a_59_75# 0
C6902 _1054_/a_27_47# net75 0
C6903 _0817_/a_585_47# clknet_1_1__leaf__0465_ 0
C6904 _0180_ _1061_/a_193_47# 0
C6905 net8 _1061_/a_27_47# 0
C6906 _0343_ _1000_/a_1017_47# 0
C6907 hold67/a_391_47# _0292_ 0
C6908 _0293_ _0275_ 0.00933f
C6909 _0465_ hold71/a_391_47# 0.01562f
C6910 _1012_/a_27_47# net98 0.22685f
C6911 _0178_ net17 0
C6912 _1012_/a_634_159# clknet_1_1__leaf__0461_ 0
C6913 _1046_/a_27_47# _1046_/a_634_159# 0.13601f
C6914 hold86/a_391_47# hold100/a_49_47# 0
C6915 hold86/a_49_47# hold100/a_391_47# 0
C6916 hold86/a_285_47# hold100/a_285_47# 0.00245f
C6917 _0978_/a_27_297# _0488_ 0.09085f
C6918 hold55/a_49_47# _0208_ 0
C6919 net55 clknet_0__0462_ 0
C6920 clknet_1_0__leaf__0462_ output51/a_27_47# 0.00139f
C6921 _0219_ net91 0
C6922 net241 _0103_ 0
C6923 _0772_/a_510_47# _0099_ 0
C6924 net61 _0642_/a_215_297# 0
C6925 _1056_/a_27_47# _0517_/a_81_21# 0
C6926 net231 control0.sh 0.00343f
C6927 _1016_/a_891_413# net221 0.02614f
C6928 _1016_/a_27_47# _0115_ 0.03143f
C6929 _1032_/a_27_47# clknet_1_0__leaf__0457_ 0.00437f
C6930 _0432_ net65 0
C6931 _0752_/a_384_47# _0375_ 0
C6932 _0752_/a_27_413# _0376_ 0.15167f
C6933 acc0.A\[2\] hold71/a_391_47# 0
C6934 output56/a_27_47# _0219_ 0
C6935 _0322_ _0360_ 0.00275f
C6936 net23 comp0.B\[15\] 0.00525f
C6937 _0131_ _0472_ 0.00775f
C6938 _0664_/a_79_21# _0422_ 0
C6939 _0724_/a_199_47# _0345_ 0
C6940 VPWR _0542_/a_240_47# 0.00597f
C6941 _0983_/a_975_413# _0183_ 0
C6942 _0775_/a_79_21# _0393_ 0.15509f
C6943 output66/a_27_47# _0189_ 0.00324f
C6944 _0260_ _0255_ 0.0049f
C6945 _0327_ _0360_ 0
C6946 _0996_/a_193_47# acc0.A\[15\] 0.01168f
C6947 _1043_/a_193_47# net19 0.00106f
C6948 _0211_ _1036_/a_193_47# 0
C6949 clknet_0__0458_ hold75/a_49_47# 0
C6950 hold38/a_49_47# _0175_ 0.06744f
C6951 acc0.A\[12\] _1057_/a_193_47# 0.00776f
C6952 hold27/a_285_47# _0473_ 0.0139f
C6953 _1001_/a_975_413# net206 0
C6954 _0467_ _0564_/a_68_297# 0
C6955 net63 _0518_/a_109_297# 0
C6956 _0539_/a_68_297# _0176_ 0.11014f
C6957 _1019_/a_193_47# _0208_ 0
C6958 net44 _0999_/a_193_47# 0.0042f
C6959 _0120_ net48 0.01431f
C6960 _1030_/a_1059_315# _0333_ 0
C6961 _0206_ net153 0
C6962 clknet_1_1__leaf__0459_ _0999_/a_1059_315# 0
C6963 _0229_ _0750_/a_27_47# 0.09271f
C6964 hold34/a_49_47# VPWR 0.25013f
C6965 hold23/a_285_47# clknet_1_0__leaf__0464_ 0.00214f
C6966 net103 _0294_ 0
C6967 _1000_/a_27_47# net46 0
C6968 acc0.A\[3\] clknet_1_1__leaf__0457_ 0
C6969 VPWR _0406_ 0.24754f
C6970 net196 net20 0.04189f
C6971 _1052_/a_634_159# _0522_/a_27_297# 0
C6972 _1052_/a_193_47# _0522_/a_109_297# 0
C6973 hold26/a_285_47# net7 0
C6974 _0216_ _0345_ 0.75671f
C6975 _0401_ _0421_ 0
C6976 _0467_ clknet_1_1__leaf_clk 0.16959f
C6977 _0731_/a_81_21# _0318_ 0
C6978 _0259_ _0824_/a_59_75# 0
C6979 _0092_ _0218_ 0.0244f
C6980 _0598_/a_79_21# acc0.A\[21\] 0.00135f
C6981 control0.sh clknet_1_1__leaf__0457_ 0
C6982 _0518_/a_27_297# _0191_ 0.14973f
C6983 _1039_/a_27_47# net8 0.08057f
C6984 hold41/a_285_47# VPWR 0.27389f
C6985 hold100/a_391_47# acc0.A\[14\] 0
C6986 _0712_/a_561_47# _0195_ 0
C6987 _0985_/a_1059_315# _0985_/a_1017_47# 0
C6988 _0985_/a_27_47# _0083_ 0.09744f
C6989 net116 net209 0.00104f
C6990 acc0.A\[10\] clknet_1_1__leaf__0465_ 0.15497f
C6991 net186 comp0.B\[3\] 0
C6992 acc0.A\[22\] net176 0.00272f
C6993 comp0.B\[0\] _0564_/a_68_297# 0.17078f
C6994 _1018_/a_466_413# _1018_/a_592_47# 0.00553f
C6995 _1018_/a_634_159# _1018_/a_1017_47# 0
C6996 net136 _0218_ 0
C6997 net36 _1014_/a_891_413# 0
C6998 _0300_ net6 0.09586f
C6999 hold19/a_285_47# _1016_/a_466_413# 0.00145f
C7000 comp0.B\[14\] _1046_/a_381_47# 0
C7001 _0404_ _0302_ 0
C7002 hold21/a_49_47# clknet_1_1__leaf__0458_ 0
C7003 _0789_/a_201_297# _0409_ 0.03134f
C7004 _0404_ _0795_/a_299_297# 0
C7005 _0298_ _0795_/a_81_21# 0
C7006 hold47/a_49_47# acc0.A\[4\] 0
C7007 _0716_/a_27_47# hold81/a_49_47# 0
C7008 net36 _0492_/a_27_47# 0.04165f
C7009 _0982_/a_466_413# _0982_/a_381_47# 0.03733f
C7010 _0982_/a_193_47# _0982_/a_975_413# 0
C7011 _0982_/a_1059_315# _0982_/a_891_413# 0.31086f
C7012 _0222_ acc0.A\[23\] 0
C7013 _1011_/a_466_413# clknet_1_1__leaf__0462_ 0
C7014 _1049_/a_634_159# _1049_/a_381_47# 0
C7015 _0983_/a_975_413# acc0.A\[15\] 0
C7016 _0869_/a_27_47# _0350_ 0.01197f
C7017 clknet_1_1__leaf_clk comp0.B\[0\] 0.17582f
C7018 net12 _0522_/a_109_297# 0.00923f
C7019 net105 _0459_ 0.00168f
C7020 pp[10] input3/a_75_212# 0
C7021 _0343_ _0233_ 0.05162f
C7022 VPWR _0319_ 0.54346f
C7023 _0462_ _0315_ 0.0499f
C7024 _0399_ _0841_/a_215_47# 0.00506f
C7025 _1053_/a_27_47# _1053_/a_193_47# 0.97453f
C7026 _0760_/a_47_47# _0460_ 0.00124f
C7027 _0172_ _0138_ 0.74723f
C7028 _0276_ _0301_ 0.04169f
C7029 acc0.A\[1\] _0634_/a_113_47# 0
C7030 _1019_/a_466_413# _0218_ 0
C7031 hold98/a_391_47# net245 0.1316f
C7032 comp0.B\[13\] comp0.B\[9\] 0.002f
C7033 net204 _0135_ 0
C7034 _0195_ _1008_/a_27_47# 0
C7035 net203 net23 0
C7036 hold16/a_391_47# _0195_ 0.00343f
C7037 _1066_/a_634_159# _1066_/a_381_47# 0
C7038 clknet_0__0459_ hold74/a_391_47# 0
C7039 acc0.A\[14\] _0094_ 0
C7040 _0849_/a_79_21# _0263_ 0.00308f
C7041 net1 _1066_/a_634_159# 0
C7042 _0101_ _0382_ 0
C7043 net45 _0999_/a_975_413# 0
C7044 pp[9] A[11] 0.42175f
C7045 net9 net195 0
C7046 _0401_ _0809_/a_81_21# 0
C7047 _1068_/a_634_159# _1068_/a_381_47# 0
C7048 _0346_ hold70/a_285_47# 0.00151f
C7049 _0290_ _0809_/a_299_297# 0
C7050 _1030_/a_27_47# _1030_/a_466_413# 0.26957f
C7051 _1030_/a_193_47# _1030_/a_634_159# 0.11897f
C7052 _0449_ _0843_/a_68_297# 0.01196f
C7053 acc0.A\[22\] hold68/a_49_47# 0
C7054 _0217_ hold68/a_285_47# 0.0333f
C7055 _0557_/a_240_47# comp0.B\[4\] 0.00576f
C7056 net71 _0844_/a_297_47# 0
C7057 _0402_ _0807_/a_68_297# 0.00104f
C7058 _1017_/a_27_47# _0347_ 0
C7059 _0218_ net219 0.14078f
C7060 net207 clknet_1_0__leaf__0461_ 0.0481f
C7061 _0299_ net81 0
C7062 net187 _0461_ 0.00609f
C7063 net157 clknet_1_1__leaf__0457_ 0.09245f
C7064 net205 comp0.B\[5\] 0
C7065 net150 _0462_ 0
C7066 _0752_/a_27_413# _0224_ 0.00167f
C7067 _0476_ _0959_/a_80_21# 0.02639f
C7068 _0251_ _0519_/a_81_21# 0
C7069 _0416_ _0279_ 0.0934f
C7070 _0415_ _0278_ 0
C7071 _0174_ hold5/a_285_47# 0
C7072 _0312_ _1009_/a_466_413# 0
C7073 _0313_ net113 0.0024f
C7074 net148 _0523_/a_81_21# 0.06287f
C7075 _1035_/a_466_413# clknet_1_1__leaf__0463_ 0.00489f
C7076 _1035_/a_193_47# net122 0
C7077 _0992_/a_1059_315# hold70/a_49_47# 0.00923f
C7078 _0992_/a_634_159# hold70/a_391_47# 0.00982f
C7079 _0992_/a_466_413# hold70/a_285_47# 0.01371f
C7080 control0.count\[1\] _0975_/a_59_75# 0
C7081 VPWR control0.state\[2\] 2.05474f
C7082 _0195_ _0611_/a_68_297# 0
C7083 hold53/a_49_47# net200 0.00106f
C7084 hold53/a_391_47# _0123_ 0
C7085 _0598_/a_79_21# _0598_/a_297_47# 0.03259f
C7086 net120 VPWR 0.33375f
C7087 _0204_ _0140_ 0
C7088 _1015_/a_193_47# _0181_ 0.02459f
C7089 _0183_ net87 0.49457f
C7090 net71 _1048_/a_1059_315# 0
C7091 VPWR _0307_ 0.35838f
C7092 _0238_ _0748_/a_81_21# 0
C7093 _0222_ _0602_/a_113_47# 0
C7094 hold47/a_49_47# _1051_/a_466_413# 0
C7095 _1034_/a_891_413# comp0.B\[2\] 0.04217f
C7096 hold6/a_391_47# _0140_ 0.0014f
C7097 net247 _0345_ 0.00119f
C7098 _0533_/a_27_297# _1047_/a_27_47# 0
C7099 pp[7] net65 0.06208f
C7100 _0254_ net76 0
C7101 _0125_ _1008_/a_193_47# 0
C7102 acc0.A\[27\] _1008_/a_1059_315# 0
C7103 _0992_/a_193_47# net67 0.00141f
C7104 _1000_/a_193_47# VPWR 0.28319f
C7105 _0326_ clkbuf_1_0__f__0462_/a_110_47# 0
C7106 net24 _0562_/a_68_297# 0
C7107 VPWR _0513_/a_384_47# 0
C7108 _0796_/a_79_21# net41 0.00358f
C7109 _0983_/a_1059_315# _0181_ 0.02268f
C7110 clknet_0__0464_ _1044_/a_466_413# 0
C7111 _1072_/a_466_413# _0466_ 0.00113f
C7112 net137 clknet_0__0464_ 0
C7113 acc0.A\[14\] _0508_/a_299_297# 0
C7114 hold89/a_49_47# clk 0.00625f
C7115 _0404_ net6 0.06334f
C7116 _0219_ _0505_/a_109_297# 0.05088f
C7117 control0.state\[1\] control0.sh 0
C7118 net190 _0126_ 0.16554f
C7119 B[12] input21/a_75_212# 0.00253f
C7120 input20/a_75_212# B[13] 0.00556f
C7121 _0346_ _1006_/a_381_47# 0.01173f
C7122 net46 _0374_ 0.00327f
C7123 _0756_/a_285_47# net50 0.0503f
C7124 hold2/a_49_47# net247 0
C7125 acc0.A\[12\] _0803_/a_68_297# 0
C7126 hold52/a_285_47# _0216_ 0
C7127 net176 _0379_ 0
C7128 net168 hold21/a_391_47# 0.13574f
C7129 pp[30] _1031_/a_592_47# 0
C7130 _0227_ _0606_/a_109_53# 0
C7131 _1032_/a_891_413# clknet_1_0__leaf__0461_ 0.00291f
C7132 _0686_/a_219_297# _0364_ 0
C7133 net175 _0530_/a_299_297# 0.05953f
C7134 net104 _0242_ 0
C7135 net83 _0791_/a_113_297# 0.00144f
C7136 _0343_ _0998_/a_466_413# 0.00205f
C7137 _0581_/a_27_297# _0393_ 0
C7138 _1008_/a_1059_315# _0364_ 0.02163f
C7139 _0815_/a_113_297# net47 0
C7140 _0218_ _0637_/a_56_297# 0.00581f
C7141 _0645_/a_285_47# _0996_/a_27_47# 0
C7142 clknet_1_0__leaf__0465_ _0536_/a_51_297# 0.00485f
C7143 acc0.A\[12\] _0672_/a_215_47# 0.00485f
C7144 clknet_1_0__leaf__0463_ _0550_/a_51_297# 0.08085f
C7145 _1017_/a_193_47# _1016_/a_1059_315# 0.00808f
C7146 _1017_/a_27_47# _1016_/a_891_413# 0.00309f
C7147 _1017_/a_466_413# _1016_/a_634_159# 0
C7148 hold55/a_285_47# _0178_ 0
C7149 _0520_/a_27_297# _0180_ 0.11937f
C7150 _0661_/a_27_297# _0661_/a_277_297# 0.00876f
C7151 net178 _0516_/a_109_297# 0
C7152 _0233_ _0376_ 0.00161f
C7153 _0509_/a_27_47# hold71/a_49_47# 0
C7154 acc0.A\[8\] _0988_/a_891_413# 0
C7155 _0268_ _0186_ 0
C7156 _0402_ net217 0
C7157 _0998_/a_634_159# acc0.A\[17\] 0
C7158 _0310_ _0312_ 0
C7159 _0681_/a_113_47# VPWR 0
C7160 input25/a_75_212# net25 0.10849f
C7161 _0578_/a_109_297# acc0.A\[20\] 0
C7162 _0643_/a_103_199# _0255_ 0.00335f
C7163 _0216_ net52 0.14495f
C7164 VPWR B[11] 0.21667f
C7165 _1037_/a_27_47# clknet_1_1__leaf__0463_ 0.00163f
C7166 _0465_ _0986_/a_193_47# 0
C7167 _0998_/a_27_47# clkbuf_1_1__f__0461_/a_110_47# 0.01732f
C7168 _0555_/a_51_297# _0555_/a_512_297# 0.0116f
C7169 _0533_/a_27_297# clknet_1_0__leaf__0461_ 0
C7170 _0462_ control0.add 0.0698f
C7171 _0733_/a_448_47# VPWR 0.00307f
C7172 _1067_/a_27_47# _1065_/a_1059_315# 0
C7173 _0399_ _0790_/a_35_297# 0.0019f
C7174 net58 _0986_/a_27_47# 0.03741f
C7175 pp[28] _0221_ 0.04333f
C7176 _0299_ _0797_/a_207_413# 0.21357f
C7177 _0298_ _0797_/a_297_47# 0
C7178 _0476_ _0173_ 0.05682f
C7179 hold47/a_285_47# clknet_1_0__leaf__0465_ 0.00644f
C7180 _0308_ _1009_/a_27_47# 0
C7181 _1033_/a_27_47# _0131_ 0.08937f
C7182 _1033_/a_193_47# net119 0.00727f
C7183 _1033_/a_1059_315# _1033_/a_1017_47# 0
C7184 _0192_ net230 0.1903f
C7185 net234 acc0.A\[19\] 0
C7186 _0248_ _0617_/a_150_297# 0
C7187 _0372_ _0617_/a_68_297# 0
C7188 hold87/a_391_47# _0261_ 0
C7189 hold87/a_285_47# _0263_ 0
C7190 _0083_ _0197_ 0
C7191 net63 _0987_/a_193_47# 0.00489f
C7192 _0841_/a_79_21# _0345_ 0.06431f
C7193 hold68/a_49_47# _0379_ 0
C7194 _1012_/a_1059_315# _1012_/a_1017_47# 0
C7195 VPWR _0780_/a_285_297# 0.25434f
C7196 _0130_ _1033_/a_634_159# 0
C7197 _0148_ net154 0
C7198 _0196_ net11 0.00393f
C7199 net64 pp[8] 0.00196f
C7200 _0693_/a_68_297# _0368_ 0
C7201 pp[9] net66 0.00294f
C7202 _0545_/a_150_297# _0202_ 0
C7203 _0343_ clknet_1_1__leaf__0459_ 0.25989f
C7204 _0529_/a_109_297# _0261_ 0.00588f
C7205 _0529_/a_109_47# _0262_ 0
C7206 net226 _0484_ 0.00385f
C7207 _0352_ _0105_ 0
C7208 _0102_ net93 0
C7209 net3 _0186_ 0.00274f
C7210 _1056_/a_634_159# _0187_ 0
C7211 acc0.A\[20\] net202 0
C7212 _0172_ net134 0
C7213 net46 acc0.A\[19\] 0.43852f
C7214 _0753_/a_79_21# VPWR 0.18668f
C7215 _0719_/a_27_47# _0350_ 0.18773f
C7216 _1054_/a_27_47# hold83/a_285_47# 0
C7217 _1009_/a_1059_315# _0219_ 0.04102f
C7218 hold86/a_285_47# net233 0.01507f
C7219 _0964_/a_109_297# _0481_ 0
C7220 _0460_ _0350_ 0.05791f
C7221 _0269_ _0265_ 0
C7222 net44 _0677_/a_285_47# 0.06726f
C7223 _1050_/a_891_413# acc0.A\[4\] 0.04689f
C7224 _0459_ hold72/a_49_47# 0.01075f
C7225 _0729_/a_68_297# _0334_ 0.00159f
C7226 net106 clknet_1_0__leaf__0461_ 0.19048f
C7227 _0343_ _1030_/a_975_413# 0
C7228 net35 _0382_ 0
C7229 _1055_/a_381_47# acc0.A\[9\] 0
C7230 _0854_/a_79_21# _0853_/a_68_297# 0
C7231 _1041_/a_1059_315# net152 0.00115f
C7232 hold100/a_285_47# _0458_ 0
C7233 net100 _0345_ 0
C7234 _0854_/a_510_47# _0346_ 0
C7235 _0122_ net50 0.09964f
C7236 _0625_/a_59_75# clknet_1_0__leaf__0465_ 0.00178f
C7237 _0946_/a_30_53# _0485_ 0.02481f
C7238 _0446_ _0347_ 0
C7239 _0794_/a_326_47# acc0.A\[15\] 0
C7240 _0244_ _0869_/a_27_47# 0
C7241 _0836_/a_150_297# _0369_ 0
C7242 _0993_/a_27_47# net79 0.22616f
C7243 net158 hold26/a_391_47# 0
C7244 VPWR _0544_/a_512_297# 0.00628f
C7245 _0358_ _0350_ 0.03417f
C7246 net231 _0955_/a_32_297# 0
C7247 _0983_/a_193_47# _1018_/a_466_413# 0
C7248 hold96/a_49_47# pp[24] 0
C7249 hold96/a_391_47# net52 0.00235f
C7250 control0.state\[1\] _0483_ 0
C7251 net149 _0116_ 0
C7252 _0218_ _0352_ 0.42246f
C7253 VPWR _1034_/a_466_413# 0.24086f
C7254 clknet_1_0__leaf__0460_ _1067_/a_193_47# 0.00361f
C7255 _0179_ _1057_/a_27_47# 0
C7256 net198 _1043_/a_27_47# 0.02767f
C7257 _0129_ acc0.A\[30\] 0
C7258 _0369_ _0437_ 0.09296f
C7259 _0383_ clknet_1_0__leaf__0460_ 0
C7260 net169 _1052_/a_891_413# 0
C7261 _0188_ clknet_1_1__leaf__0465_ 0.01512f
C7262 _0465_ _0845_/a_109_47# 0.0024f
C7263 _0531_/a_27_297# _0531_/a_109_297# 0.17136f
C7264 comp0.B\[7\] net36 0.44526f
C7265 _0996_/a_27_47# _0507_/a_27_297# 0
C7266 net61 net63 0.02021f
C7267 hold6/a_285_47# _1043_/a_466_413# 0
C7268 _1053_/a_1059_315# input12/a_75_212# 0
C7269 _1053_/a_193_47# A[5] 0
C7270 net87 hold40/a_285_47# 0
C7271 net46 _0249_ 0.20857f
C7272 _1002_/a_27_47# acc0.A\[20\] 0
C7273 _0998_/a_27_47# _0998_/a_1059_315# 0.04875f
C7274 _0998_/a_193_47# _0998_/a_466_413# 0.07593f
C7275 hold32/a_285_47# VPWR 0.31946f
C7276 _0956_/a_220_297# _0208_ 0.00371f
C7277 clknet_1_0__leaf__0458_ net58 0.02268f
C7278 net64 _0988_/a_891_413# 0.03009f
C7279 _1059_/a_634_159# _0459_ 0.00802f
C7280 _0498_/a_51_297# _0935_/a_27_47# 0.07709f
C7281 hold64/a_285_47# _0345_ 0.00586f
C7282 _1031_/a_592_47# _0339_ 0.0015f
C7283 _0343_ _0292_ 0
C7284 _1003_/a_27_47# _0369_ 0
C7285 _0498_/a_51_297# _1061_/a_193_47# 0
C7286 _0410_ _0792_/a_80_21# 0
C7287 net85 _0998_/a_891_413# 0.00124f
C7288 clknet_1_0__leaf__0459_ _0307_ 0
C7289 _0662_/a_299_297# _0986_/a_27_47# 0
C7290 _0662_/a_81_21# _0986_/a_193_47# 0
C7291 net193 _1046_/a_1017_47# 0
C7292 hold87/a_285_47# clknet_1_0__leaf__0461_ 0.00258f
C7293 hold38/a_285_47# _0955_/a_32_297# 0
C7294 _0960_/a_27_47# clkbuf_1_0__f_clk/a_110_47# 0.00874f
C7295 VPWR _0507_/a_109_297# 0.19727f
C7296 _1019_/a_27_47# _1019_/a_634_159# 0.13601f
C7297 net44 _1012_/a_466_413# 0
C7298 _1046_/a_891_413# _1046_/a_975_413# 0.00851f
C7299 _1046_/a_27_47# net132 0.2197f
C7300 _1046_/a_381_47# _1046_/a_561_413# 0.00123f
C7301 _1019_/a_466_413# _0099_ 0.00327f
C7302 _0227_ hold3/a_285_47# 0
C7303 acc0.A\[21\] hold3/a_391_47# 0.07402f
C7304 _1000_/a_193_47# clknet_1_0__leaf__0459_ 0
C7305 _0809_/a_81_21# hold70/a_49_47# 0
C7306 pp[26] net197 0
C7307 net54 net190 0.02638f
C7308 _1056_/a_466_413# _0153_ 0
C7309 net133 _0533_/a_27_297# 0
C7310 net123 input29/a_75_212# 0.00167f
C7311 control0.state\[1\] control0.count\[1\] 0
C7312 VPWR hold82/a_49_47# 0.30903f
C7313 net154 _0525_/a_384_47# 0.00928f
C7314 net215 net110 0
C7315 _1039_/a_891_413# clkbuf_1_0__f__0463_/a_110_47# 0.00712f
C7316 _0783_/a_79_21# _0307_ 0.02503f
C7317 _0565_/a_51_297# _0175_ 0
C7318 _0957_/a_32_297# _0176_ 0.12707f
C7319 clknet_1_0__leaf__0462_ _0123_ 0.03067f
C7320 clknet_1_0__leaf_clk _0468_ 0.13151f
C7321 _0266_ _0181_ 0.11114f
C7322 net175 _1049_/a_1059_315# 0.00565f
C7323 net9 _1049_/a_193_47# 0.01486f
C7324 hold34/a_391_47# A[9] 0
C7325 output64/a_27_47# net62 0
C7326 _0343_ _0435_ 0.2345f
C7327 hold87/a_391_47# net47 0.00785f
C7328 VPWR _0333_ 0.72892f
C7329 pp[2] pp[3] 0.1811f
C7330 _0275_ _0840_/a_150_297# 0
C7331 _0259_ _0425_ 0
C7332 hold32/a_285_47# output62/a_27_47# 0
C7333 net160 comp0.B\[5\] 0.09811f
C7334 comp0.B\[1\] net17 0.19925f
C7335 _0775_/a_215_47# _0352_ 0.05702f
C7336 _0457_ _1032_/a_592_47# 0
C7337 _0220_ net209 0
C7338 net34 clkbuf_1_0__f_clk/a_110_47# 0
C7339 hold76/a_49_47# _0247_ 0.0039f
C7340 pp[30] net163 0.00465f
C7341 _0278_ _0347_ 0
C7342 clknet_1_0__leaf__0465_ comp0.B\[14\] 0.00766f
C7343 _0857_/a_27_47# clknet_1_1__leaf__0463_ 0.03769f
C7344 acc0.A\[1\] clknet_1_0__leaf__0457_ 0
C7345 _1056_/a_975_413# _0189_ 0
C7346 hold88/a_49_47# hold88/a_285_47# 0.22264f
C7347 _0758_/a_79_21# _0758_/a_510_47# 0.00844f
C7348 _0758_/a_297_297# _0758_/a_215_47# 0
C7349 _1024_/a_1059_315# output52/a_27_47# 0.00635f
C7350 _1024_/a_193_47# net52 0.01223f
C7351 VPWR _0999_/a_975_413# 0.00491f
C7352 _1052_/a_634_159# _0193_ 0
C7353 _1052_/a_561_413# acc0.A\[6\] 0.00141f
C7354 _0984_/a_891_413# _0465_ 0
C7355 _0581_/a_27_297# net206 0.09768f
C7356 _0581_/a_109_47# net219 0
C7357 _0990_/a_27_47# _0990_/a_466_413# 0.26005f
C7358 _0990_/a_193_47# _0990_/a_634_159# 0.11897f
C7359 clkbuf_0__0463_/a_110_47# _0173_ 0.01079f
C7360 _0245_ _0347_ 0.0239f
C7361 _0732_/a_80_21# VPWR 0.1488f
C7362 _0287_ acc0.A\[13\] 0.00273f
C7363 _0179_ acc0.A\[6\] 0.12156f
C7364 _1002_/a_27_47# _0880_/a_27_47# 0
C7365 _0534_/a_384_47# net149 0.00912f
C7366 net168 _0519_/a_81_21# 0.09688f
C7367 _0260_ _0843_/a_68_297# 0.17389f
C7368 _0733_/a_222_93# clkbuf_0__0462_/a_110_47# 0.01227f
C7369 _0326_ net51 0
C7370 _0464_ _0142_ 0.00343f
C7371 hold7/a_285_47# _0525_/a_81_21# 0
C7372 _0984_/a_1059_315# net58 0.08733f
C7373 hold27/a_285_47# comp0.B\[8\] 0.01018f
C7374 _0264_ _0261_ 0
C7375 VPWR net4 0.35966f
C7376 net8 _0953_/a_32_297# 0
C7377 _0348_ _0353_ 0
C7378 net232 _0476_ 0.28009f
C7379 _0672_/a_215_47# net42 0.0059f
C7380 net203 _0213_ 0
C7381 hold19/a_285_47# net166 0.01139f
C7382 _0985_/a_891_413# acc0.A\[3\] 0
C7383 _0463_ _0475_ 0
C7384 hold56/a_285_47# _0132_ 0
C7385 _0346_ _1014_/a_1059_315# 0.02758f
C7386 acc0.A\[25\] _1007_/a_27_47# 0
C7387 _0967_/a_215_297# _0484_ 0
C7388 _0967_/a_109_93# _0485_ 0
C7389 _0485_ _0487_ 0.00827f
C7390 net44 net98 0
C7391 _0343_ _0793_/a_512_297# 0
C7392 pp[2] _0273_ 0.00118f
C7393 _1053_/a_381_47# _0191_ 0
C7394 _0982_/a_381_47# _0080_ 0.12808f
C7395 VPWR hold83/a_391_47# 0.17613f
C7396 clknet_1_1__leaf__0463_ _1062_/a_27_47# 0
C7397 hold88/a_49_47# _0086_ 0
C7398 _1049_/a_891_413# _0147_ 0.03819f
C7399 _1049_/a_634_159# acc0.A\[3\] 0
C7400 _1049_/a_381_47# net135 0
C7401 VPWR net118 0.72327f
C7402 clknet_1_1__leaf__0459_ net38 0.00478f
C7403 _0552_/a_68_297# _0175_ 0
C7404 VPWR clkbuf_1_0__f__0460_/a_110_47# 1.45197f
C7405 hold25/a_391_47# _1040_/a_193_47# 0
C7406 hold25/a_49_47# _1040_/a_466_413# 0
C7407 _0459_ clknet_0__0461_ 0.04507f
C7408 _1011_/a_193_47# hold80/a_391_47# 0
C7409 _0818_/a_109_47# acc0.A\[9\] 0
C7410 hold9/a_285_47# _0347_ 0
C7411 net57 _0703_/a_109_297# 0.00176f
C7412 _0747_/a_297_297# _0104_ 0
C7413 _0226_ _0373_ 1.07503f
C7414 _0747_/a_510_47# _0371_ 0.00122f
C7415 _0838_/a_109_297# VPWR 0.00442f
C7416 net248 _0989_/a_193_47# 0
C7417 VPWR _0250_ 1.02737f
C7418 acc0.A\[1\] _0635_/a_27_47# 0
C7419 _0949_/a_59_75# _1062_/a_891_413# 0
C7420 _1070_/a_634_159# _1070_/a_381_47# 0
C7421 _1052_/a_193_47# _0150_ 0.53509f
C7422 _1053_/a_466_413# _1053_/a_592_47# 0.00553f
C7423 _1053_/a_634_159# _1053_/a_1017_47# 0
C7424 hold98/a_391_47# VPWR 0.18458f
C7425 _0575_/a_373_47# net199 0.00122f
C7426 net44 _1030_/a_466_413# 0.02625f
C7427 pp[17] _1030_/a_193_47# 0
C7428 _1057_/a_381_47# acc0.A\[10\] 0.00825f
C7429 _0269_ _0267_ 0
C7430 clknet_1_0__leaf__0463_ _0913_/a_27_47# 0.00681f
C7431 net207 _0218_ 0
C7432 clknet_1_0__leaf__0465_ _1050_/a_381_47# 0
C7433 _0532_/a_384_47# _0465_ 0
C7434 hold77/a_49_47# _0685_/a_68_297# 0
C7435 _0960_/a_27_47# control0.count\[2\] 0.21532f
C7436 net45 _0998_/a_891_413# 0.00598f
C7437 acc0.A\[22\] _1023_/a_466_413# 0.00324f
C7438 _0120_ _1023_/a_27_47# 0
C7439 _0217_ _1023_/a_1059_315# 0
C7440 _0816_/a_68_297# clknet_1_1__leaf__0465_ 0.0046f
C7441 _0198_ _1061_/a_466_413# 0
C7442 _1032_/a_466_413# _0208_ 0
C7443 hold43/a_285_47# _0216_ 0.03837f
C7444 _1066_/a_634_159# control0.sh 0.00493f
C7445 _1066_/a_381_47# clknet_1_1__leaf_clk 0
C7446 _0217_ hold59/a_285_47# 0.06949f
C7447 clknet_1_1__leaf__0463_ _0561_/a_51_297# 0.00559f
C7448 _0314_ _1007_/a_381_47# 0
C7449 _0559_/a_51_297# _1034_/a_1059_315# 0.00862f
C7450 _0261_ net170 0.04751f
C7451 net1 clknet_1_1__leaf_clk 0
C7452 _0502_/a_27_47# _0500_/a_27_47# 0.01996f
C7453 _1061_/a_27_47# _0492_/a_27_47# 0
C7454 net109 _1022_/a_561_413# 0
C7455 _1068_/a_891_413# _0166_ 0
C7456 _0259_ _0432_ 0
C7457 _1030_/a_1059_315# _1030_/a_1017_47# 0
C7458 _0997_/a_193_47# net83 0.00347f
C7459 _1038_/a_1059_315# _0552_/a_68_297# 0.00179f
C7460 hold78/a_391_47# _0339_ 0.00964f
C7461 hold63/a_285_47# hold53/a_285_47# 0.00306f
C7462 _0747_/a_79_21# _0745_/a_193_47# 0
C7463 clkbuf_1_1__f__0465_/a_110_47# _0424_ 0
C7464 clknet_1_0__leaf__0458_ _0262_ 0.01585f
C7465 _0272_ _0399_ 0
C7466 clknet_0__0463_ _0494_/a_27_47# 0.00242f
C7467 clknet_1_0__leaf__0462_ _0758_/a_510_47# 0
C7468 _0330_ net227 0
C7469 hold27/a_285_47# _1046_/a_466_413# 0
C7470 input4/a_75_212# net4 0.11027f
C7471 _1014_/a_891_413# hold60/a_391_47# 0.00206f
C7472 _0430_ _0186_ 0.02257f
C7473 net12 _0150_ 0.02951f
C7474 hold100/a_49_47# _0268_ 0
C7475 acc0.A\[14\] _0637_/a_139_47# 0.0012f
C7476 acc0.A\[27\] clknet_1_1__leaf__0462_ 0.15807f
C7477 _0133_ clknet_1_1__leaf__0463_ 0.07696f
C7478 _0231_ net46 0.03351f
C7479 _1056_/a_27_47# _1056_/a_466_413# 0.27314f
C7480 _1056_/a_193_47# _1056_/a_634_159# 0.11072f
C7481 _1032_/a_634_159# net17 0.00971f
C7482 _0143_ net10 0
C7483 _0243_ _0242_ 0.02233f
C7484 _0294_ _0815_/a_113_297# 0
C7485 _0458_ _0270_ 0
C7486 net34 control0.count\[2\] 0
C7487 _0229_ _0230_ 0.00318f
C7488 hold28/a_49_47# hold71/a_285_47# 0
C7489 _0987_/a_634_159# _0987_/a_592_47# 0
C7490 _0312_ _0315_ 0
C7491 _0305_ _0399_ 0.02124f
C7492 acc0.A\[5\] _0186_ 0.00565f
C7493 clknet_1_1__leaf__0459_ hold81/a_285_47# 0.01456f
C7494 _0218_ _0613_/a_109_297# 0.00362f
C7495 _0855_/a_299_297# _0855_/a_384_47# 0
C7496 _0558_/a_68_297# clknet_1_1__leaf__0463_ 0.00194f
C7497 acc0.A\[1\] _1047_/a_891_413# 0.00676f
C7498 _1052_/a_381_47# input14/a_75_212# 0
C7499 _0180_ _1047_/a_466_413# 0
C7500 _0182_ _1047_/a_1059_315# 0
C7501 _0199_ _1047_/a_27_47# 0.03358f
C7502 _0858_/a_27_47# _0458_ 0.11032f
C7503 hold15/a_391_47# _0345_ 0
C7504 clknet_0_clk _0163_ 0.00193f
C7505 output54/a_27_47# net54 0.1765f
C7506 _1004_/a_634_159# _1004_/a_381_47# 0
C7507 _0218_ _0849_/a_79_21# 0.00495f
C7508 _0195_ _0729_/a_150_297# 0
C7509 net163 _0339_ 0.09068f
C7510 clknet_1_0__leaf__0459_ _0507_/a_109_297# 0
C7511 _1027_/a_27_47# _1008_/a_466_413# 0
C7512 pp[16] _0340_ 0
C7513 _0557_/a_240_47# _1035_/a_193_47# 0
C7514 _0557_/a_51_297# _1035_/a_891_413# 0
C7515 net157 _1049_/a_634_159# 0
C7516 acc0.A\[30\] hold61/a_285_47# 0.08394f
C7517 _0953_/a_32_297# net10 0
C7518 _1021_/a_891_413# _0382_ 0
C7519 hold18/a_285_47# _0465_ 0.0181f
C7520 output66/a_27_47# net67 0
C7521 hold23/a_285_47# clkbuf_1_0__f__0464_/a_110_47# 0.00254f
C7522 _1067_/a_27_47# hold93/a_49_47# 0
C7523 net170 _0509_/a_27_47# 0
C7524 _0337_ net56 0.00349f
C7525 _0369_ hold93/a_285_47# 0
C7526 net47 _0264_ 0.27312f
C7527 acc0.A\[1\] _0850_/a_68_297# 0.1882f
C7528 clknet_1_1__leaf__0462_ _0364_ 0.0032f
C7529 _0447_ _0843_/a_150_297# 0
C7530 _0172_ net22 0.23585f
C7531 clknet_1_0__leaf__0465_ _1053_/a_193_47# 0.00236f
C7532 net82 clkbuf_0__0459_/a_110_47# 0.01357f
C7533 _1039_/a_27_47# _0492_/a_27_47# 0
C7534 _1029_/a_634_159# _1029_/a_592_47# 0
C7535 acc0.A\[16\] _0582_/a_109_297# 0
C7536 net58 hold18/a_49_47# 0
C7537 _0583_/a_27_297# net102 0
C7538 _0503_/a_109_297# VPWR 0.00677f
C7539 _0352_ _0099_ 0.09483f
C7540 _0577_/a_109_297# clknet_1_0__leaf__0460_ 0
C7541 clknet_0__0464_ _0148_ 0
C7542 comp0.B\[11\] hold51/a_391_47# 0
C7543 _0448_ _0219_ 0.02329f
C7544 net62 _0268_ 0
C7545 _0999_/a_1059_315# _0095_ 0
C7546 _0268_ _0450_ 0.28165f
C7547 _0328_ _0737_/a_35_297# 0.01728f
C7548 _0817_/a_266_297# _0345_ 0.00121f
C7549 _0116_ _0393_ 0.0011f
C7550 clknet_1_1__leaf__0463_ net107 0
C7551 _0110_ clknet_1_1__leaf__0462_ 0.00151f
C7552 _0462_ _0610_/a_145_75# 0
C7553 hold67/a_391_47# clkbuf_1_1__f__0465_/a_110_47# 0
C7554 comp0.B\[13\] _1045_/a_1017_47# 0.00191f
C7555 hold66/a_285_47# _0377_ 0
C7556 acc0.A\[4\] _0987_/a_891_413# 0.01088f
C7557 _0961_/a_113_297# _0479_ 0.14117f
C7558 _1015_/a_27_47# net201 0
C7559 _0716_/a_27_47# _0286_ 0.00468f
C7560 net233 _0458_ 0.00166f
C7561 _1020_/a_27_47# _0217_ 0.00104f
C7562 _1020_/a_193_47# net150 0
C7563 clknet_1_0__leaf__0463_ _0172_ 0.35752f
C7564 _0359_ _0352_ 0
C7565 _0182_ _0186_ 0.01102f
C7566 net103 _1016_/a_466_413# 0.00923f
C7567 _0661_/a_277_297# _0293_ 0
C7568 _0398_ net43 0.12921f
C7569 _0381_ net51 0
C7570 _1016_/a_27_47# _1016_/a_193_47# 0.96163f
C7571 net84 acc0.A\[17\] 0
C7572 input2/a_75_212# net2 0.10968f
C7573 hold13/a_49_47# _0496_/a_27_47# 0.00125f
C7574 _0856_/a_215_47# _0465_ 0.00177f
C7575 acc0.A\[27\] net242 0
C7576 control0.count\[3\] _1068_/a_1059_315# 0
C7577 _0483_ _1068_/a_634_159# 0.00187f
C7578 clknet_1_1__leaf__0460_ hold69/a_49_47# 0.00792f
C7579 _0101_ net91 0
C7580 net243 acc0.A\[23\] 0.02916f
C7581 _1028_/a_466_413# _1028_/a_561_413# 0.00772f
C7582 _1028_/a_634_159# _1028_/a_975_413# 0
C7583 _0555_/a_240_47# net204 0.05177f
C7584 net188 hold42/a_49_47# 0.03843f
C7585 _0343_ _0996_/a_466_413# 0.00193f
C7586 acc0.A\[2\] _0856_/a_215_47# 0
C7587 _0252_ _0369_ 0.03736f
C7588 hold31/a_49_47# _0989_/a_27_47# 0
C7589 _0369_ _0989_/a_381_47# 0.00435f
C7590 _0812_/a_79_21# _0812_/a_215_47# 0.04584f
C7591 _0765_/a_215_47# clknet_1_0__leaf__0457_ 0
C7592 _0765_/a_79_21# _0460_ 0.02492f
C7593 _0999_/a_27_47# _0398_ 0
C7594 _0306_ _1009_/a_1017_47# 0
C7595 _1033_/a_975_413# comp0.B\[1\] 0
C7596 _0369_ _0992_/a_381_47# 0
C7597 _0553_/a_240_47# _0176_ 0.00336f
C7598 clknet_1_1__leaf__0459_ _0282_ 0.02234f
C7599 VPWR _1018_/a_592_47# 0
C7600 _0130_ net119 0
C7601 hold55/a_285_47# comp0.B\[1\] 0
C7602 _0351_ _0720_/a_150_297# 0
C7603 clknet_1_1__leaf__0460_ _0109_ 0
C7604 _0693_/a_68_297# clknet_0__0460_ 0
C7605 net230 clknet_1_0__leaf__0465_ 0.02419f
C7606 VPWR _1049_/a_561_413# 0.00292f
C7607 _0581_/a_27_297# _0774_/a_150_297# 0
C7608 _0538_/a_51_297# _0540_/a_51_297# 0
C7609 net200 _0352_ 0
C7610 _0516_/a_27_297# _0181_ 0.17518f
C7611 _0812_/a_510_47# net228 0
C7612 _0647_/a_47_47# VPWR 0.38193f
C7613 _0575_/a_373_47# VPWR 0
C7614 _1041_/a_891_413# net31 0.06825f
C7615 pp[15] _0797_/a_297_47# 0
C7616 _0460_ _1006_/a_634_159# 0.0102f
C7617 hold97/a_49_47# _1008_/a_891_413# 0.00386f
C7618 hold97/a_285_47# _1008_/a_1059_315# 0.00108f
C7619 hold97/a_391_47# _1008_/a_466_413# 0.00388f
C7620 VPWR _1066_/a_561_413# 0.00579f
C7621 _0751_/a_183_297# _0460_ 0
C7622 net120 comp0.B\[3\] 0
C7623 net167 _1072_/a_27_47# 0
C7624 _1010_/a_193_47# clknet_1_1__leaf__0462_ 0
C7625 net235 clkbuf_1_1__f__0458_/a_110_47# 0
C7626 hold37/a_49_47# clknet_1_0__leaf__0465_ 0.00676f
C7627 VPWR _1068_/a_561_413# 0.00213f
C7628 clkload0/a_27_47# _0217_ 0
C7629 _0218_ hold72/a_285_47# 0.09382f
C7630 _0241_ clkbuf_1_0__f__0461_/a_110_47# 0.02269f
C7631 _0367_ _0219_ 0.00586f
C7632 _0387_ _0775_/a_79_21# 0.00135f
C7633 hold14/a_49_47# clknet_1_1__leaf__0463_ 0.00956f
C7634 _0229_ _0236_ 0
C7635 _0993_/a_466_413# _0091_ 0.0019f
C7636 VPWR _0140_ 0.39093f
C7637 _0175_ _0493_/a_27_47# 0.08932f
C7638 hold87/a_285_47# _0848_/a_27_47# 0
C7639 _0661_/a_205_297# clknet_1_1__leaf__0465_ 0
C7640 net213 _0228_ 0.00329f
C7641 _0769_/a_299_297# _0218_ 0
C7642 _0204_ net129 0
C7643 _0107_ _0305_ 0
C7644 clknet_1_0__leaf__0465_ _1046_/a_561_413# 0
C7645 _1018_/a_27_47# _0612_/a_59_75# 0.00388f
C7646 hold87/a_285_47# _0218_ 0
C7647 _0697_/a_80_21# _0319_ 0.05198f
C7648 _0343_ _0983_/a_1017_47# 0.00115f
C7649 _0531_/a_373_47# net9 0.00164f
C7650 _0433_ _0438_ 0
C7651 _0767_/a_59_75# _0246_ 0
C7652 hold57/a_49_47# _1039_/a_27_47# 0
C7653 _0996_/a_634_159# net5 0.03486f
C7654 _0996_/a_891_413# acc0.A\[13\] 0
C7655 _0996_/a_27_47# _0185_ 0
C7656 _0680_/a_80_21# _0219_ 0
C7657 _0136_ _0463_ 0.0013f
C7658 _0337_ _0345_ 0
C7659 clknet_0_clk _1068_/a_27_47# 0.03194f
C7660 net56 _0319_ 0.00211f
C7661 VPWR _0834_/a_109_297# 0.00618f
C7662 _1019_/a_381_47# clkbuf_0__0457_/a_110_47# 0.00126f
C7663 _0998_/a_891_413# _0998_/a_1017_47# 0.00617f
C7664 _0998_/a_634_159# net84 0.00639f
C7665 net45 _0793_/a_240_47# 0
C7666 comp0.B\[2\] _1015_/a_27_47# 0
C7667 net211 hold40/a_49_47# 0.00632f
C7668 acc0.A\[12\] _0511_/a_81_21# 0
C7669 _0804_/a_215_47# net80 0
C7670 _1020_/a_193_47# control0.add 0
C7671 _0305_ _0295_ 0
C7672 clknet_1_0__leaf__0460_ _0756_/a_129_47# 0
C7673 acc0.A\[11\] _0281_ 0.03344f
C7674 _0396_ _0308_ 0
C7675 _0961_/a_199_47# VPWR 0
C7676 net247 _1061_/a_466_413# 0
C7677 _0217_ _0219_ 0
C7678 _1024_/a_381_47# acc0.A\[23\] 0
C7679 net203 _1033_/a_466_413# 0.00228f
C7680 _0399_ _0181_ 0.18911f
C7681 _0788_/a_68_297# _0345_ 0.00296f
C7682 _0551_/a_27_47# _0112_ 0
C7683 _0984_/a_466_413# net47 0.01243f
C7684 net31 net147 0
C7685 net190 _0569_/a_109_297# 0.0015f
C7686 _0968_/a_193_297# net236 0.00125f
C7687 net34 _0966_/a_27_47# 0
C7688 hold38/a_285_47# _0474_ 0.00245f
C7689 _0176_ _0213_ 0.01431f
C7690 _1019_/a_891_413# _1019_/a_975_413# 0.00851f
C7691 _1019_/a_27_47# net105 0.27741f
C7692 _1019_/a_381_47# _1019_/a_561_413# 0.00123f
C7693 _0714_/a_51_297# _0714_/a_149_47# 0.02487f
C7694 clknet_1_0__leaf__0462_ hold63/a_49_47# 0
C7695 _0123_ _0574_/a_373_47# 0
C7696 _0965_/a_47_47# _0965_/a_285_47# 0.01755f
C7697 hold42/a_49_47# _0155_ 0.36572f
C7698 clknet_1_1__leaf__0463_ _0959_/a_300_47# 0
C7699 _0442_ _0172_ 0.2052f
C7700 net133 _0199_ 0
C7701 VPWR _1012_/a_1017_47# 0
C7702 comp0.B\[7\] _1061_/a_27_47# 0
C7703 _0149_ _1050_/a_891_413# 0.00437f
C7704 net201 _0215_ 0.01506f
C7705 hold83/a_49_47# acc0.A\[6\] 0.29541f
C7706 _0548_/a_51_297# net174 0.06964f
C7707 _0183_ hold2/a_391_47# 0.00137f
C7708 hold24/a_391_47# net171 0.15815f
C7709 hold24/a_285_47# _0207_ 0.01856f
C7710 _0575_/a_27_297# net176 0
C7711 _1033_/a_891_413# _1032_/a_891_413# 0.00333f
C7712 _0600_/a_103_199# net51 0.03297f
C7713 net242 _1010_/a_193_47# 0
C7714 net67 _0420_ 0
C7715 _0316_ _0739_/a_297_297# 0
C7716 _1013_/a_466_413# _0220_ 0
C7717 hold5/a_49_47# hold5/a_391_47# 0.00188f
C7718 _0326_ _0324_ 0.42351f
C7719 net55 _0352_ 0.0237f
C7720 _0337_ hold16/a_49_47# 0
C7721 hold58/a_49_47# _1035_/a_1059_315# 0.00435f
C7722 _0655_/a_215_53# hold81/a_285_47# 0
C7723 _0982_/a_1059_315# _0350_ 0.0237f
C7724 _0902_/a_27_47# acc0.A\[19\] 0
C7725 VPWR _0998_/a_891_413# 0.19426f
C7726 _0716_/a_27_47# _0672_/a_79_21# 0.01138f
C7727 acc0.A\[29\] hold50/a_285_47# 0
C7728 clknet_1_0__leaf__0465_ _0987_/a_381_47# 0.00315f
C7729 _0212_ _0176_ 0.00651f
C7730 hold3/a_285_47# _0352_ 0
C7731 _0347_ _0739_/a_297_297# 0
C7732 _0990_/a_634_159# clknet_1_1__leaf__0465_ 0
C7733 _0465_ _1048_/a_27_47# 0.0047f
C7734 clknet_0__0458_ _0434_ 0.0652f
C7735 _0294_ _0991_/a_975_413# 0
C7736 hold23/a_49_47# _0458_ 0.00133f
C7737 _0176_ _0547_/a_68_297# 0.10432f
C7738 net206 _0116_ 0.06464f
C7739 _0990_/a_27_47# _0088_ 0.09751f
C7740 _0990_/a_1059_315# _0990_/a_1017_47# 0
C7741 _0357_ _0334_ 0
C7742 _0244_ _0614_/a_29_53# 0.12613f
C7743 hold81/a_391_47# _0281_ 0
C7744 hold81/a_49_47# _0418_ 0
C7745 _0546_/a_149_47# net127 0
C7746 _0406_ _0345_ 0.03161f
C7747 _0267_ _0082_ 0
C7748 _1002_/a_381_47# _0460_ 0.00591f
C7749 _0218_ _0392_ 0
C7750 net46 _0225_ 0.23829f
C7751 _1032_/a_634_159# _0165_ 0
C7752 acc0.A\[2\] _1048_/a_27_47# 0.00387f
C7753 _0174_ net8 0.0244f
C7754 _0793_/a_51_297# _0793_/a_512_297# 0.0116f
C7755 _0343_ _0617_/a_150_297# 0
C7756 _0366_ acc0.A\[23\] 0
C7757 pp[30] _0720_/a_68_297# 0
C7758 output59/a_27_47# net239 0
C7759 output46/a_27_47# hold29/a_285_47# 0
C7760 net42 _0669_/a_29_53# 0
C7761 _1050_/a_193_47# _0180_ 0.03744f
C7762 _0174_ net32 0.24316f
C7763 hold35/a_285_47# _0153_ 0
C7764 _0743_/a_51_297# _0368_ 0.09199f
C7765 _0967_/a_297_297# _0476_ 0.01809f
C7766 _0770_/a_297_47# net46 0.00295f
C7767 _0260_ _0257_ 0.00158f
C7768 _0343_ _0095_ 0.0093f
C7769 clknet_1_0__leaf__0460_ net110 0
C7770 comp0.B\[7\] _1039_/a_27_47# 0
C7771 _0110_ hold92/a_49_47# 0
C7772 output42/a_27_47# net42 0.16607f
C7773 _0123_ _1025_/a_891_413# 0.01133f
C7774 net200 _1025_/a_466_413# 0.02568f
C7775 _0195_ _0869_/a_27_47# 0
C7776 net135 acc0.A\[3\] 0
C7777 clkload4/a_268_47# _0369_ 0.00105f
C7778 _0183_ _0611_/a_68_297# 0.00398f
C7779 _1034_/a_27_47# comp0.B\[6\] 0.02302f
C7780 _1034_/a_193_47# comp0.B\[5\] 0
C7781 _0465_ _0846_/a_512_297# 0
C7782 _0743_/a_149_47# _0319_ 0
C7783 hold25/a_49_47# net174 0
C7784 _1051_/a_634_159# _1051_/a_466_413# 0.23992f
C7785 _1051_/a_193_47# _1051_/a_1059_315# 0.03405f
C7786 _1051_/a_27_47# _1051_/a_891_413# 0.03224f
C7787 hold9/a_285_47# _0106_ 0.00137f
C7788 _0451_ _0350_ 0.3953f
C7789 _1056_/a_634_159# clknet_1_1__leaf__0465_ 0
C7790 _0742_/a_299_297# _0219_ 0.00244f
C7791 input20/a_75_212# net128 0
C7792 acc0.A\[14\] _0849_/a_215_47# 0.04862f
C7793 hold100/a_49_47# net222 0
C7794 net106 _1033_/a_891_413# 0
C7795 _1070_/a_891_413# _0168_ 0
C7796 _1070_/a_634_159# control0.count\[1\] 0.00167f
C7797 _1045_/a_1059_315# _1045_/a_891_413# 0.31086f
C7798 _1045_/a_193_47# _1045_/a_975_413# 0
C7799 _1045_/a_466_413# _1045_/a_381_47# 0.03733f
C7800 _1070_/a_561_413# VPWR 0.00579f
C7801 _0811_/a_81_21# acc0.A\[10\] 0
C7802 _0113_ net118 0
C7803 hold90/a_49_47# _0360_ 0.05271f
C7804 clknet_1_0__leaf__0465_ acc0.A\[4\] 0.04846f
C7805 _0680_/a_80_21# _0746_/a_81_21# 0
C7806 _1003_/a_27_47# hold66/a_391_47# 0
C7807 _0584_/a_27_297# _0566_/a_27_47# 0.00118f
C7808 _0319_ _0345_ 0.05292f
C7809 clknet_1_0__leaf__0462_ _0121_ 0.0405f
C7810 net202 _0208_ 0.01109f
C7811 _0678_/a_150_297# _0306_ 0
C7812 _0183_ net109 0.03053f
C7813 acc0.A\[22\] net177 0.13376f
C7814 VPWR _1043_/a_634_159# 0.18505f
C7815 hold21/a_49_47# net15 0
C7816 clknet_1_1__leaf_clk control0.sh 0
C7817 _0209_ input29/a_75_212# 0
C7818 hold23/a_391_47# acc0.A\[4\] 0
C7819 VPWR _1030_/a_1017_47# 0
C7820 clknet_1_1__leaf__0463_ _0208_ 0.11145f
C7821 _1029_/a_193_47# _0106_ 0
C7822 _0733_/a_448_47# _0697_/a_80_21# 0.00123f
C7823 _1043_/a_1059_315# _1043_/a_891_413# 0.31086f
C7824 _1043_/a_193_47# _1043_/a_975_413# 0
C7825 _1043_/a_466_413# _1043_/a_381_47# 0.03733f
C7826 _1018_/a_27_47# _0399_ 0.00977f
C7827 _0636_/a_59_75# _0636_/a_145_75# 0.00658f
C7828 _0848_/a_109_297# _0264_ 0
C7829 comp0.B\[2\] _0215_ 0.00136f
C7830 hold46/a_285_47# _0176_ 0.00454f
C7831 _0535_/a_68_297# net10 0.05739f
C7832 _0430_ net62 0
C7833 _0574_/a_27_297# _0347_ 0
C7834 _0248_ _0219_ 0
C7835 clknet_1_1__leaf__0459_ _0654_/a_297_47# 0.0012f
C7836 _0784_/a_113_47# _0410_ 0
C7837 _1038_/a_975_413# _0209_ 0
C7838 _0263_ _0449_ 0
C7839 _1030_/a_27_47# net208 0
C7840 clknet_1_1__leaf__0460_ _0777_/a_377_297# 0
C7841 _1004_/a_561_413# VPWR 0.00368f
C7842 _1021_/a_1059_315# _1002_/a_891_413# 0.01065f
C7843 _1021_/a_891_413# _1002_/a_1059_315# 0.00358f
C7844 VPWR input9/a_27_47# 0.26943f
C7845 _0518_/a_109_297# _0180_ 0.01148f
C7846 _1054_/a_27_47# _1054_/a_1059_315# 0.04875f
C7847 _1054_/a_193_47# _1054_/a_466_413# 0.07443f
C7848 _0775_/a_215_47# _0392_ 0.05954f
C7849 clkbuf_0__0459_/a_110_47# net146 0
C7850 _1071_/a_466_413# clknet_1_0__leaf_clk 0
C7851 _1015_/a_27_47# _1015_/a_193_47# 0.96639f
C7852 _0401_ net62 0.00504f
C7853 _0107_ _0181_ 0.30971f
C7854 hold100/a_285_47# acc0.A\[1\] 0
C7855 _0983_/a_193_47# VPWR 0.29433f
C7856 _0174_ _1042_/a_1059_315# 0.03193f
C7857 _0454_ _0261_ 0
C7858 _0730_/a_215_47# _1010_/a_27_47# 0
C7859 _0730_/a_79_21# _1010_/a_634_159# 0
C7860 net8 _0208_ 0.00192f
C7861 _0982_/a_634_159# acc0.A\[1\] 0
C7862 acc0.A\[20\] _0771_/a_27_413# 0
C7863 _0987_/a_975_413# _0085_ 0
C7864 _0792_/a_209_297# _0792_/a_303_47# 0
C7865 _0195_ _0633_/a_109_297# 0
C7866 net36 _0117_ 0
C7867 _0689_/a_68_297# _0686_/a_219_297# 0
C7868 _1038_/a_27_47# _1038_/a_634_159# 0.14145f
C7869 _0556_/a_68_297# _1037_/a_27_47# 0.00357f
C7870 _0287_ VPWR 0.64441f
C7871 hold88/a_285_47# net76 0
C7872 _0984_/a_193_47# _0267_ 0
C7873 net222 _0450_ 0
C7874 _0180_ _0145_ 0.0084f
C7875 A[12] acc0.A\[11\] 0.04663f
C7876 _0145_ net218 0
C7877 _0856_/a_79_21# net47 0.01243f
C7878 _1041_/a_27_47# net173 0
C7879 _0174_ net10 0.02376f
C7880 _0972_/a_346_47# _0471_ 0.00373f
C7881 acc0.A\[8\] _0987_/a_1059_315# 0
C7882 _0557_/a_512_297# _0133_ 0
C7883 _0727_/a_277_47# _0356_ 0.01045f
C7884 net157 net135 0
C7885 pp[29] hold80/a_49_47# 0.03852f
C7886 hold78/a_285_47# net162 0
C7887 _0515_/a_81_21# acc0.A\[10\] 0
C7888 _0157_ _1060_/a_891_413# 0.00127f
C7889 _1059_/a_891_413# _0158_ 0
C7890 _0983_/a_27_47# _0983_/a_561_413# 0.00163f
C7891 _0983_/a_634_159# _0983_/a_891_413# 0.03684f
C7892 _0983_/a_193_47# _0983_/a_381_47# 0.09799f
C7893 _0820_/a_215_47# hold67/a_285_47# 0.00236f
C7894 clknet_1_0__leaf__0465_ _1051_/a_466_413# 0.004f
C7895 _0349_ _0327_ 0
C7896 output41/a_27_47# pp[14] 0.15413f
C7897 pp[15] acc0.A\[31\] 0
C7898 hold88/a_49_47# _0350_ 0
C7899 clknet_1_0__leaf__0465_ _1045_/a_891_413# 0.00129f
C7900 _0758_/a_297_297# _0350_ 0.00224f
C7901 _0758_/a_79_21# _0380_ 0.08483f
C7902 hold37/a_49_47# net137 0.00136f
C7903 _0576_/a_109_297# net110 0.0021f
C7904 hold98/a_285_47# _0995_/a_466_413# 0.00566f
C7905 hold98/a_49_47# _0995_/a_1059_315# 0
C7906 hold98/a_391_47# _0995_/a_634_159# 0
C7907 VPWR _0526_/a_27_47# 0.41635f
C7908 _0457_ _1014_/a_27_47# 0
C7909 hold37/a_285_47# net184 0.00978f
C7910 hold37/a_391_47# net131 0.05532f
C7911 _0985_/a_27_47# net71 0.22754f
C7912 _0399_ _0507_/a_373_47# 0
C7913 _0538_/a_149_47# comp0.B\[12\] 0
C7914 net21 _0954_/a_32_297# 0
C7915 pp[30] net116 0.10736f
C7916 _0180_ _0446_ 0.00398f
C7917 VPWR net9 1.38359f
C7918 _1015_/a_634_159# _0566_/a_27_47# 0
C7919 _0606_/a_109_53# _0237_ 0.09772f
C7920 _1056_/a_27_47# hold35/a_285_47# 0.01366f
C7921 _1056_/a_193_47# hold35/a_49_47# 0.00127f
C7922 _0267_ clkbuf_0__0458_/a_110_47# 0.01722f
C7923 _0206_ _0205_ 0.00478f
C7924 net194 _0180_ 0.00508f
C7925 _0637_/a_56_297# _0268_ 0.09033f
C7926 _1020_/a_592_47# _0183_ 0.00227f
C7927 hold97/a_49_47# _0320_ 0
C7928 _1003_/a_193_47# _0183_ 0
C7929 _1003_/a_1059_315# net150 0
C7930 _1003_/a_466_413# _0217_ 0.00317f
C7931 _0104_ _0326_ 0
C7932 net103 net166 0.05281f
C7933 _1013_/a_1059_315# _0218_ 0.00378f
C7934 _1016_/a_466_413# _1016_/a_592_47# 0.00553f
C7935 _1016_/a_634_159# _1016_/a_1017_47# 0
C7936 _1004_/a_1059_315# net176 0
C7937 clkload2/Y _1050_/a_27_47# 0
C7938 _0251_ hold31/a_391_47# 0
C7939 clknet_0__0459_ _0996_/a_27_47# 0.00976f
C7940 pp[10] net37 0.02467f
C7941 _0443_ net62 0.03015f
C7942 clknet_0__0465_ _0823_/a_109_297# 0
C7943 _0378_ acc0.A\[23\] 0
C7944 _0280_ _0290_ 0
C7945 comp0.B\[1\] _0956_/a_304_297# 0.01405f
C7946 _0131_ comp0.B\[15\] 0
C7947 clknet_1_1__leaf__0462_ _1026_/a_634_159# 0
C7948 net113 _1026_/a_27_47# 0.00199f
C7949 _0195_ _0705_/a_59_75# 0
C7950 _1028_/a_1059_315# acc0.A\[28\] 0.12779f
C7951 net188 net189 0.21028f
C7952 _0176_ net127 0
C7953 _0692_/a_113_47# clknet_1_0__leaf__0460_ 0
C7954 _0329_ _0701_/a_80_21# 0.03644f
C7955 _0641_/a_113_47# acc0.A\[6\] 0
C7956 _0238_ _0352_ 0.02819f
C7957 _0176_ _0543_/a_150_297# 0
C7958 _0363_ _0361_ 0.0036f
C7959 VPWR _0990_/a_1017_47# 0
C7960 _0812_/a_510_47# _0090_ 0
C7961 net56 _0333_ 0.02548f
C7962 _0999_/a_592_47# _0096_ 0
C7963 _0327_ _0701_/a_209_297# 0.09968f
C7964 _0846_/a_51_297# _0261_ 0
C7965 hold97/a_285_47# clknet_1_1__leaf__0462_ 0
C7966 VPWR _0793_/a_240_47# 0.00621f
C7967 input30/a_75_212# B[7] 0.19873f
C7968 clkbuf_1_1__f__0460_/a_110_47# _0318_ 0.02018f
C7969 net88 clknet_1_0__leaf__0461_ 0
C7970 _0749_/a_299_297# _0346_ 0.0031f
C7971 _0326_ _0745_/a_109_47# 0
C7972 _0514_/a_27_297# net2 0.17662f
C7973 _0534_/a_81_21# _0534_/a_299_297# 0.08213f
C7974 VPWR _0175_ 2.27892f
C7975 _0454_ net47 0.23073f
C7976 _0397_ _0777_/a_285_47# 0.0091f
C7977 net39 _0994_/a_1059_315# 0.13798f
C7978 acc0.A\[26\] _1008_/a_27_47# 0
C7979 hold28/a_285_47# _0532_/a_81_21# 0
C7980 hold45/a_391_47# _0179_ 0.02643f
C7981 _0134_ _1037_/a_27_47# 0
C7982 _1032_/a_193_47# _0352_ 0
C7983 hold62/a_49_47# hold62/a_285_47# 0.22264f
C7984 _0584_/a_109_47# net157 0
C7985 _1059_/a_891_413# acc0.A\[14\] 0.05209f
C7986 _0538_/a_245_297# net20 0
C7987 clknet_1_1__leaf__0459_ _1057_/a_27_47# 0.00118f
C7988 _1041_/a_891_413# net7 0.05342f
C7989 _0216_ clknet_1_0__leaf__0457_ 0
C7990 _1057_/a_193_47# acc0.A\[11\] 0
C7991 _0978_/a_109_297# clknet_1_0__leaf_clk 0
C7992 _0190_ _0181_ 0.03915f
C7993 _0460_ net92 0.01902f
C7994 _0198_ _1047_/a_891_413# 0
C7995 _0146_ _1047_/a_634_159# 0
C7996 _1056_/a_193_47# A[9] 0
C7997 _0221_ _0701_/a_80_21# 0
C7998 clknet_1_0__leaf__0462_ _0380_ 0.007f
C7999 hold46/a_391_47# _0139_ 0
C8000 _0483_ _0479_ 0.06901f
C8001 _0753_/a_79_21# _0345_ 0
C8002 _0343_ _0754_/a_51_297# 0
C8003 output65/a_27_47# pp[3] 0.08616f
C8004 hold29/a_285_47# hold29/a_391_47# 0.41909f
C8005 hold20/a_391_47# _0468_ 0
C8006 _0399_ clknet_1_1__leaf__0461_ 0.05179f
C8007 _1054_/a_891_413# VPWR 0.18789f
C8008 _0791_/a_113_297# _0406_ 0.00758f
C8009 _0643_/a_103_199# _0257_ 0
C8010 _0305_ _0306_ 0.01723f
C8011 _0358_ _0195_ 0
C8012 _0517_/a_81_21# net16 0.02706f
C8013 output43/a_27_47# _0797_/a_27_413# 0
C8014 acc0.A\[5\] _0987_/a_634_159# 0.00311f
C8015 _1051_/a_891_413# _0085_ 0
C8016 net137 _0987_/a_381_47# 0
C8017 clknet_0__0464_ _1048_/a_27_47# 0
C8018 clkbuf_1_1__f__0461_/a_110_47# _0777_/a_47_47# 0
C8019 _0316_ acc0.A\[28\] 0.00323f
C8020 _0163_ _1065_/a_27_47# 0.11416f
C8021 net69 net104 0
C8022 _0369_ _1063_/a_27_47# 0
C8023 _1038_/a_1059_315# VPWR 0.38657f
C8024 _0457_ _0195_ 0
C8025 _0707_/a_75_199# _0336_ 0
C8026 _1041_/a_1059_315# A[15] 0
C8027 _0269_ _0347_ 0
C8028 hold45/a_391_47# _0513_/a_81_21# 0
C8029 hold45/a_285_47# _0513_/a_299_297# 0.00228f
C8030 VPWR _0655_/a_297_297# 0
C8031 _1018_/a_381_47# acc0.A\[18\] 0.02574f
C8032 _1034_/a_27_47# net26 0
C8033 _0721_/a_27_47# _0352_ 0.33078f
C8034 _1067_/a_27_47# clknet_1_0__leaf__0457_ 0.07535f
C8035 _0799_/a_80_21# net42 0
C8036 acc0.A\[28\] _0347_ 0
C8037 clkbuf_1_0__f_clk/a_110_47# _0166_ 0
C8038 _0983_/a_193_47# clknet_1_0__leaf__0459_ 0
C8039 clknet_1_0__leaf__0460_ _0618_/a_79_21# 0.0117f
C8040 _0695_/a_217_297# _0250_ 0.05373f
C8041 _0369_ _1060_/a_27_47# 0
C8042 _0824_/a_59_75# _0431_ 0.08088f
C8043 _0209_ net180 0
C8044 _0241_ _0616_/a_78_199# 0.12917f
C8045 hold86/a_285_47# _0264_ 0
C8046 _0957_/a_32_297# net28 0
C8047 _0339_ net116 0
C8048 _0479_ control0.count\[1\] 0.08594f
C8049 hold30/a_391_47# _0121_ 0
C8050 clknet_1_0__leaf__0462_ _0683_/a_113_47# 0
C8051 net7 net147 0.21809f
C8052 pp[17] _0567_/a_27_297# 0
C8053 acc0.A\[24\] acc0.A\[23\] 0.00156f
C8054 net203 _0131_ 0.4432f
C8055 _0369_ _0988_/a_891_413# 0
C8056 _1001_/a_1059_315# _0216_ 0
C8057 _1031_/a_193_47# _1030_/a_27_47# 0
C8058 _1031_/a_27_47# _1030_/a_193_47# 0
C8059 _0400_ net41 0.21143f
C8060 _0817_/a_266_47# _0346_ 0.00751f
C8061 done _1071_/a_1059_315# 0
C8062 net35 _1071_/a_381_47# 0
C8063 _1008_/a_193_47# net244 0.00506f
C8064 net51 _1005_/a_1017_47# 0
C8065 net189 _0155_ 0
C8066 comp0.B\[13\] _1042_/a_1059_315# 0
C8067 _0322_ _0181_ 0
C8068 _1012_/a_27_47# _0395_ 0
C8069 _0235_ _0219_ 0
C8070 _0136_ clkbuf_1_0__f__0463_/a_110_47# 0
C8071 clknet_1_1__leaf__0460_ _0331_ 0.04587f
C8072 _0180_ _0987_/a_193_47# 0
C8073 acc0.A\[5\] net136 0
C8074 _1038_/a_466_413# _0550_/a_51_297# 0
C8075 _1038_/a_27_47# _0550_/a_149_47# 0
C8076 clknet_1_1__leaf__0460_ _0695_/a_300_47# 0
C8077 _0237_ hold3/a_285_47# 0.05782f
C8078 _0381_ hold3/a_391_47# 0.06181f
C8079 _0260_ clknet_1_1__leaf__0458_ 0
C8080 net43 _0308_ 0.00107f
C8081 _0327_ _0181_ 0
C8082 _0154_ acc0.A\[11\] 0
C8083 _0343_ _0995_/a_381_47# 0.00695f
C8084 _0554_/a_68_297# _1037_/a_27_47# 0
C8085 _1014_/a_561_413# clknet_1_0__leaf__0461_ 0.00117f
C8086 _0858_/a_27_47# acc0.A\[1\] 0
C8087 _1025_/a_27_47# _1025_/a_634_159# 0.14145f
C8088 _0726_/a_240_47# _0109_ 0.00134f
C8089 _0354_ _0355_ 0.16928f
C8090 _0216_ _0588_/a_113_47# 0
C8091 _0668_/a_297_47# net6 0
C8092 _0458_ hold71/a_49_47# 0
C8093 clkbuf_1_0__f__0461_/a_110_47# net219 0
C8094 hold82/a_49_47# _0345_ 0.00147f
C8095 _0654_/a_207_413# _0418_ 0
C8096 comp0.B\[1\] _1032_/a_1059_315# 0
C8097 _0287_ _0283_ 0.00552f
C8098 _0437_ net75 0
C8099 _0486_ clknet_1_0__leaf__0460_ 0.006f
C8100 net34 _1064_/a_561_413# 0.002f
C8101 control0.state\[1\] _1064_/a_975_413# 0
C8102 hold55/a_49_47# net202 0.01093f
C8103 hold58/a_285_47# _0133_ 0
C8104 _1050_/a_381_47# _0148_ 0.13104f
C8105 comp0.B\[13\] net10 0.11907f
C8106 net187 net223 0
C8107 hold31/a_49_47# clknet_1_1__leaf__0458_ 0
C8108 _0740_/a_113_47# acc0.A\[25\] 0
C8109 net245 _0413_ 0.17016f
C8110 _0347_ hold72/a_49_47# 0
C8111 hold55/a_49_47# clknet_1_1__leaf__0463_ 0
C8112 _0386_ _0393_ 0
C8113 net58 _0448_ 0.28508f
C8114 _0739_/a_297_297# _0106_ 0
C8115 _0333_ _0345_ 0.20917f
C8116 _0739_/a_510_47# _0365_ 0.00189f
C8117 _1046_/a_193_47# net10 0.07623f
C8118 clknet_0__0457_ _1001_/a_891_413# 0
C8119 net71 _0197_ 0.03607f
C8120 hold76/a_285_47# control0.add 0
C8121 _0515_/a_299_297# _0181_ 0
C8122 _0467_ _1065_/a_891_413# 0.03637f
C8123 net191 net114 0
C8124 _0089_ _0450_ 0
C8125 _0216_ _1047_/a_891_413# 0
C8126 hold95/a_49_47# hold95/a_391_47# 0.00188f
C8127 net8 comp0.B\[9\] 0
C8128 _0996_/a_27_47# _0996_/a_1059_315# 0.04875f
C8129 _0996_/a_193_47# _0996_/a_466_413# 0.07402f
C8130 net36 _1018_/a_193_47# 0
C8131 net125 net7 0.11905f
C8132 _0388_ _0246_ 0
C8133 _0139_ net153 0.13488f
C8134 pp[15] net43 0.00525f
C8135 _0955_/a_32_297# clknet_1_1__leaf_clk 0
C8136 comp0.B\[5\] _1066_/a_891_413# 0
C8137 _0999_/a_1059_315# _0219_ 0.00171f
C8138 hold10/a_49_47# clknet_1_1__leaf__0457_ 0
C8139 _0793_/a_51_297# _0095_ 0.10261f
C8140 _0260_ _0263_ 0
C8141 _0646_/a_129_47# acc0.A\[13\] 0
C8142 _0537_/a_68_297# net196 0
C8143 _0752_/a_27_413# _0377_ 0
C8144 _0234_ _0754_/a_240_47# 0.00199f
C8145 _0376_ _0754_/a_51_297# 0.0761f
C8146 hold55/a_391_47# _0182_ 0
C8147 _0230_ _0382_ 0
C8148 _0559_/a_245_297# _0175_ 0.00307f
C8149 net61 _0180_ 0.01065f
C8150 acc0.A\[7\] input15/a_75_212# 0.00194f
C8151 acc0.A\[16\] _0158_ 0
C8152 VPWR _0996_/a_891_413# 0.18562f
C8153 _1065_/a_891_413# comp0.B\[0\] 0.01625f
C8154 _0743_/a_51_297# clknet_0__0460_ 0
C8155 _0272_ _0346_ 0
C8156 _0726_/a_51_297# acc0.A\[29\] 0.00879f
C8157 _0465_ _0445_ 0.00263f
C8158 VPWR input16/a_75_212# 0.18521f
C8159 _1051_/a_27_47# _1044_/a_381_47# 0
C8160 _1051_/a_381_47# _1044_/a_27_47# 0
C8161 comp0.B\[7\] _0953_/a_32_297# 0.11343f
C8162 _1037_/a_561_413# net28 0
C8163 hold65/a_285_47# _0830_/a_215_47# 0
C8164 _1051_/a_466_413# net137 0
C8165 _1051_/a_634_159# _0149_ 0
C8166 hold22/a_285_47# _1054_/a_27_47# 0.00123f
C8167 _1045_/a_891_413# _1044_/a_466_413# 0
C8168 _1045_/a_1059_315# _1044_/a_1059_315# 0.00135f
C8169 _0302_ _0420_ 0.00247f
C8170 net58 _0444_ 0.01416f
C8171 net104 net102 0
C8172 _0762_/a_79_21# net51 0.0344f
C8173 _0992_/a_634_159# acc0.A\[10\] 0.01088f
C8174 _1030_/a_634_159# _0353_ 0
C8175 _1051_/a_891_413# net131 0
C8176 acc0.A\[9\] _0218_ 0.08143f
C8177 _0210_ _0207_ 0
C8178 net62 _0986_/a_891_413# 0.04318f
C8179 net22 _1040_/a_193_47# 0
C8180 _1045_/a_381_47# net184 0.11464f
C8181 _1045_/a_561_413# net131 0
C8182 net78 _0422_ 0.02921f
C8183 clknet_1_1__leaf__0459_ _0789_/a_544_297# 0.00224f
C8184 _0480_ clknet_1_0__leaf_clk 0.06622f
C8185 _0305_ _0346_ 0.00154f
C8186 net61 _0432_ 0.02426f
C8187 _1072_/a_891_413# clknet_1_0__leaf_clk 0
C8188 _0399_ _0990_/a_193_47# 0.04965f
C8189 VPWR net129 0.39089f
C8190 _0693_/a_68_297# _0693_/a_150_297# 0.00477f
C8191 _0250_ _0345_ 0
C8192 _0643_/a_253_47# _0465_ 0.00197f
C8193 net40 _0298_ 0
C8194 clknet_1_0__leaf__0458_ acc0.A\[14\] 0.02834f
C8195 clknet_1_1__leaf__0459_ _0673_/a_253_297# 0
C8196 net191 _0365_ 0
C8197 _1002_/a_634_159# net240 0
C8198 _1043_/a_381_47# net196 0.12341f
C8199 _1060_/a_466_413# _0506_/a_299_297# 0
C8200 hold49/a_285_47# clknet_1_1__leaf__0464_ 0.00106f
C8201 VPWR _1015_/a_592_47# 0
C8202 _1003_/a_27_47# _0467_ 0
C8203 _0181_ _0306_ 0
C8204 _0458_ _0529_/a_109_297# 0.00405f
C8205 clknet_0__0464_ _0540_/a_149_47# 0
C8206 clknet_1_0__leaf__0463_ _1040_/a_193_47# 0.00837f
C8207 _0275_ _0427_ 0.42054f
C8208 hold3/a_285_47# _1005_/a_27_47# 0
C8209 _0435_ acc0.A\[6\] 0.00634f
C8210 _1021_/a_561_413# net88 0.00169f
C8211 _1021_/a_381_47# _0100_ 0
C8212 _1032_/a_634_159# _1032_/a_1059_315# 0
C8213 _1032_/a_27_47# _1032_/a_381_47# 0.06222f
C8214 _1032_/a_193_47# _1032_/a_891_413# 0.19685f
C8215 _1054_/a_891_413# _1054_/a_1017_47# 0.00617f
C8216 _1054_/a_193_47# net169 0.47759f
C8217 _1054_/a_634_159# net140 0
C8218 _0231_ _0601_/a_68_297# 0.01239f
C8219 _0568_/a_27_297# _0568_/a_109_47# 0.00393f
C8220 _0233_ _0601_/a_150_297# 0
C8221 _1015_/a_466_413# _1015_/a_592_47# 0.00553f
C8222 _1015_/a_634_159# _1015_/a_1017_47# 0
C8223 net46 _0462_ 0.04312f
C8224 _1038_/a_193_47# net29 0.00293f
C8225 _0717_/a_80_21# hold80/a_285_47# 0
C8226 _0717_/a_209_297# hold80/a_49_47# 0
C8227 _0713_/a_27_47# _1015_/a_27_47# 0
C8228 _0748_/a_384_47# _0369_ 0
C8229 clknet_1_1__leaf__0462_ _0689_/a_68_297# 0
C8230 clknet_0__0457_ _0586_/a_27_47# 0
C8231 _0307_ _0394_ 0
C8232 _0108_ _1010_/a_466_413# 0.00187f
C8233 net68 acc0.A\[1\] 0.1516f
C8234 _0753_/a_297_297# clknet_1_0__leaf__0460_ 0.00474f
C8235 clknet_1_1__leaf__0462_ _1027_/a_1017_47# 0
C8236 _0343_ _1031_/a_381_47# 0
C8237 _1014_/a_193_47# net149 0.06053f
C8238 net10 comp0.B\[9\] 0
C8239 net247 _1047_/a_891_413# 0
C8240 _0180_ _1045_/a_27_47# 0
C8241 _1038_/a_891_413# _1038_/a_975_413# 0.00851f
C8242 _1038_/a_27_47# net124 0.22924f
C8243 _1038_/a_381_47# _1038_/a_561_413# 0.00123f
C8244 net19 _0541_/a_68_297# 0.04966f
C8245 _1039_/a_1059_315# _0210_ 0
C8246 _0211_ _1037_/a_1059_315# 0
C8247 _0473_ net7 0.03353f
C8248 _0765_/a_79_21# _0373_ 0
C8249 acc0.A\[14\] acc0.A\[16\] 0
C8250 hold35/a_49_47# clknet_1_1__leaf__0465_ 0
C8251 _0442_ _0836_/a_150_297# 0
C8252 _0319_ _1008_/a_592_47# 0
C8253 _1067_/a_891_413# clknet_1_0__leaf__0461_ 0.01636f
C8254 _1057_/a_193_47# _0281_ 0
C8255 hold19/a_391_47# _0369_ 0
C8256 _0655_/a_109_93# _0286_ 0.06485f
C8257 _0655_/a_297_297# _0283_ 0
C8258 pp[30] _0220_ 0.04246f
C8259 input20/a_75_212# comp0.B\[11\] 0.03737f
C8260 _0268_ _0849_/a_79_21# 0.00248f
C8261 _0637_/a_56_297# net222 0
C8262 _0346_ hold73/a_49_47# 0.00402f
C8263 _0269_ _0824_/a_59_75# 0
C8264 _0983_/a_891_413# net69 0
C8265 _0490_ control0.state\[2\] 0
C8266 clknet_1_0__leaf__0465_ _0149_ 0.02707f
C8267 hold36/a_49_47# hold36/a_285_47# 0.22264f
C8268 _0289_ _0673_/a_103_199# 0.11028f
C8269 hold37/a_285_47# net130 0
C8270 _0661_/a_109_297# _0295_ 0
C8271 _0200_ net31 0
C8272 clknet_1_0__leaf__0462_ _0590_/a_113_47# 0
C8273 _0218_ _0449_ 0
C8274 _0752_/a_27_413# net109 0
C8275 VPWR output50/a_27_47# 0.292f
C8276 net9 _0523_/a_81_21# 0
C8277 clknet_0__0461_ _0347_ 0.04834f
C8278 clkbuf_1_0__f__0461_/a_110_47# _0352_ 0
C8279 _0891_/a_27_47# _0181_ 0.00312f
C8280 _0262_ _0448_ 0
C8281 net40 _0995_/a_1017_47# 0
C8282 VPWR _0840_/a_68_297# 0.16763f
C8283 _0286_ _0418_ 0.14303f
C8284 _0461_ hold40/a_49_47# 0
C8285 _0454_ _0294_ 0
C8286 _0984_/a_1059_315# acc0.A\[14\] 0
C8287 clknet_1_1__leaf__0460_ _1008_/a_27_47# 0
C8288 net31 comp0.B\[8\] 0
C8289 hold45/a_49_47# net4 0
C8290 hold64/a_285_47# clknet_1_0__leaf__0457_ 0.00224f
C8291 _0997_/a_1059_315# net42 0.15991f
C8292 hold37/a_49_47# _0148_ 0
C8293 _0230_ _0600_/a_253_47# 0.0556f
C8294 _0550_/a_51_297# _0550_/a_240_47# 0.03076f
C8295 _0113_ _0526_/a_27_47# 0
C8296 net216 _1006_/a_27_47# 0.00288f
C8297 control0.reset acc0.A\[15\] 0
C8298 _0238_ _0237_ 0
C8299 net106 _1032_/a_193_47# 0.00109f
C8300 _0466_ _1068_/a_592_47# 0.00306f
C8301 acc0.A\[12\] _1058_/a_634_159# 0.03564f
C8302 _0459_ net6 0.07417f
C8303 _1031_/a_891_413# net60 0
C8304 _0835_/a_215_47# acc0.A\[3\] 0
C8305 hold32/a_285_47# _1055_/a_27_47# 0.00403f
C8306 _0452_ _0266_ 0.06626f
C8307 _0101_ _0217_ 0.02612f
C8308 hold14/a_49_47# _0556_/a_68_297# 0
C8309 _1054_/a_466_413# acc0.A\[6\] 0
C8310 _1054_/a_27_47# net13 0
C8311 A[9] clknet_1_1__leaf__0465_ 0.00143f
C8312 _0330_ _0329_ 1.22317f
C8313 _0294_ _0505_/a_27_297# 0.00673f
C8314 clknet_1_0__leaf__0462_ _1005_/a_891_413# 0.01681f
C8315 VPWR _0955_/a_114_297# 0.01299f
C8316 _0643_/a_103_199# clknet_1_1__leaf__0458_ 0.01306f
C8317 hold33/a_49_47# _0953_/a_32_297# 0.00159f
C8318 _0553_/a_240_47# net28 0
C8319 _0386_ net206 0
C8320 _1061_/a_891_413# acc0.A\[15\] 0.00379f
C8321 _0247_ _0614_/a_183_297# 0
C8322 _1036_/a_27_47# _0175_ 0.00352f
C8323 _0313_ _0739_/a_79_21# 0.00108f
C8324 clknet_1_1__leaf__0462_ net112 0
C8325 net76 net66 0
C8326 _0998_/a_381_47# _0096_ 0.12675f
C8327 _0998_/a_561_413# _0399_ 0
C8328 _0567_/a_27_297# _0567_/a_109_297# 0.17136f
C8329 _0230_ _0751_/a_29_53# 0
C8330 control0.count\[2\] _0168_ 0
C8331 hold22/a_391_47# VPWR 0.17343f
C8332 comp0.B\[4\] _0552_/a_68_297# 0
C8333 _0780_/a_285_297# _0394_ 0.00396f
C8334 _0732_/a_80_21# net52 0
C8335 clknet_0__0465_ acc0.A\[8\] 0
C8336 _0216_ _0499_/a_59_75# 0
C8337 _0186_ _0825_/a_150_297# 0
C8338 _1036_/a_193_47# control0.sh 0
C8339 comp0.B\[4\] _1066_/a_193_47# 0
C8340 hold54/a_49_47# comp0.B\[15\] 0.00421f
C8341 _0399_ clkbuf_1_1__f__0459_/a_110_47# 0.00398f
C8342 _0131_ _0176_ 0.00761f
C8343 _0773_/a_35_297# _0773_/a_285_47# 0.00723f
C8344 _0532_/a_299_297# clkbuf_1_0__f__0464_/a_110_47# 0
C8345 net167 _0467_ 0
C8346 _0217_ hold4/a_285_47# 0.03206f
C8347 acc0.A\[22\] hold4/a_49_47# 0.03552f
C8348 net2 _0189_ 0.01672f
C8349 acc0.A\[20\] _0749_/a_384_47# 0
C8350 _0330_ _0221_ 0
C8351 _1008_/a_466_413# hold50/a_391_47# 0
C8352 net61 pp[7] 0.00226f
C8353 _1052_/a_466_413# net11 0
C8354 input10/a_75_212# B[11] 0
C8355 _0082_ _0347_ 0
C8356 _0645_/a_285_47# _0301_ 0
C8357 _0982_/a_27_47# _1014_/a_1059_315# 0.00102f
C8358 _0985_/a_381_47# _0219_ 0
C8359 net193 net31 0
C8360 net183 _0142_ 0
C8361 _0195_ _1017_/a_1059_315# 0.05801f
C8362 net160 _1035_/a_975_413# 0
C8363 _0397_ _0219_ 0.02415f
C8364 hold64/a_49_47# _1001_/a_891_413# 0
C8365 clknet_1_0__leaf__0460_ _0242_ 0
C8366 net70 _0218_ 0
C8367 _0618_/a_79_21# hold94/a_285_47# 0
C8368 hold39/a_391_47# _0173_ 0.03555f
C8369 hold42/a_285_47# VPWR 0.2667f
C8370 _0180_ net132 0
C8371 _0294_ _0506_/a_81_21# 0.00232f
C8372 _1016_/a_891_413# clknet_0__0461_ 0
C8373 _1057_/a_1059_315# VPWR 0.39023f
C8374 _1048_/a_1059_315# _0186_ 0
C8375 _0346_ _0181_ 0.67839f
C8376 _0732_/a_209_297# clknet_1_0__leaf__0460_ 0
C8377 clkbuf_1_0__f__0460_/a_110_47# net52 0.03602f
C8378 hold29/a_285_47# net50 0.07997f
C8379 clkbuf_1_1__f__0462_/a_110_47# _1008_/a_193_47# 0
C8380 _0233_ _0377_ 0
C8381 _0343_ _0219_ 0.33505f
C8382 _0598_/a_79_21# _0762_/a_79_21# 0
C8383 _0808_/a_81_21# _0806_/a_113_297# 0
C8384 clkbuf_0__0459_/a_110_47# net41 0
C8385 net47 _0184_ 0
C8386 _0464_ _0147_ 0
C8387 _0362_ _1009_/a_193_47# 0
C8388 net44 _0096_ 0
C8389 _0274_ _0258_ 0.02235f
C8390 _0548_/a_51_297# _0543_/a_68_297# 0
C8391 _0222_ _0606_/a_109_53# 0
C8392 _0250_ net52 0.02661f
C8393 acc0.A\[5\] net73 0
C8394 net95 _0219_ 0
C8395 VPWR acc0.A\[29\] 2.28054f
C8396 net63 _0152_ 0.00167f
C8397 _0399_ _0438_ 0.09917f
C8398 acc0.A\[12\] _0787_/a_209_297# 0
C8399 _0366_ _1007_/a_466_413# 0.05602f
C8400 _0315_ _1007_/a_634_159# 0
C8401 _0367_ _1007_/a_193_47# 0
C8402 comp0.B\[10\] _0540_/a_51_297# 0
C8403 hold5/a_391_47# net152 0.13587f
C8404 hold5/a_285_47# net32 0
C8405 net1 _1064_/a_1059_315# 0
C8406 _0339_ _0220_ 0.38458f
C8407 _0992_/a_466_413# _0181_ 0
C8408 _0338_ _0336_ 0.1876f
C8409 net11 _0194_ 0
C8410 net76 _0350_ 0.33263f
C8411 pp[6] _0621_/a_285_297# 0
C8412 hold69/a_49_47# hold69/a_391_47# 0.00188f
C8413 _0522_/a_27_297# _0522_/a_373_47# 0.01338f
C8414 _0252_ net75 0.20495f
C8415 _0805_/a_109_47# _0402_ 0.00151f
C8416 _0179_ _1061_/a_891_413# 0
C8417 _1001_/a_193_47# _0580_/a_27_297# 0
C8418 _0800_/a_51_297# _0800_/a_245_297# 0.01218f
C8419 _0989_/a_381_47# net75 0
C8420 net35 _1072_/a_975_413# 0
C8421 clknet_0__0457_ net149 0.1271f
C8422 hold57/a_49_47# _0174_ 0.04567f
C8423 _0181_ _0935_/a_27_47# 0
C8424 _0314_ _0574_/a_27_297# 0
C8425 _1017_/a_466_413# _0369_ 0.01148f
C8426 _0225_ _1023_/a_193_47# 0
C8427 _1052_/a_1059_315# hold7/a_285_47# 0.0011f
C8428 net44 _1031_/a_193_47# 0
C8429 _0304_ _0671_/a_113_297# 0.07454f
C8430 _0458_ net170 0.00415f
C8431 _0473_ comp0.B\[11\] 0
C8432 VPWR _0699_/a_68_297# 0.17799f
C8433 _0672_/a_215_47# _0303_ 0.00331f
C8434 _0607_/a_373_47# _0347_ 0
C8435 _0607_/a_27_297# _0352_ 0.05881f
C8436 _0965_/a_377_297# _0466_ 0
C8437 hold14/a_49_47# _0134_ 0.37302f
C8438 _0275_ _0818_/a_193_47# 0.00378f
C8439 _0760_/a_285_47# _0237_ 0.08574f
C8440 _0760_/a_377_297# _0382_ 0.00214f
C8441 _0172_ control0.sh 0
C8442 net178 _0988_/a_466_413# 0.02276f
C8443 net126 net8 0
C8444 _0217_ _0582_/a_109_297# 0.02104f
C8445 _0803_/a_68_297# _0281_ 0
C8446 _0458_ _0845_/a_109_297# 0.00105f
C8447 _0982_/a_1059_315# hold18/a_391_47# 0
C8448 _0982_/a_891_413# hold18/a_285_47# 0.00147f
C8449 _0476_ _0950_/a_75_212# 0
C8450 _1053_/a_891_413# _0152_ 0
C8451 _1012_/a_193_47# _0306_ 0.00131f
C8452 _0983_/a_466_413# _0399_ 0.03102f
C8453 _0217_ net23 0
C8454 _0457_ _1067_/a_592_47# 0
C8455 net51 _1022_/a_634_159# 0
C8456 hold58/a_285_47# _0208_ 0
C8457 _0328_ _0367_ 0
C8458 hold35/a_391_47# input16/a_75_212# 0
C8459 clknet_1_0__leaf__0463_ _1061_/a_1059_315# 0
C8460 hold68/a_49_47# net176 0.13693f
C8461 net64 clknet_0__0465_ 0.0019f
C8462 net8 input8/a_75_212# 0.11546f
C8463 net187 clkbuf_0__0457_/a_110_47# 0.00119f
C8464 _0498_/a_149_47# _0177_ 0.00154f
C8465 net7 _0497_/a_68_297# 0
C8466 _1038_/a_466_413# _0172_ 0
C8467 net172 _0550_/a_51_297# 0.003f
C8468 _1038_/a_193_47# _0137_ 0
C8469 clknet_1_0__leaf__0463_ _0207_ 0.09062f
C8470 _0210_ _1037_/a_1059_315# 0
C8471 net160 _1037_/a_891_413# 0
C8472 _1025_/a_891_413# _1025_/a_975_413# 0.00851f
C8473 _1025_/a_381_47# _1025_/a_561_413# 0.00123f
C8474 _0499_/a_59_75# net247 0
C8475 net5 _0669_/a_29_53# 0
C8476 _1012_/a_1017_47# _0345_ 0
C8477 _1030_/a_27_47# _0221_ 0
C8478 _0984_/a_193_47# _0347_ 0
C8479 _0183_ _0869_/a_27_47# 0.00361f
C8480 _0973_/a_27_297# _1067_/a_634_159# 0
C8481 clknet_0__0458_ _0186_ 0.04091f
C8482 clknet_0__0465_ _0423_ 0
C8483 net120 net24 0
C8484 hold25/a_285_47# _0136_ 0.00355f
C8485 _0982_/a_1059_315# _0195_ 0.00448f
C8486 hold54/a_391_47# _0551_/a_27_47# 0
C8487 _1055_/a_592_47# _0181_ 0
C8488 output42/a_27_47# net5 0
C8489 comp0.B\[0\] _0214_ 0
C8490 _0247_ _0391_ 0.00199f
C8491 control0.count\[1\] _0976_/a_218_47# 0.00155f
C8492 _1070_/a_1017_47# _0488_ 0
C8493 acc0.A\[4\] _0148_ 0.15373f
C8494 _0413_ VPWR 0.29964f
C8495 acc0.A\[12\] _0664_/a_297_47# 0
C8496 _0516_/a_27_297# clknet_1_1__leaf__0465_ 0.0577f
C8497 _0157_ net228 0.01178f
C8498 comp0.B\[3\] _0175_ 0.21205f
C8499 _0236_ _1006_/a_27_47# 0
C8500 net123 B[1] 0
C8501 _0972_/a_584_47# _1063_/a_27_47# 0
C8502 _0403_ _0994_/a_381_47# 0
C8503 _0217_ net35 0.04596f
C8504 acc0.A\[0\] _0265_ 0
C8505 _0314_ _0326_ 0
C8506 acc0.A\[14\] _0670_/a_215_47# 0.05353f
C8507 _0557_/a_51_297# net25 0
C8508 _0539_/a_150_297# net19 0
C8509 _0473_ _0202_ 0
C8510 _0996_/a_891_413# _0996_/a_1017_47# 0.00617f
C8511 _0812_/a_215_47# hold70/a_285_47# 0
C8512 _0432_ _0431_ 0.03552f
C8513 _0998_/a_193_47# _0219_ 0
C8514 VPWR _0827_/a_109_297# 0.0034f
C8515 _0314_ _1025_/a_634_159# 0
C8516 VPWR _0255_ 4.23448f
C8517 hold5/a_285_47# net10 0.02192f
C8518 output47/a_27_47# net47 0.20028f
C8519 clkload2/a_268_47# clknet_1_0__leaf__0465_ 0
C8520 _0218_ _0771_/a_298_297# 0
C8521 _0472_ _0138_ 0
C8522 _0581_/a_27_297# _0247_ 0.02243f
C8523 _1018_/a_27_47# _0346_ 0
C8524 _0294_ _0310_ 0.21817f
C8525 _0376_ _0219_ 0.00246f
C8526 _0172_ net157 0.12636f
C8527 _0158_ _0505_/a_109_297# 0.00746f
C8528 net146 _0505_/a_109_47# 0.00265f
C8529 _1060_/a_381_47# net6 0
C8530 acc0.A\[16\] _1016_/a_634_159# 0
C8531 pp[0] _0209_ 0
C8532 hold79/a_49_47# _0978_/a_27_297# 0.01013f
C8533 _0714_/a_51_297# _0342_ 0.08381f
C8534 _0812_/a_79_21# net67 0.07255f
C8535 acc0.A\[27\] _0359_ 0
C8536 net182 input16/a_75_212# 0
C8537 clkbuf_0__0458_/a_110_47# _0347_ 0
C8538 clknet_1_0__leaf__0463_ _1039_/a_1059_315# 0.00304f
C8539 clkbuf_1_1__f__0464_/a_110_47# _0202_ 0
C8540 VPWR _1036_/a_381_47# 0.07547f
C8541 hold54/a_391_47# _0533_/a_27_297# 0
C8542 comp0.B\[7\] _0174_ 0.05235f
C8543 hold24/a_49_47# _0136_ 0
C8544 clknet_0__0457_ _0982_/a_466_413# 0
C8545 clknet_1_1__leaf__0461_ _0306_ 0.0011f
C8546 _1044_/a_193_47# _1044_/a_381_47# 0.09799f
C8547 _1044_/a_634_159# _1044_/a_891_413# 0.03684f
C8548 _1044_/a_27_47# _1044_/a_561_413# 0.0027f
C8549 _0596_/a_145_75# _0227_ 0.00256f
C8550 net101 _0584_/a_27_297# 0.00331f
C8551 B[7] _0176_ 0
C8552 _1038_/a_193_47# comp0.B\[6\] 0.03389f
C8553 net145 _0347_ 0
C8554 _0815_/a_113_297# _0290_ 0.05008f
C8555 _1056_/a_193_47# _0190_ 0
C8556 net137 _0149_ 0.05923f
C8557 _1051_/a_1017_47# acc0.A\[5\] 0
C8558 net44 _0395_ 0.02536f
C8559 net131 _1044_/a_381_47# 0
C8560 _0222_ hold3/a_285_47# 0
C8561 hold59/a_391_47# net234 0
C8562 clknet_1_0__leaf__0462_ _0592_/a_150_297# 0
C8563 _0548_/a_149_47# _0206_ 0.00154f
C8564 _0399_ clknet_1_1__leaf__0465_ 0.50021f
C8565 _0278_ output40/a_27_47# 0
C8566 _0363_ VPWR 0.37425f
C8567 net46 _1023_/a_891_413# 0.0174f
C8568 _1067_/a_634_159# net17 0.00385f
C8569 hold49/a_49_47# _0202_ 0.00582f
C8570 _0442_ _0252_ 0
C8571 _1057_/a_27_47# _1057_/a_634_159# 0.14145f
C8572 _0259_ _0627_/a_297_297# 0
C8573 VPWR _0754_/a_512_297# 0.00705f
C8574 net88 net240 0.07284f
C8575 _1039_/a_561_413# clknet_0__0463_ 0
C8576 _0369_ _0094_ 0.05288f
C8577 _0158_ _0506_/a_299_297# 0.00194f
C8578 _0260_ _0218_ 0.06914f
C8579 _0854_/a_79_21# net206 0
C8580 _1059_/a_27_47# _1059_/a_634_159# 0.14145f
C8581 _0800_/a_51_297# _0995_/a_27_47# 0
C8582 _0575_/a_109_297# pp[24] 0
C8583 _0575_/a_373_47# net52 0
C8584 acc0.A\[14\] _0455_ 0
C8585 net166 hold72/a_391_47# 0
C8586 comp0.B\[2\] _1065_/a_193_47# 0
C8587 hold101/a_285_47# _0271_ 0
C8588 _0259_ _0817_/a_266_47# 0
C8589 _0458_ _0532_/a_81_21# 0
C8590 _0858_/a_27_47# _0198_ 0
C8591 _0849_/a_79_21# net222 0.11722f
C8592 hold100/a_285_47# net247 0.00868f
C8593 _0517_/a_81_21# net142 0.00533f
C8594 _0267_ _0447_ 0
C8595 _0500_/a_27_47# _1047_/a_193_47# 0.00143f
C8596 _1032_/a_466_413# net202 0
C8597 pp[15] net40 0.01113f
C8598 _1015_/a_592_47# _0113_ 0.00188f
C8599 _0344_ _1030_/a_27_47# 0
C8600 _0982_/a_634_159# net247 0
C8601 _0317_ _0729_/a_68_297# 0
C8602 _1032_/a_466_413# clknet_1_1__leaf__0463_ 0
C8603 net67 _0347_ 0.11249f
C8604 VPWR A[7] 0.21796f
C8605 _0134_ _0208_ 0.01099f
C8606 net178 _0186_ 0.0021f
C8607 _0179_ _1058_/a_193_47# 0
C8608 _0328_ _0742_/a_299_297# 0
C8609 _1051_/a_592_47# _0180_ 0.00157f
C8610 acc0.A\[14\] _0505_/a_109_297# 0.0015f
C8611 hold46/a_49_47# _0540_/a_149_47# 0
C8612 _0649_/a_113_47# VPWR 0
C8613 net214 _0990_/a_27_47# 0
C8614 _0570_/a_27_297# _0320_ 0
C8615 _0386_ _0773_/a_35_297# 0.15174f
C8616 net33 _1066_/a_1017_47# 0.00161f
C8617 hold46/a_391_47# net173 0.00151f
C8618 comp0.B\[7\] _0208_ 0
C8619 _0718_/a_47_47# _0220_ 0.0567f
C8620 _0765_/a_510_47# _0352_ 0.00251f
C8621 hold86/a_285_47# _0846_/a_51_297# 0
C8622 _0551_/a_27_47# _0182_ 0.00241f
C8623 _0343_ _1055_/a_1059_315# 0
C8624 _0125_ _1028_/a_27_47# 0.00504f
C8625 acc0.A\[27\] _1028_/a_466_413# 0.00815f
C8626 comp0.B\[14\] _0954_/a_220_297# 0.00188f
C8627 _0287_ _0345_ 0.11725f
C8628 _0292_ _0814_/a_181_47# 0
C8629 control0.count\[2\] _0976_/a_439_47# 0
C8630 _1034_/a_466_413# net24 0
C8631 _0536_/a_240_47# _0159_ 0
C8632 _0200_ net7 0
C8633 acc0.A\[20\] hold73/a_285_47# 0.01795f
C8634 _0373_ net92 0.00139f
C8635 _0129_ _1030_/a_891_413# 0.00349f
C8636 net163 _1030_/a_466_413# 0
C8637 net97 _0347_ 0
C8638 _0768_/a_27_47# _0294_ 0
C8639 net168 _1052_/a_891_413# 0
C8640 _0375_ acc0.A\[23\] 0.10855f
C8641 _0997_/a_592_47# net43 0.00248f
C8642 net205 net27 0
C8643 _0227_ _0383_ 0.20608f
C8644 _0352_ _1006_/a_891_413# 0.017f
C8645 _0570_/a_109_297# clknet_1_1__leaf__0462_ 0.00553f
C8646 pp[1] _0988_/a_1059_315# 0
C8647 VPWR _0995_/a_975_413# 0.00489f
C8648 _0284_ _0993_/a_891_413# 0.00108f
C8649 _0399_ _0452_ 0
C8650 _0769_/a_299_297# clkbuf_1_0__f__0461_/a_110_47# 0
C8651 _0216_ _0246_ 0.01399f
C8652 _0343_ _0799_/a_209_297# 0.00658f
C8653 hold78/a_285_47# net45 0.01239f
C8654 net23 _0164_ 0
C8655 hold101/a_49_47# acc0.A\[4\] 0
C8656 hold64/a_49_47# net149 0
C8657 _1056_/a_27_47# net214 0
C8658 net7 comp0.B\[8\] 0.16163f
C8659 net192 _0187_ 0.09086f
C8660 _0156_ net4 0.22611f
C8661 clkbuf_0__0465_/a_110_47# clkbuf_0__0458_/a_110_47# 0
C8662 _0663_/a_207_413# _0290_ 0.20633f
C8663 _0663_/a_27_413# _0401_ 0
C8664 _0183_ _0460_ 0.03484f
C8665 _0550_/a_240_47# _0172_ 0.03767f
C8666 _0550_/a_512_297# _0137_ 0.00257f
C8667 clknet_1_0__leaf__0458_ _0534_/a_384_47# 0
C8668 _0240_ _0393_ 0.03701f
C8669 _0533_/a_27_297# _0182_ 0.09638f
C8670 _0533_/a_109_297# acc0.A\[1\] 0.0015f
C8671 hold43/a_49_47# net190 0
C8672 _0951_/a_209_311# _1062_/a_193_47# 0
C8673 _0951_/a_109_93# _1062_/a_634_159# 0.00498f
C8674 _0355_ _0353_ 0.02753f
C8675 _0369_ _0393_ 0
C8676 _0180_ _0269_ 0
C8677 acc0.A\[1\] hold71/a_49_47# 0.30279f
C8678 acc0.A\[12\] net144 0
C8679 _0183_ _1060_/a_193_47# 0.03898f
C8680 clknet_0__0463_ _0957_/a_32_297# 0.00139f
C8681 acc0.A\[24\] _1007_/a_466_413# 0
C8682 hold33/a_49_47# _0174_ 0
C8683 _0723_/a_297_47# _0334_ 0.001f
C8684 hold24/a_391_47# _0206_ 0
C8685 net169 acc0.A\[6\] 0.00815f
C8686 B[12] _0542_/a_512_297# 0
C8687 hold64/a_391_47# _0241_ 0
C8688 _1000_/a_592_47# _0461_ 0
C8689 hold53/a_285_47# _1024_/a_193_47# 0
C8690 hold53/a_391_47# _1024_/a_27_47# 0
C8691 _0511_/a_81_21# acc0.A\[11\] 0.01357f
C8692 _0294_ _0184_ 0
C8693 net55 acc0.A\[27\] 0.4342f
C8694 _0261_ clknet_1_1__leaf__0457_ 0.00229f
C8695 _1031_/a_27_47# _0567_/a_27_297# 0.00819f
C8696 _0616_/a_78_199# _0352_ 0
C8697 _0274_ net72 0
C8698 hold33/a_391_47# comp0.B\[10\] 0
C8699 _0546_/a_51_297# net152 0.09302f
C8700 _1047_/a_1059_315# clkbuf_1_1__f__0457_/a_110_47# 0.00985f
C8701 VPWR _1023_/a_381_47# 0.07577f
C8702 clknet_1_0__leaf__0464_ _0142_ 0.00424f
C8703 hold100/a_391_47# _0846_/a_240_47# 0
C8704 net248 net63 0.10285f
C8705 hold38/a_391_47# net23 0
C8706 clknet_1_1__leaf__0462_ hold50/a_285_47# 0.00803f
C8707 _0183_ _0457_ 0.18518f
C8708 _0991_/a_466_413# _0991_/a_561_413# 0.00772f
C8709 _0991_/a_634_159# _0991_/a_975_413# 0
C8710 _0992_/a_466_413# _0187_ 0
C8711 comp0.B\[14\] _0540_/a_149_47# 0.00598f
C8712 _0554_/a_68_297# _0208_ 0.00411f
C8713 _0627_/a_109_93# _0186_ 0
C8714 net21 net19 0.60035f
C8715 _0370_ _1006_/a_27_47# 0
C8716 _0195_ _0727_/a_109_47# 0
C8717 _0794_/a_27_47# _0297_ 0.04861f
C8718 _0432_ _0269_ 0.32115f
C8719 _0902_/a_27_47# _0462_ 0.11064f
C8720 _0216_ _1029_/a_466_413# 0.01353f
C8721 hold11/a_285_47# _0177_ 0
C8722 clkbuf_0__0463_/a_110_47# _0562_/a_68_297# 0.00115f
C8723 _0210_ _0472_ 0.00805f
C8724 net160 _0475_ 0.0107f
C8725 _0375_ _0602_/a_113_47# 0
C8726 hold78/a_285_47# _0587_/a_27_47# 0
C8727 net193 net7 0
C8728 _0295_ clknet_1_1__leaf__0465_ 0
C8729 _0799_/a_80_21# net5 0.0839f
C8730 _0404_ _0407_ 0
C8731 _0793_/a_240_47# _0345_ 0
C8732 _0793_/a_51_297# _0219_ 0.13981f
C8733 _0080_ _1014_/a_193_47# 0.00432f
C8734 net68 _1014_/a_634_159# 0.00124f
C8735 _0982_/a_634_159# net100 0
C8736 _1004_/a_193_47# acc0.A\[23\] 0.0011f
C8737 clkbuf_1_0__f__0459_/a_110_47# _0219_ 0.03339f
C8738 _0159_ _1046_/a_27_47# 0
C8739 _1001_/a_381_47# _0183_ 0.00747f
C8740 _0195_ _1016_/a_27_47# 0
C8741 clknet_1_0__leaf__0462_ net155 0
C8742 clkbuf_1_1__f__0462_/a_110_47# _0318_ 0.07479f
C8743 net123 _1037_/a_634_159# 0.00174f
C8744 output50/a_27_47# pp[22] 0.15955f
C8745 _0399_ _0996_/a_561_413# 0
C8746 _0731_/a_81_21# _0350_ 0
C8747 _0276_ _0405_ 0
C8748 _0530_/a_299_297# _0465_ 0
C8749 _0230_ _0762_/a_510_47# 0
C8750 _0739_/a_79_21# _0321_ 0
C8751 _0229_ _0369_ 0
C8752 _1021_/a_891_413# _0217_ 0.00426f
C8753 clknet_0__0458_ hold100/a_49_47# 0
C8754 _1041_/a_561_413# clknet_1_0__leaf__0463_ 0
C8755 net173 net153 0
C8756 _1060_/a_193_47# acc0.A\[15\] 0.00621f
C8757 _0348_ _0336_ 0.00807f
C8758 acc0.A\[2\] _0530_/a_299_297# 0.06825f
C8759 _0315_ net93 0.01443f
C8760 _0366_ _0105_ 0.22613f
C8761 hold57/a_285_47# _0555_/a_51_297# 0.00124f
C8762 _0579_/a_27_297# _0713_/a_27_47# 0.01269f
C8763 net53 _1007_/a_27_47# 0.00345f
C8764 _0522_/a_373_47# _0193_ 0.00197f
C8765 _0976_/a_76_199# _0466_ 0.1903f
C8766 _0976_/a_505_21# _0488_ 0.05957f
C8767 hold87/a_391_47# acc0.A\[1\] 0.00424f
C8768 _0800_/a_149_47# _0413_ 0.00869f
C8769 _0800_/a_240_47# _0412_ 0.01395f
C8770 _0305_ net221 0.03534f
C8771 pp[17] _1031_/a_1017_47# 0
C8772 _1011_/a_27_47# _1011_/a_634_159# 0.13832f
C8773 _0655_/a_297_297# _0345_ 0
C8774 net201 _0563_/a_149_47# 0
C8775 _0981_/a_27_297# _0166_ 0.01229f
C8776 VPWR _0830_/a_215_47# 0.00252f
C8777 hold86/a_391_47# _0260_ 0
C8778 A[3] net18 0
C8779 net232 _0972_/a_93_21# 0
C8780 VPWR _1031_/a_975_413# 0.00488f
C8781 _0504_/a_27_47# hold2/a_391_47# 0.00112f
C8782 _0350_ _1006_/a_193_47# 0.05306f
C8783 clknet_0__0465_ _0986_/a_466_413# 0.00477f
C8784 _0216_ _1019_/a_1059_315# 0
C8785 _0643_/a_103_199# _0218_ 0
C8786 acc0.A\[12\] _0648_/a_277_297# 0
C8787 net140 input14/a_75_212# 0.00629f
C8788 _0137_ net29 0
C8789 _1043_/a_1059_315# hold51/a_285_47# 0.00197f
C8790 _1043_/a_891_413# hold51/a_49_47# 0.01135f
C8791 net44 _0221_ 0
C8792 clknet_1_0__leaf__0462_ hold96/a_285_47# 0.01995f
C8793 _0200_ comp0.B\[11\] 0
C8794 hold74/a_49_47# _0459_ 0.00331f
C8795 _1020_/a_634_159# VPWR 0.18237f
C8796 _0350_ _0986_/a_193_47# 0.00959f
C8797 hold12/a_49_47# VPWR 0.3029f
C8798 clknet_0__0458_ net62 0.01257f
C8799 net181 acc0.A\[11\] 0.00361f
C8800 _0971_/a_299_297# _1063_/a_634_159# 0
C8801 clknet_0__0458_ _0450_ 0.28147f
C8802 clkbuf_1_0__f__0458_/a_110_47# _0451_ 0.00146f
C8803 _0835_/a_493_297# _0255_ 0.01135f
C8804 _0183_ _0796_/a_79_21# 0
C8805 _0955_/a_114_297# comp0.B\[3\] 0.00181f
C8806 control0.state\[2\] control0.count\[0\] 0
C8807 _0858_/a_27_47# net247 0
C8808 acc0.A\[31\] _0336_ 0
C8809 net97 hold95/a_49_47# 0
C8810 _0356_ _0334_ 0
C8811 _0789_/a_201_297# _0297_ 0.00594f
C8812 _0150_ _0522_/a_109_47# 0
C8813 _1004_/a_975_413# clknet_1_0__leaf__0460_ 0
C8814 net49 _1022_/a_193_47# 0
C8815 _0429_ hold65/a_285_47# 0
C8816 net55 _1010_/a_193_47# 0.00198f
C8817 control0.reset _0565_/a_240_47# 0
C8818 hold101/a_285_47# clknet_1_0__leaf__0465_ 0.01115f
C8819 net240 _1067_/a_891_413# 0
C8820 _0165_ _1067_/a_634_159# 0.00713f
C8821 _0179_ _1060_/a_193_47# 0
C8822 _0712_/a_79_21# _0567_/a_27_297# 0.00828f
C8823 clknet_1_0__leaf__0458_ _0991_/a_193_47# 0
C8824 control0.state\[2\] _0974_/a_544_297# 0.00161f
C8825 _0486_ _0974_/a_222_93# 0.06821f
C8826 net54 _1008_/a_891_413# 0.04092f
C8827 net194 comp0.B\[12\] 0
C8828 _0278_ _0797_/a_207_413# 0
C8829 _0190_ clknet_1_1__leaf__0465_ 0.12325f
C8830 _0255_ _0523_/a_81_21# 0
C8831 _1010_/a_27_47# _0347_ 0.03635f
C8832 _0632_/a_113_47# _0264_ 0.00963f
C8833 _0972_/a_250_297# _0161_ 0
C8834 hold91/a_391_47# net41 0.07584f
C8835 _1051_/a_27_47# clknet_1_1__leaf__0464_ 0.00932f
C8836 _0531_/a_27_297# _1061_/a_193_47# 0
C8837 _0800_/a_51_297# _0299_ 0
C8838 _0413_ _0789_/a_75_199# 0
C8839 net16 _0088_ 0
C8840 net55 _1009_/a_634_159# 0
C8841 _0384_ _0352_ 0
C8842 _1045_/a_634_159# clknet_1_1__leaf__0464_ 0
C8843 _1036_/a_634_159# _1036_/a_1059_315# 0
C8844 _1036_/a_27_47# _1036_/a_381_47# 0.06222f
C8845 _1036_/a_193_47# _1036_/a_891_413# 0.19685f
C8846 _1056_/a_466_413# _1056_/a_592_47# 0.00553f
C8847 _0218_ _0097_ 0.27901f
C8848 _0346_ _0990_/a_193_47# 0
C8849 _1012_/a_1059_315# clknet_1_1__leaf__0462_ 0
C8850 _1030_/a_891_413# hold61/a_285_47# 0
C8851 _1030_/a_1059_315# hold61/a_391_47# 0.00145f
C8852 _0116_ _0247_ 0.0925f
C8853 _0480_ _0970_/a_27_297# 0
C8854 _0517_/a_81_21# _0988_/a_27_47# 0
C8855 _1012_/a_193_47# _0778_/a_68_297# 0
C8856 hold90/a_391_47# _0319_ 0
C8857 _0459_ _0583_/a_27_297# 0
C8858 _0578_/a_27_297# _0578_/a_109_47# 0.00393f
C8859 net199 acc0.A\[23\] 0
C8860 _1049_/a_193_47# net11 0
C8861 comp0.B\[7\] comp0.B\[9\] 0
C8862 comp0.B\[6\] net29 0.39853f
C8863 _0725_/a_80_21# _0725_/a_209_47# 0.01013f
C8864 _0259_ _0181_ 0.09048f
C8865 pp[9] _0179_ 0
C8866 _0200_ _0202_ 0
C8867 net225 _0342_ 0.00611f
C8868 pp[28] _0723_/a_27_413# 0.01046f
C8869 clknet_1_0__leaf__0463_ _0553_/a_245_297# 0
C8870 _0343_ _0251_ 0
C8871 _1041_/a_1059_315# _0544_/a_240_47# 0
C8872 _1041_/a_891_413# _0544_/a_149_47# 0
C8873 _0845_/a_109_47# _0350_ 0
C8874 VPWR comp0.B\[4\] 0.76062f
C8875 net2 net67 0
C8876 _1050_/a_466_413# net148 0
C8877 _0437_ _0436_ 0.11572f
C8878 _0796_/a_79_21# acc0.A\[15\] 0.00565f
C8879 clknet_0__0457_ _0080_ 0
C8880 _0144_ net173 0
C8881 _0654_/a_207_413# _0417_ 0.00151f
C8882 net160 net27 0.0907f
C8883 _0178_ _1048_/a_561_413# 0
C8884 output56/a_27_47# hold62/a_391_47# 0.00236f
C8885 net193 comp0.B\[11\] 0
C8886 hold11/a_391_47# _0144_ 0.05204f
C8887 _1041_/a_634_159# hold6/a_285_47# 0
C8888 clkbuf_1_0__f__0457_/a_110_47# _0236_ 0.00217f
C8889 _0172_ net13 0
C8890 hold49/a_285_47# _0542_/a_240_47# 0
C8891 _0343_ _0997_/a_891_413# 0
C8892 _0181_ _1062_/a_193_47# 0
C8893 _0995_/a_466_413# _0297_ 0.00476f
C8894 clknet_1_0__leaf__0462_ _1024_/a_27_47# 0.00621f
C8895 _0682_/a_68_297# _1007_/a_1059_315# 0.01364f
C8896 _0467_ _1063_/a_27_47# 0.04954f
C8897 _0402_ acc0.A\[15\] 0
C8898 VPWR _0843_/a_68_297# 0.15385f
C8899 _1052_/a_27_47# _0518_/a_109_297# 0
C8900 pp[0] _1038_/a_891_413# 0
C8901 clknet_1_1__leaf_clk _1065_/a_592_47# 0
C8902 _1049_/a_1059_315# _0465_ 0
C8903 hold47/a_391_47# _0142_ 0.07131f
C8904 _0428_ _0990_/a_634_159# 0
C8905 _0427_ _0990_/a_466_413# 0
C8906 _0467_ _0974_/a_448_47# 0.03486f
C8907 hold86/a_49_47# _0448_ 0.11847f
C8908 _0722_/a_215_47# _0350_ 0
C8909 _0670_/a_510_47# net41 0.00392f
C8910 _0216_ _1028_/a_975_413# 0
C8911 _0195_ _1028_/a_1017_47# 0
C8912 hold34/a_285_47# _0186_ 0
C8913 output67/a_27_47# _0188_ 0.18284f
C8914 _0736_/a_311_297# _0363_ 0.01462f
C8915 _0327_ _0354_ 0
C8916 _0458_ _0846_/a_51_297# 0.00229f
C8917 _1057_/a_891_413# _1057_/a_975_413# 0.00851f
C8918 _1057_/a_381_47# _1057_/a_561_413# 0.00123f
C8919 acc0.A\[2\] _1049_/a_1059_315# 0
C8920 _0502_/a_27_47# _0924_/a_27_47# 0.10738f
C8921 _0553_/a_240_47# clknet_0__0463_ 0
C8922 B[13] _1042_/a_381_47# 0
C8923 _0269_ _0986_/a_381_47# 0
C8924 net44 _0344_ 0
C8925 _0090_ acc0.A\[9\] 0
C8926 pp[30] _0347_ 0
C8927 _0195_ _0534_/a_81_21# 0
C8928 _0343_ net58 0.02464f
C8929 VPWR _1064_/a_592_47# 0
C8930 _0607_/a_109_297# clknet_0__0461_ 0
C8931 _0579_/a_27_297# _0579_/a_109_297# 0.17136f
C8932 _0195_ hold62/a_49_47# 0.00226f
C8933 net57 hold62/a_285_47# 0
C8934 _1059_/a_381_47# _1059_/a_561_413# 0.00123f
C8935 _1059_/a_27_47# net145 0.22944f
C8936 _1059_/a_891_413# _1059_/a_975_413# 0.00851f
C8937 acc0.A\[1\] _0264_ 0.10767f
C8938 net178 net62 0.02917f
C8939 _1041_/a_634_159# _1041_/a_1017_47# 0
C8940 comp0.B\[0\] _1063_/a_27_47# 0
C8941 hold78/a_285_47# VPWR 0.26521f
C8942 net231 _1062_/a_975_413# 0
C8943 hold76/a_391_47# net45 0
C8944 hold41/a_391_47# _0186_ 0
C8945 net36 _0266_ 0.12855f
C8946 _0528_/a_299_297# _0196_ 0.00955f
C8947 _0528_/a_81_21# net170 0.06169f
C8948 _0568_/a_27_297# _0219_ 0.01686f
C8949 hold23/a_391_47# _0195_ 0.00476f
C8950 _0981_/a_109_47# VPWR 0
C8951 _0433_ _0989_/a_634_159# 0
C8952 net68 net247 0
C8953 _0176_ _1042_/a_27_47# 0
C8954 net22 _0472_ 0
C8955 net202 clknet_1_1__leaf__0463_ 0.00914f
C8956 clknet_1_0__leaf_clk _1068_/a_27_47# 0.21626f
C8957 _0673_/a_253_297# _0673_/a_253_47# 0.00137f
C8958 _0181_ net221 0.02295f
C8959 net193 _0202_ 0
C8960 _1002_/a_193_47# _0578_/a_27_297# 0
C8961 comp0.B\[13\] hold48/a_49_47# 0
C8962 net160 _0136_ 0
C8963 _0398_ _0399_ 0.70562f
C8964 _0997_/a_1059_315# net5 0
C8965 _1030_/a_1059_315# clknet_1_1__leaf__0462_ 0
C8966 hold35/a_285_47# net16 0
C8967 hold32/a_49_47# pp[8] 0.04334f
C8968 hold65/a_285_47# clknet_1_1__leaf__0458_ 0.00747f
C8969 _0984_/a_891_413# _0350_ 0.00468f
C8970 _0734_/a_47_47# _0181_ 0
C8971 _0285_ _0403_ 0.00205f
C8972 VPWR _0686_/a_219_297# 0.11276f
C8973 _0496_/a_27_47# _0560_/a_68_297# 0.00183f
C8974 input10/a_75_212# input9/a_27_47# 0.01246f
C8975 _0324_ _1026_/a_193_47# 0
C8976 _1054_/a_634_159# _0087_ 0
C8977 _0138_ _1046_/a_891_413# 0
C8978 VPWR _1008_/a_1059_315# 0.39082f
C8979 net158 _1046_/a_1059_315# 0
C8980 net56 acc0.A\[29\] 0.05827f
C8981 clknet_1_0__leaf__0463_ _0472_ 0.03021f
C8982 _0891_/a_27_47# _1015_/a_27_47# 0.01015f
C8983 _0467_ _1062_/a_1059_315# 0.0025f
C8984 net117 _0341_ 0
C8985 _0216_ _0102_ 0.14125f
C8986 _0682_/a_68_297# clkbuf_1_0__f__0462_/a_110_47# 0.00932f
C8987 _0305_ _1017_/a_27_47# 0
C8988 _0179_ hold47/a_49_47# 0.00714f
C8989 _0268_ _0449_ 0.00201f
C8990 clknet_0__0463_ _0213_ 0.0232f
C8991 _0346_ clkbuf_1_1__f__0459_/a_110_47# 0.01788f
C8992 _0699_/a_68_297# net56 0.10128f
C8993 hold38/a_285_47# _0173_ 0
C8994 hold38/a_391_47# _0213_ 0
C8995 _0399_ _0277_ 0.08696f
C8996 hold33/a_49_47# comp0.B\[9\] 0.05047f
C8997 _0840_/a_68_297# _0345_ 0
C8998 _1010_/a_27_47# hold95/a_49_47# 0
C8999 net162 _0218_ 0
C9000 _0637_/a_311_297# net247 0
C9001 _0467_ _0561_/a_240_47# 0
C9002 _0302_ _0347_ 0
C9003 _0182_ _0199_ 0.74943f
C9004 control0.state\[0\] clk 0.07404f
C9005 comp0.B\[0\] _1062_/a_1059_315# 0
C9006 net213 net51 0.00851f
C9007 _0782_/a_27_47# _0181_ 0
C9008 net45 clknet_1_1__leaf__0462_ 0
C9009 clknet_1_1__leaf__0457_ _0173_ 0
C9010 hold69/a_49_47# _0219_ 0
C9011 pp[18] hold78/a_391_47# 0.00119f
C9012 hold28/a_285_47# clknet_1_1__leaf__0457_ 0
C9013 acc0.A\[24\] _0105_ 0.00919f
C9014 _0275_ _0267_ 0
C9015 VPWR _0563_/a_245_297# 0.00471f
C9016 _0457_ _1034_/a_193_47# 0
C9017 _0804_/a_79_21# _0788_/a_68_297# 0.00157f
C9018 control0.state\[1\] _1063_/a_1059_315# 0.13203f
C9019 net105 _1014_/a_1059_315# 0
C9020 clknet_1_0__leaf__0462_ _1022_/a_975_413# 0
C9021 _1005_/a_27_47# _1005_/a_561_413# 0.0027f
C9022 _1005_/a_634_159# _1005_/a_891_413# 0.03684f
C9023 _1005_/a_193_47# _1005_/a_381_47# 0.09799f
C9024 _0731_/a_81_21# _0731_/a_299_297# 0.08213f
C9025 _0383_ _0352_ 0.08218f
C9026 _0519_/a_299_297# _0519_/a_384_47# 0
C9027 VPWR acc0.A\[23\] 1.16367f
C9028 _0205_ _0139_ 0
C9029 _1047_/a_1017_47# clknet_1_1__leaf__0457_ 0.00148f
C9030 _0984_/a_634_159# net222 0
C9031 net9 input10/a_75_212# 0.00342f
C9032 control0.state\[1\] net159 0
C9033 _1060_/a_27_47# _0507_/a_27_297# 0
C9034 _1013_/a_27_47# _1013_/a_1059_315# 0.04875f
C9035 _1013_/a_193_47# _1013_/a_466_413# 0.07855f
C9036 _0195_ _0400_ 0
C9037 _0438_ _0346_ 0
C9038 _0991_/a_1059_315# net67 0.08398f
C9039 VPWR _0541_/a_150_297# 0.00129f
C9040 _0109_ _0219_ 0.03566f
C9041 VPWR _0746_/a_384_47# 0
C9042 _0339_ _0347_ 0
C9043 _0212_ hold38/a_391_47# 0
C9044 _0399_ _0808_/a_81_21# 0
C9045 _0830_/a_79_21# acc0.A\[6\] 0.06579f
C9046 _0366_ _0359_ 0.1198f
C9047 net65 _0438_ 0
C9048 _0985_/a_891_413# _0261_ 0.02123f
C9049 _0985_/a_1059_315# _0263_ 0
C9050 clknet_1_1__leaf__0459_ _0997_/a_466_413# 0.00534f
C9051 _0286_ _0417_ 0.01079f
C9052 net165 _1060_/a_27_47# 0.009f
C9053 _0583_/a_27_297# _1060_/a_381_47# 0
C9054 _0770_/a_79_21# _0461_ 0
C9055 _0216_ net191 0.25437f
C9056 _0728_/a_59_75# _0109_ 0
C9057 VPWR _0620_/a_113_47# 0
C9058 clknet_1_1__leaf__0459_ _0992_/a_561_413# 0
C9059 VPWR _0989_/a_27_47# 0.73931f
C9060 VPWR hold1/a_49_47# 0.2961f
C9061 _0357_ _0317_ 0
C9062 _0559_/a_240_47# net26 0.06213f
C9063 net68 net100 0.03497f
C9064 _0274_ _0642_/a_298_297# 0
C9065 hold64/a_285_47# _1019_/a_1059_315# 0.01349f
C9066 _0174_ _0203_ 0.06708f
C9067 VPWR _1065_/a_1017_47# 0
C9068 _1038_/a_466_413# _1040_/a_193_47# 0
C9069 _1038_/a_1059_315# _1040_/a_27_47# 0
C9070 VPWR _0992_/a_27_47# 0.67483f
C9071 _0600_/a_337_297# _0223_ 0.00835f
C9072 hold56/a_285_47# hold39/a_285_47# 0.00344f
C9073 _0217_ _0391_ 0
C9074 _0764_/a_299_297# _0373_ 0.06049f
C9075 _1018_/a_891_413# _0582_/a_109_297# 0
C9076 hold35/a_49_47# _0515_/a_81_21# 0
C9077 comp0.B\[10\] net195 0
C9078 clkbuf_0__0462_/a_110_47# _0219_ 0.0878f
C9079 net70 _0268_ 0
C9080 _0995_/a_193_47# _0995_/a_592_47# 0.00135f
C9081 _0995_/a_466_413# _0995_/a_561_413# 0.00772f
C9082 _0995_/a_634_159# _0995_/a_975_413# 0
C9083 clknet_0__0459_ _0301_ 0
C9084 hold10/a_285_47# VPWR 0.28058f
C9085 hold76/a_285_47# net46 0.10026f
C9086 _0137_ comp0.B\[6\] 0
C9087 _0983_/a_27_47# _0853_/a_68_297# 0
C9088 net17 _0951_/a_209_311# 0
C9089 _0119_ _0183_ 0.02309f
C9090 _0565_/a_51_297# clknet_1_0__leaf__0461_ 0.00244f
C9091 _0343_ _0582_/a_109_297# 0.0098f
C9092 hold59/a_49_47# acc0.A\[18\] 0.29155f
C9093 _0983_/a_466_413# _0346_ 0
C9094 hold18/a_285_47# _0350_ 0.02516f
C9095 pp[30] hold95/a_49_47# 0
C9096 net59 hold95/a_391_47# 0
C9097 input6/a_75_212# _0668_/a_297_47# 0
C9098 _1070_/a_634_159# _0489_ 0
C9099 _0534_/a_81_21# _1048_/a_193_47# 0
C9100 VPWR _0549_/a_150_297# 0.00223f
C9101 _1017_/a_193_47# _0675_/a_68_297# 0
C9102 hold64/a_49_47# net206 0
C9103 _0217_ _0581_/a_27_297# 0.10019f
C9104 hold9/a_391_47# _1027_/a_381_47# 0.00142f
C9105 clknet_0_clk _1065_/a_466_413# 0.00332f
C9106 clknet_1_0__leaf__0465_ _1048_/a_193_47# 0
C9107 _0217_ acc0.A\[14\] 0
C9108 net152 _1042_/a_891_413# 0
C9109 net32 _1042_/a_1059_315# 0.00564f
C9110 _0139_ _1042_/a_193_47# 0
C9111 A[12] _0511_/a_81_21# 0
C9112 _1018_/a_634_159# _0459_ 0.00357f
C9113 hold85/a_391_47# control0.state\[2\] 0.00133f
C9114 acc0.A\[29\] _0345_ 0.04148f
C9115 VPWR _1069_/a_193_47# 0.29925f
C9116 _1070_/a_27_47# clknet_1_0__leaf_clk 0.26812f
C9117 control0.reset _0171_ 0.38631f
C9118 _0488_ _0466_ 0.45913f
C9119 control0.state\[0\] _1062_/a_592_47# 0
C9120 VPWR hold60/a_49_47# 0.25944f
C9121 _0982_/a_1059_315# _0183_ 0
C9122 _0298_ _0399_ 0
C9123 comp0.B\[12\] _1045_/a_27_47# 0
C9124 net118 clknet_1_0__leaf__0457_ 0.04057f
C9125 net54 _0320_ 0.2062f
C9126 _0622_/a_109_47# _0252_ 0
C9127 _1011_/a_891_413# _1011_/a_975_413# 0.00851f
C9128 _1011_/a_27_47# net97 0.23034f
C9129 _1011_/a_381_47# _1011_/a_561_413# 0.00123f
C9130 _0608_/a_27_47# _0352_ 0
C9131 _0985_/a_27_47# _0186_ 0.07018f
C9132 _1016_/a_1017_47# _0369_ 0.00146f
C9133 _0133_ _1034_/a_381_47# 0
C9134 _0171_ _1061_/a_891_413# 0
C9135 _0343_ pp[16] 0.11687f
C9136 net176 net177 0
C9137 net57 _0350_ 0
C9138 output37/a_27_47# net4 0.0061f
C9139 _1006_/a_193_47# _1006_/a_634_159# 0.11072f
C9140 _1006_/a_27_47# _1006_/a_466_413# 0.27314f
C9141 clkload2/a_268_47# _0148_ 0
C9142 _0538_/a_51_297# VPWR 0.4786f
C9143 _0240_ _0773_/a_35_297# 0
C9144 _0247_ _0773_/a_285_47# 0
C9145 net32 net10 0.04454f
C9146 _0287_ _0992_/a_891_413# 0
C9147 net45 _0997_/a_561_413# 0
C9148 _0972_/a_256_47# _0487_ 0
C9149 net211 acc0.A\[18\] 0
C9150 _0258_ _0433_ 0.23425f
C9151 _0699_/a_68_297# _0345_ 0
C9152 _0305_ net238 0
C9153 _0316_ hold97/a_49_47# 0
C9154 _0425_ net67 0
C9155 _0201_ _1043_/a_27_47# 0
C9156 hold14/a_391_47# net123 0
C9157 clknet_1_0__leaf__0462_ _0756_/a_47_47# 0.00669f
C9158 _0500_/a_27_47# _0178_ 0.21201f
C9159 _0124_ _1025_/a_634_159# 0
C9160 _0808_/a_81_21# _0808_/a_266_297# 0.01575f
C9161 _1055_/a_381_47# VPWR 0.07818f
C9162 net196 hold51/a_391_47# 0
C9163 _1018_/a_466_413# clknet_1_0__leaf__0461_ 0.01163f
C9164 _0123_ _0217_ 0
C9165 _1001_/a_891_413# acc0.A\[19\] 0.00129f
C9166 net150 output49/a_27_47# 0
C9167 _0102_ _1024_/a_193_47# 0
C9168 _1003_/a_891_413# VPWR 0.19128f
C9169 _0971_/a_81_21# _0161_ 0.01545f
C9170 hold77/a_49_47# hold77/a_285_47# 0.22264f
C9171 net9 _0527_/a_373_47# 0
C9172 hold69/a_49_47# _0746_/a_81_21# 0
C9173 hold97/a_49_47# _0347_ 0
C9174 hold74/a_285_47# _0218_ 0
C9175 _0986_/a_193_47# _0986_/a_634_159# 0.11072f
C9176 _0986_/a_27_47# _0986_/a_466_413# 0.27314f
C9177 net78 _0369_ 0.02448f
C9178 _0585_/a_373_47# _0181_ 0.00164f
C9179 _0299_ _0277_ 0.17432f
C9180 clknet_0__0465_ _0369_ 0
C9181 net148 _0987_/a_466_413# 0.00211f
C9182 _0384_ _0237_ 0
C9183 _0252_ _0436_ 0
C9184 _0432_ clkbuf_0__0458_/a_110_47# 0.01363f
C9185 net236 _0488_ 0.34738f
C9186 _1020_/a_634_159# _0113_ 0
C9187 _0732_/a_209_297# hold90/a_285_47# 0
C9188 clknet_1_1__leaf__0460_ _0460_ 0.11484f
C9189 _1017_/a_27_47# _0181_ 0.02839f
C9190 _1023_/a_193_47# _1023_/a_891_413# 0.19685f
C9191 _1023_/a_27_47# _1023_/a_381_47# 0.06222f
C9192 _1023_/a_634_159# _1023_/a_1059_315# 0
C9193 _0183_ _0451_ 0
C9194 VPWR _0799_/a_303_47# 0
C9195 hold24/a_391_47# A[1] 0
C9196 input22/a_75_212# net153 0
C9197 _1042_/a_634_159# _1042_/a_381_47# 0
C9198 net192 clknet_1_1__leaf__0465_ 0.00489f
C9199 _0181_ _1060_/a_975_413# 0.00124f
C9200 _0403_ _0218_ 0.36438f
C9201 _0516_/a_109_297# net16 0.00906f
C9202 _0423_ _0288_ 0.07221f
C9203 _0401_ acc0.A\[9\] 0.16758f
C9204 _1010_/a_975_413# _0352_ 0
C9205 output50/a_27_47# net52 0
C9206 net50 output52/a_27_47# 0.00126f
C9207 _0982_/a_1059_315# acc0.A\[15\] 0
C9208 _0734_/a_285_47# _0317_ 0
C9209 clknet_1_1__leaf__0464_ _1044_/a_193_47# 0.10671f
C9210 _1011_/a_193_47# _0707_/a_75_199# 0
C9211 _1045_/a_193_47# _0202_ 0
C9212 VPWR hold61/a_391_47# 0.18911f
C9213 net175 _0465_ 0.00504f
C9214 _0346_ clknet_1_1__leaf__0465_ 0.02501f
C9215 _0164_ _0161_ 0
C9216 clknet_1_1__leaf__0460_ _0358_ 0.0013f
C9217 _0093_ _0404_ 0
C9218 _0413_ _0345_ 0.00301f
C9219 net131 clknet_1_1__leaf__0464_ 0.1199f
C9220 _1021_/a_193_47# net118 0
C9221 _1036_/a_27_47# comp0.B\[4\] 0.00105f
C9222 _1036_/a_466_413# net161 0.00391f
C9223 _0466_ _1064_/a_27_47# 0
C9224 control0.sh _0214_ 0
C9225 net59 net209 0.00382f
C9226 net10 _1042_/a_1059_315# 0
C9227 acc0.A\[2\] net175 0.03668f
C9228 _0229_ hold66/a_391_47# 0
C9229 _0107_ hold77/a_49_47# 0
C9230 _0153_ _0988_/a_466_413# 0
C9231 _0459_ _0114_ 0.00273f
C9232 _0248_ _0391_ 0
C9233 hold76/a_391_47# VPWR 0.17792f
C9234 _0372_ net223 0
C9235 _1057_/a_193_47# _0511_/a_81_21# 0
C9236 _1057_/a_27_47# _0511_/a_299_297# 0
C9237 _0767_/a_59_75# _0310_ 0.01892f
C9238 VPWR _1040_/a_381_47# 0.07435f
C9239 _0992_/a_466_413# clknet_1_1__leaf__0465_ 0
C9240 hold27/a_391_47# _0159_ 0
C9241 _0218_ _0583_/a_109_297# 0
C9242 _0294_ _0583_/a_109_47# 0.00243f
C9243 A[12] net181 0.00225f
C9244 hold31/a_285_47# clkbuf_1_1__f__0458_/a_110_47# 0.00142f
C9245 pp[10] _0155_ 0
C9246 _0743_/a_51_297# _0743_/a_245_297# 0.01218f
C9247 hold38/a_391_47# _0161_ 0
C9248 _1011_/a_891_413# _0334_ 0
C9249 _0483_ net167 0.07873f
C9250 _0163_ _1062_/a_1017_47# 0
C9251 _1058_/a_1017_47# net4 0
C9252 hold28/a_49_47# _0530_/a_81_21# 0.01564f
C9253 net223 hold40/a_49_47# 0
C9254 _0511_/a_384_47# _0286_ 0
C9255 _0451_ acc0.A\[15\] 0.03144f
C9256 _0725_/a_80_21# _0219_ 0
C9257 _0571_/a_27_297# _0571_/a_109_297# 0.17136f
C9258 _1032_/a_193_47# _1067_/a_891_413# 0
C9259 _0195_ hold71/a_391_47# 0.01205f
C9260 _1032_/a_466_413# _1067_/a_466_413# 0
C9261 _1032_/a_891_413# _1067_/a_193_47# 0
C9262 net36 _0399_ 0.05433f
C9263 _0646_/a_285_47# _0093_ 0
C9264 _0476_ net186 0
C9265 control0.state\[2\] _0160_ 0
C9266 net221 clknet_1_1__leaf__0461_ 0.0595f
C9267 _0999_/a_634_159# _0218_ 0.04525f
C9268 _1012_/a_592_47# net239 0
C9269 _1054_/a_1059_315# _0252_ 0
C9270 _0856_/a_79_21# acc0.A\[1\] 0.05216f
C9271 _0618_/a_510_47# net51 0
C9272 _0126_ hold8/a_49_47# 0
C9273 _0728_/a_59_75# _0725_/a_80_21# 0.00147f
C9274 _1057_/a_1017_47# net189 0
C9275 clkbuf_1_1__f__0463_/a_110_47# _1033_/a_381_47# 0
C9276 _0305_ _0245_ 0
C9277 clknet_1_0__leaf__0464_ _1049_/a_466_413# 0.00175f
C9278 net133 _1049_/a_193_47# 0
C9279 _0257_ VPWR 0.96285f
C9280 hold41/a_49_47# A[10] 0.00149f
C9281 clkbuf_0__0463_/a_110_47# net247 0
C9282 _1058_/a_634_159# acc0.A\[11\] 0
C9283 _0984_/a_466_413# net77 0
C9284 net70 _0991_/a_466_413# 0
C9285 _0457_ _0565_/a_240_47# 0.00146f
C9286 input2/a_75_212# _0510_/a_27_297# 0
C9287 VPWR _1035_/a_193_47# 0.31194f
C9288 _1053_/a_193_47# _1052_/a_381_47# 0
C9289 _1053_/a_381_47# _1052_/a_193_47# 0
C9290 _0550_/a_240_47# _1040_/a_193_47# 0
C9291 _0550_/a_149_47# _1040_/a_634_159# 0
C9292 hold22/a_285_47# _0437_ 0
C9293 _0298_ _0299_ 0.4192f
C9294 _0224_ hold4/a_285_47# 0.00238f
C9295 _0260_ _0268_ 0.26131f
C9296 _0789_/a_544_297# _0219_ 0
C9297 _0754_/a_512_297# _0345_ 0
C9298 _0467_ _1033_/a_27_47# 0
C9299 _0754_/a_51_297# _0377_ 0.09866f
C9300 _0982_/a_27_47# _0181_ 0.10978f
C9301 control0.sh _0207_ 0.0199f
C9302 _0330_ clknet_0__0462_ 0
C9303 _0179_ _1053_/a_27_47# 0
C9304 _0992_/a_27_47# _0283_ 0
C9305 hold37/a_285_47# _0142_ 0
C9306 net24 _0175_ 0.26544f
C9307 _1034_/a_193_47# net27 0
C9308 _0404_ _0304_ 0
C9309 _0452_ _0346_ 0.02795f
C9310 _0313_ _0321_ 0.14927f
C9311 _1064_/a_27_47# _1064_/a_193_47# 0.96976f
C9312 _1055_/a_592_47# clknet_1_1__leaf__0465_ 0
C9313 _0191_ net12 0
C9314 _0181_ _0145_ 0.00188f
C9315 _0837_/a_81_21# _0270_ 0.00123f
C9316 net44 _0778_/a_150_297# 0.00189f
C9317 _0387_ _0240_ 0.04106f
C9318 _0313_ clkbuf_0__0460_/a_110_47# 0.00123f
C9319 _0340_ _0342_ 0.22374f
C9320 _0508_/a_384_47# acc0.A\[15\] 0
C9321 clk input1/a_27_47# 0
C9322 clk _1068_/a_193_47# 0
C9323 _1018_/a_27_47# _1017_/a_27_47# 0.00133f
C9324 _0387_ _0369_ 0.13201f
C9325 VPWR clknet_1_1__leaf__0462_ 3.5699f
C9326 clknet_0__0457_ hold71/a_285_47# 0.00169f
C9327 _1038_/a_1059_315# net171 0.00707f
C9328 _1038_/a_466_413# _0207_ 0
C9329 _1026_/a_193_47# _1025_/a_27_47# 0
C9330 _1026_/a_27_47# _1025_/a_193_47# 0
C9331 VPWR _0818_/a_109_47# 0
C9332 _0587_/a_27_47# hold92/a_49_47# 0
C9333 _0829_/a_109_297# _0434_ 0
C9334 _1051_/a_27_47# net148 0
C9335 _1051_/a_381_47# _0524_/a_27_297# 0
C9336 net1 _1063_/a_27_47# 0
C9337 _0748_/a_299_297# _0250_ 0
C9338 clkload3/Y _0459_ 0.00301f
C9339 _1033_/a_27_47# comp0.B\[0\] 0.02648f
C9340 _1053_/a_381_47# net12 0.01551f
C9341 _0181_ net17 0.02535f
C9342 _0535_/a_68_297# hold6/a_49_47# 0.00521f
C9343 _0181_ net238 0
C9344 _0197_ _0186_ 0.07126f
C9345 control0.state\[1\] net232 0.00253f
C9346 VPWR _0994_/a_381_47# 0.07542f
C9347 _0343_ _1060_/a_466_413# 0.00126f
C9348 _0359_ net112 0.00202f
C9349 net159 _1068_/a_634_159# 0.00124f
C9350 clk _0478_ 0
C9351 net45 clkload4/Y 0
C9352 clknet_1_0__leaf__0458_ _0854_/a_79_21# 0.00284f
C9353 _0179_ _0451_ 0
C9354 _0359_ acc0.A\[24\] 0
C9355 _0461_ _1015_/a_381_47# 0.00927f
C9356 _1010_/a_1059_315# _0350_ 0.03866f
C9357 _0557_/a_512_297# clknet_1_1__leaf__0463_ 0
C9358 pp[27] _1011_/a_1059_315# 0
C9359 _0181_ _0446_ 0
C9360 _0737_/a_35_297# _0737_/a_285_47# 0.00723f
C9361 hold13/a_285_47# _1034_/a_1059_315# 0
C9362 input2/a_75_212# _0181_ 0.0115f
C9363 _0259_ _0990_/a_193_47# 0.00116f
C9364 net45 _0582_/a_373_47# 0
C9365 _1039_/a_1059_315# control0.sh 0
C9366 _0565_/a_245_297# _0173_ 0
C9367 _0287_ _0809_/a_299_297# 0.00644f
C9368 _0289_ _0809_/a_384_47# 0
C9369 _0341_ _1013_/a_1017_47# 0
C9370 _0663_/a_297_47# _0369_ 0
C9371 net61 _0272_ 0
C9372 net157 _1061_/a_1059_315# 0.01464f
C9373 hold87/a_391_47# _0216_ 0
C9374 _0961_/a_199_47# control0.count\[0\] 0
C9375 _0699_/a_150_297# _0329_ 0
C9376 _0846_/a_512_297# _0350_ 0
C9377 _0454_ acc0.A\[1\] 0
C9378 _0369_ _0382_ 0.24199f
C9379 _0383_ _0237_ 0.04326f
C9380 _0995_/a_1059_315# _0219_ 0
C9381 _0227_ _0618_/a_79_21# 0.00113f
C9382 comp0.B\[4\] comp0.B\[3\] 0.07407f
C9383 _0192_ _0179_ 0.09018f
C9384 _0695_/a_472_297# _0312_ 0.00307f
C9385 _0695_/a_80_21# _0323_ 0.16009f
C9386 _1009_/a_891_413# _0350_ 0
C9387 _1034_/a_193_47# _1033_/a_193_47# 0.00464f
C9388 net247 hold71/a_49_47# 0.04371f
C9389 _0183_ _1016_/a_27_47# 0.00157f
C9390 net108 acc0.A\[22\] 0.01029f
C9391 comp0.B\[10\] _0204_ 0.06389f
C9392 _1031_/a_466_413# _1031_/a_561_413# 0.00772f
C9393 _1031_/a_634_159# _1031_/a_975_413# 0
C9394 _0531_/a_109_297# _1047_/a_634_159# 0
C9395 _0531_/a_27_297# _1047_/a_466_413# 0
C9396 _0174_ hold6/a_49_47# 0.01478f
C9397 net63 A[8] 0
C9398 net200 net112 0
C9399 _0153_ _0186_ 0
C9400 net67 hold70/a_285_47# 0.05662f
C9401 hold30/a_391_47# _0756_/a_47_47# 0.00139f
C9402 _1041_/a_193_47# VPWR 0.28576f
C9403 B[8] _0139_ 0
C9404 net65 _0829_/a_27_47# 0
C9405 comp0.B\[10\] hold6/a_391_47# 0
C9406 pp[15] _0995_/a_27_47# 0.00481f
C9407 _0722_/a_215_47# _0722_/a_510_47# 0.00529f
C9408 _0645_/a_47_47# acc0.A\[14\] 0.05765f
C9409 net200 acc0.A\[24\] 0.00183f
C9410 _1005_/a_891_413# net91 0
C9411 _1005_/a_1059_315# _0103_ 0.0671f
C9412 _0179_ _0508_/a_384_47# 0
C9413 _0465_ _0842_/a_145_75# 0
C9414 _0331_ _0589_/a_113_47# 0
C9415 _0386_ _0247_ 0
C9416 _0130_ _0183_ 0
C9417 _0325_ _0366_ 0
C9418 comp0.B\[6\] net26 0
C9419 VPWR net242 0.3372f
C9420 net70 net222 0
C9421 acc0.A\[12\] net41 0
C9422 acc0.A\[21\] _0181_ 0
C9423 _1060_/a_634_159# net5 0
C9424 _1060_/a_27_47# _0185_ 0
C9425 _1013_/a_891_413# _1013_/a_1017_47# 0.00617f
C9426 _0976_/a_76_199# _1069_/a_1059_315# 0.01104f
C9427 net58 _0842_/a_59_75# 0.00506f
C9428 net1 _1062_/a_1059_315# 0
C9429 _1002_/a_634_159# _1002_/a_592_47# 0
C9430 VPWR net11 0.49202f
C9431 _1027_/a_27_47# _0365_ 0
C9432 _0429_ VPWR 0.71191f
C9433 _1059_/a_27_47# _0302_ 0
C9434 _0227_ _0486_ 0
C9435 _0319_ _0687_/a_145_75# 0.00198f
C9436 _0758_/a_215_47# _0379_ 0.05119f
C9437 _0640_/a_392_297# VPWR 0
C9438 net63 _0837_/a_585_47# 0
C9439 net45 clknet_1_0__leaf__0461_ 0.00532f
C9440 net22 _1046_/a_891_413# 0
C9441 _0679_/a_68_297# _0392_ 0
C9442 _0144_ clknet_1_1__leaf__0457_ 0
C9443 _0749_/a_81_21# _0352_ 0
C9444 _0965_/a_285_47# clknet_1_0__leaf_clk 0.03297f
C9445 hold28/a_391_47# _1049_/a_193_47# 0
C9446 acc0.A\[18\] _0611_/a_150_297# 0
C9447 _0552_/a_150_297# _0173_ 0
C9448 hold87/a_391_47# _0852_/a_285_297# 0
C9449 _0361_ _0105_ 0
C9450 VPWR _0997_/a_561_413# 0.00232f
C9451 _0678_/a_68_297# _0352_ 0
C9452 _0836_/a_68_297# _0255_ 0
C9453 _0409_ _0405_ 0.19375f
C9454 _1038_/a_193_47# net174 0
C9455 output58/a_27_47# _0274_ 0
C9456 _0662_/a_81_21# _0785_/a_81_21# 0
C9457 _1059_/a_891_413# _0369_ 0.01291f
C9458 _0766_/a_109_297# _0352_ 0
C9459 net149 acc0.A\[19\] 0.15876f
C9460 net54 hold8/a_49_47# 0.01971f
C9461 acc0.A\[12\] A[11] 0.00248f
C9462 _0154_ net181 0.00665f
C9463 _1041_/a_27_47# _0550_/a_51_297# 0
C9464 _0664_/a_382_297# clknet_1_1__leaf__0459_ 0
C9465 _0765_/a_215_47# _0385_ 0.00761f
C9466 _1035_/a_381_47# _0175_ 0.00487f
C9467 _0753_/a_561_47# net51 0
C9468 pp[28] _1011_/a_466_413# 0
C9469 input23/a_75_212# _0175_ 0
C9470 VPWR _1061_/a_592_47# 0
C9471 _0089_ acc0.A\[9\] 0.00335f
C9472 clknet_1_0__leaf__0463_ _1046_/a_891_413# 0
C9473 _0837_/a_81_21# _1051_/a_27_47# 0
C9474 net82 net5 0.14044f
C9475 _0398_ _0306_ 0
C9476 _0399_ _0308_ 0
C9477 output44/a_27_47# _0705_/a_59_75# 0
C9478 VPWR _0668_/a_382_297# 0.00516f
C9479 _1034_/a_1059_315# _0132_ 0
C9480 _0971_/a_299_297# _0487_ 0.06336f
C9481 net89 control0.count\[3\] 0
C9482 _0241_ _0242_ 0.2906f
C9483 _0217_ _0116_ 0.18443f
C9484 _0176_ _0548_/a_512_297# 0
C9485 _0363_ net52 0
C9486 VPWR hold7/a_391_47# 0.17532f
C9487 _1000_/a_27_47# _0393_ 0.15144f
C9488 net117 acc0.A\[30\] 0.10689f
C9489 output38/a_27_47# net246 0
C9490 _0343_ _0796_/a_215_47# 0.00327f
C9491 acc0.A\[17\] _0115_ 0
C9492 hold31/a_391_47# acc0.A\[8\] 0.0019f
C9493 net104 _0459_ 0.00135f
C9494 hold10/a_391_47# _0924_/a_27_47# 0
C9495 acc0.A\[12\] _0744_/a_27_47# 0
C9496 clknet_1_0__leaf__0458_ _1014_/a_193_47# 0
C9497 _0975_/a_59_75# _0162_ 0.00491f
C9498 _0327_ _0353_ 0
C9499 _0168_ _1069_/a_1017_47# 0
C9500 _1018_/a_466_413# _0218_ 0
C9501 _0212_ _1066_/a_466_413# 0
C9502 _1030_/a_634_159# _0336_ 0
C9503 _0990_/a_27_47# _0186_ 0
C9504 hold30/a_49_47# net110 0
C9505 _0312_ _0743_/a_240_47# 0
C9506 _0695_/a_80_21# net237 0
C9507 _1011_/a_561_413# net57 0
C9508 _1017_/a_27_47# clknet_1_1__leaf__0461_ 0
C9509 _1000_/a_466_413# _0245_ 0.00103f
C9510 _1000_/a_193_47# _0246_ 0
C9511 pp[22] acc0.A\[23\] 0.00164f
C9512 _0572_/a_27_297# _0572_/a_109_47# 0.00393f
C9513 _0133_ comp0.B\[2\] 0.01606f
C9514 _0601_/a_150_297# _0219_ 0
C9515 _0276_ hold91/a_285_47# 0
C9516 _1006_/a_1059_315# _1006_/a_1017_47# 0
C9517 _1006_/a_193_47# net92 0.0042f
C9518 _0656_/a_145_75# acc0.A\[9\] 0
C9519 _0993_/a_1059_315# net246 0.0061f
C9520 init input26/a_75_212# 0.00376f
C9521 input33/a_75_212# B[3] 0
C9522 output59/a_27_47# _0340_ 0
C9523 pp[30] _0710_/a_109_47# 0
C9524 clknet_1_0__leaf__0460_ _0754_/a_149_47# 0
C9525 _0695_/a_300_47# _0219_ 0.00121f
C9526 _0984_/a_634_159# _0984_/a_592_47# 0
C9527 _0579_/a_27_297# _0891_/a_27_47# 0
C9528 net8 _0492_/a_27_47# 0
C9529 _0195_ acc0.A\[25\] 0.00404f
C9530 _0808_/a_81_21# _0091_ 0.08791f
C9531 _0438_ _0988_/a_634_159# 0
C9532 net79 _0417_ 0.00892f
C9533 acc0.A\[9\] _0986_/a_891_413# 0
C9534 input11/a_75_212# net12 0
C9535 _0664_/a_79_21# _0289_ 0
C9536 _0550_/a_240_47# _0207_ 0
C9537 hold97/a_391_47# _0365_ 0
C9538 comp0.B\[6\] hold84/a_285_47# 0
C9539 net35 _0166_ 0
C9540 _1039_/a_592_47# VPWR 0
C9541 _0730_/a_297_297# VPWR 0.01098f
C9542 hold78/a_391_47# _1031_/a_193_47# 0
C9543 net34 net226 0
C9544 _0986_/a_1059_315# _0986_/a_1017_47# 0
C9545 net168 _1054_/a_193_47# 0.06941f
C9546 net148 _0085_ 0.00143f
C9547 _1056_/a_27_47# _0186_ 0.00715f
C9548 VPWR hold92/a_49_47# 0.30946f
C9549 _1023_/a_466_413# net177 0.02296f
C9550 _1023_/a_1059_315# net109 0
C9551 hold43/a_285_47# acc0.A\[29\] 0
C9552 _1023_/a_27_47# acc0.A\[23\] 0
C9553 _1037_/a_466_413# _0175_ 0.00292f
C9554 _0369_ _1006_/a_27_47# 0
C9555 net248 _0432_ 0.00121f
C9556 _0512_/a_27_297# acc0.A\[10\] 0.00158f
C9557 hold25/a_391_47# _0176_ 0.01852f
C9558 hold32/a_49_47# A[10] 0
C9559 _1042_/a_381_47# net128 0
C9560 _0094_ _0507_/a_27_297# 0
C9561 _0753_/a_297_297# _0227_ 0
C9562 _0684_/a_59_75# _0733_/a_448_47# 0
C9563 _1044_/a_27_47# _0202_ 0
C9564 net104 _0265_ 0
C9565 _0337_ _0723_/a_207_413# 0
C9566 _0697_/a_80_21# _0686_/a_219_297# 0
C9567 net23 _0584_/a_373_47# 0
C9568 hold58/a_285_47# clknet_1_1__leaf__0463_ 0.01841f
C9569 _0195_ _0571_/a_27_297# 0.1343f
C9570 net34 _0946_/a_112_297# 0.00234f
C9571 _0691_/a_68_297# _0359_ 0
C9572 _1011_/a_27_47# _0339_ 0
C9573 output55/a_27_47# pp[27] 0.15389f
C9574 _0675_/a_68_297# net219 0
C9575 _1037_/a_1059_315# control0.sh 0.01841f
C9576 _0439_ clknet_1_1__leaf__0458_ 0.02857f
C9577 hold55/a_285_47# _0181_ 0.03562f
C9578 _0763_/a_193_47# _0384_ 0.01172f
C9579 output56/a_27_47# _0334_ 0
C9580 VPWR clknet_1_1__leaf__0458_ 3.71431f
C9581 _0218_ acc0.A\[13\] 0.34642f
C9582 clkbuf_1_0__f__0463_/a_110_47# _0548_/a_51_297# 0
C9583 net163 _1031_/a_193_47# 0.24592f
C9584 _0195_ _0148_ 0
C9585 net133 _0531_/a_373_47# 0
C9586 _0129_ _1031_/a_466_413# 0
C9587 hold36/a_49_47# clkbuf_0__0464_/a_110_47# 0.01705f
C9588 _0183_ _0534_/a_81_21# 0
C9589 _0341_ _0216_ 0.03432f
C9590 _0128_ hold61/a_49_47# 0
C9591 net64 hold31/a_391_47# 0.05857f
C9592 _0430_ hold31/a_49_47# 0
C9593 _1059_/a_466_413# net229 0.02419f
C9594 _0457_ _0171_ 0
C9595 _0578_/a_27_297# _1067_/a_1059_315# 0
C9596 hold22/a_285_47# _0252_ 0
C9597 hold31/a_285_47# _0621_/a_285_297# 0.00234f
C9598 clkbuf_1_1__f_clk/a_110_47# clknet_1_0__leaf__0461_ 0.0113f
C9599 hold42/a_285_47# _0156_ 0.01335f
C9600 _1057_/a_1059_315# _0156_ 0.01173f
C9601 _0257_ _0835_/a_493_297# 0.00122f
C9602 _0274_ clkbuf_1_0__f__0465_/a_110_47# 0
C9603 _0486_ _0477_ 0
C9604 acc0.A\[12\] net66 0
C9605 clkbuf_0__0457_/a_110_47# hold40/a_49_47# 0
C9606 _0997_/a_466_413# _0095_ 0
C9607 _0556_/a_68_297# clknet_1_1__leaf__0463_ 0.00207f
C9608 _0574_/a_109_297# net110 0
C9609 hold99/a_285_47# net246 0.01139f
C9610 net234 net47 0.02259f
C9611 _0456_ _0633_/a_109_297# 0
C9612 _0347_ _0738_/a_150_297# 0
C9613 _0165_ _0181_ 0.02598f
C9614 _0852_/a_285_297# _0264_ 0.0225f
C9615 hold24/a_285_47# _0176_ 0
C9616 _0228_ clknet_1_0__leaf__0460_ 0.39402f
C9617 _0275_ _0347_ 0
C9618 clknet_1_0__leaf__0457_ _0526_/a_27_47# 0
C9619 net161 net26 0
C9620 _1053_/a_27_47# hold83/a_49_47# 0.00835f
C9621 _0837_/a_266_47# clkbuf_1_0__f__0465_/a_110_47# 0
C9622 _0579_/a_27_297# _0346_ 0.00408f
C9623 _0458_ clknet_1_1__leaf__0457_ 0.00348f
C9624 _0530_/a_81_21# clkbuf_1_0__f__0464_/a_110_47# 0
C9625 net42 net41 1.19259f
C9626 _0100_ _0765_/a_215_47# 0
C9627 _0146_ net10 0
C9628 _1065_/a_27_47# _1065_/a_466_413# 0.26005f
C9629 _1065_/a_193_47# _1065_/a_634_159# 0.11072f
C9630 net140 net154 0
C9631 net232 _1066_/a_634_159# 0
C9632 hold30/a_285_47# _0120_ 0.00632f
C9633 _0121_ _0217_ 0.25657f
C9634 _0787_/a_209_297# _0281_ 0.04094f
C9635 _0571_/a_109_297# _0125_ 0.00169f
C9636 _0428_ _0516_/a_27_297# 0
C9637 _0107_ _0308_ 0
C9638 _1036_/a_27_47# _1035_/a_193_47# 0
C9639 _1036_/a_193_47# _1035_/a_27_47# 0
C9640 _0584_/a_109_297# clknet_1_0__leaf__0461_ 0.0235f
C9641 _0532_/a_81_21# _0198_ 0.18163f
C9642 VPWR _0263_ 0.82433f
C9643 _0216_ _0722_/a_79_21# 0
C9644 clkload4/Y VPWR 0.42509f
C9645 _1033_/a_891_413# _0565_/a_51_297# 0.00145f
C9646 _0954_/a_32_297# _1042_/a_193_47# 0
C9647 _0954_/a_114_297# _1042_/a_27_47# 0
C9648 _0311_ _0347_ 0
C9649 net85 _0218_ 0.25466f
C9650 hold17/a_49_47# clknet_1_0__leaf_clk 0
C9651 VPWR _1047_/a_27_47# 0.6568f
C9652 _0811_/a_81_21# _0811_/a_299_297# 0.08213f
C9653 _0343_ _0833_/a_79_21# 0
C9654 _0195_ _1013_/a_561_413# 0
C9655 VPWR _0957_/a_220_297# 0.00426f
C9656 _0236_ _0248_ 0.19677f
C9657 _0843_/a_68_297# _0345_ 0
C9658 clkbuf_1_1__f__0463_/a_110_47# comp0.B\[1\] 0
C9659 clknet_0__0463_ _0131_ 0.0191f
C9660 clknet_1_0__leaf__0464_ _0147_ 0.01144f
C9661 _0139_ clknet_1_1__leaf__0464_ 0
C9662 _0332_ hold95/a_285_47# 0
C9663 hold101/a_49_47# hold101/a_285_47# 0.22264f
C9664 net173 _0205_ 0
C9665 VPWR _0582_/a_373_47# 0
C9666 net144 acc0.A\[11\] 0.41722f
C9667 net70 _0089_ 0
C9668 net247 _0264_ 0
C9669 clknet_0__0457_ clknet_1_0__leaf__0458_ 0.01504f
C9670 VPWR _1007_/a_466_413# 0.26458f
C9671 _0399_ _0989_/a_634_159# 0.00859f
C9672 _0172_ _1040_/a_891_413# 0
C9673 _0137_ _1040_/a_466_413# 0
C9674 net30 _1040_/a_381_47# 0
C9675 _1058_/a_891_413# VPWR 0.18657f
C9676 hold34/a_391_47# _0514_/a_27_297# 0
C9677 _0179_ _1051_/a_634_159# 0.01313f
C9678 _0710_/a_109_47# _0339_ 0
C9679 _0377_ _0219_ 0.003f
C9680 _0534_/a_81_21# acc0.A\[15\] 0.0503f
C9681 clknet_0__0465_ _0817_/a_81_21# 0
C9682 _0261_ _0630_/a_109_297# 0
C9683 _0178_ _1049_/a_27_47# 0
C9684 clkbuf_1_1__f__0460_/a_110_47# _0350_ 0.00218f
C9685 _1064_/a_466_413# _1064_/a_592_47# 0.00553f
C9686 _1064_/a_634_159# _1064_/a_1017_47# 0
C9687 _0272_ _0431_ 0
C9688 hold78/a_285_47# _0345_ 0
C9689 clknet_1_0__leaf__0458_ _0852_/a_117_297# 0
C9690 _0442_ _0256_ 0
C9691 _0441_ _0271_ 0
C9692 _0376_ _0750_/a_27_47# 0
C9693 _1015_/a_891_413# net23 0.00648f
C9694 clknet_1_1__leaf__0459_ _0402_ 0.05718f
C9695 pp[15] _0299_ 0.00126f
C9696 clknet_1_1__leaf_clk _1063_/a_1059_315# 0
C9697 _0827_/a_27_47# _0434_ 0.0394f
C9698 net172 _0207_ 0
C9699 _0707_/a_315_47# _0334_ 0
C9700 _0837_/a_81_21# _0085_ 0.08934f
C9701 _0346_ _0277_ 0.02052f
C9702 VPWR hold80/a_49_47# 0.29509f
C9703 _0475_ _0171_ 0
C9704 _0325_ acc0.A\[24\] 0.0904f
C9705 comp0.B\[14\] net18 0
C9706 _0243_ _1001_/a_27_47# 0
C9707 _0388_ _0310_ 0.15564f
C9708 _0260_ _0443_ 0
C9709 clkbuf_1_0__f__0459_/a_110_47# _1060_/a_466_413# 0.00605f
C9710 _0959_/a_80_21# clknet_1_1__leaf_clk 0.00115f
C9711 _0149_ _0524_/a_373_47# 0
C9712 _0428_ _0399_ 0.37682f
C9713 _1002_/a_1059_315# _0369_ 0.02088f
C9714 _0192_ hold83/a_49_47# 0
C9715 acc0.A\[16\] _0240_ 0
C9716 net245 _0218_ 0.01551f
C9717 acc0.A\[16\] _0369_ 0.44294f
C9718 net220 _0384_ 0
C9719 net1 net149 0.01444f
C9720 _0680_/a_80_21# _0370_ 0
C9721 net200 net111 0.0356f
C9722 _0692_/a_113_47# _0352_ 0
C9723 _0343_ _0158_ 0
C9724 control0.state\[0\] _0967_/a_403_297# 0.00188f
C9725 net34 _0967_/a_215_297# 0
C9726 control0.state\[1\] _0967_/a_297_297# 0.00176f
C9727 _0399_ hold60/a_391_47# 0.06624f
C9728 control0.state\[1\] _0162_ 0
C9729 _0229_ _0374_ 0.01641f
C9730 done VPWR 0.21694f
C9731 _0985_/a_193_47# net61 0
C9732 _1013_/a_193_47# _0339_ 0
C9733 _0596_/a_145_75# _0222_ 0
C9734 acc0.A\[12\] net80 0
C9735 _0701_/a_303_47# _0347_ 0
C9736 _0701_/a_80_21# _0352_ 0
C9737 clknet_0__0465_ _0084_ 0.00446f
C9738 _0804_/a_79_21# _0647_/a_47_47# 0
C9739 _1017_/a_891_413# acc0.A\[17\] 0.0026f
C9740 _0664_/a_297_47# _0281_ 0.06294f
C9741 _0259_ clknet_1_1__leaf__0465_ 0.00119f
C9742 input11/a_75_212# pp[5] 0
C9743 _0251_ acc0.A\[6\] 0.02927f
C9744 _0134_ clknet_1_1__leaf__0463_ 0.00965f
C9745 output55/a_27_47# _0216_ 0
C9746 _1008_/a_1059_315# _0345_ 0
C9747 hold16/a_391_47# _0219_ 0
C9748 _0854_/a_79_21# _0455_ 0.0776f
C9749 _0963_/a_285_297# _1070_/a_1059_315# 0
C9750 VPWR clknet_1_0__leaf__0461_ 3.69811f
C9751 _0350_ _0445_ 0
C9752 _0313_ _1026_/a_27_47# 0
C9753 net201 _0208_ 0.25011f
C9754 _0836_/a_68_297# _0830_/a_215_47# 0
C9755 hold74/a_285_47# _1016_/a_1059_315# 0.0054f
C9756 hold56/a_391_47# clkbuf_1_1__f__0463_/a_110_47# 0.00112f
C9757 clkbuf_1_1__f_clk/a_110_47# _1063_/a_891_413# 0.00187f
C9758 control0.reset _0494_/a_27_47# 0
C9759 _0153_ net62 0
C9760 _0593_/a_113_47# net51 0
C9761 _0346_ _0808_/a_81_21# 0.12696f
C9762 _0999_/a_193_47# _0347_ 0.00193f
C9763 net198 _0543_/a_150_297# 0
C9764 net18 _0543_/a_68_297# 0
C9765 _0413_ _0997_/a_193_47# 0
C9766 hold78/a_285_47# hold16/a_49_47# 0
C9767 hold63/a_391_47# net112 0
C9768 hold36/a_285_47# _0143_ 0.05443f
C9769 _0498_/a_51_297# _0498_/a_512_297# 0.0116f
C9770 _0830_/a_215_47# net212 0.06338f
C9771 _1015_/a_466_413# clknet_1_0__leaf__0461_ 0
C9772 _0180_ _0159_ 0
C9773 _0461_ acc0.A\[18\] 0.02269f
C9774 clknet_1_0__leaf__0462_ _0374_ 0
C9775 net1 _0958_/a_197_47# 0.00197f
C9776 clknet_1_0__leaf__0465_ _1052_/a_561_413# 0
C9777 _0275_ clkbuf_0__0465_/a_110_47# 0
C9778 _1038_/a_1059_315# _0553_/a_51_297# 0.00126f
C9779 _1038_/a_27_47# _0553_/a_240_47# 0
C9780 _1034_/a_27_47# net119 0.00173f
C9781 _0195_ _0532_/a_384_47# 0
C9782 _0557_/a_51_297# _0557_/a_240_47# 0.03076f
C9783 _1037_/a_592_47# VPWR 0
C9784 _0577_/a_27_297# _1005_/a_193_47# 0
C9785 _0440_ acc0.A\[4\] 0
C9786 _0531_/a_27_297# _0145_ 0
C9787 _0514_/a_27_297# _0181_ 0.16997f
C9788 acc0.A\[7\] _0827_/a_27_47# 0
C9789 _0179_ clknet_1_0__leaf__0465_ 0.26506f
C9790 _0175_ _1062_/a_466_413# 0
C9791 _0715_/a_27_47# _0399_ 0
C9792 _0682_/a_68_297# _0347_ 0
C9793 _0361_ _0359_ 0
C9794 net40 A[13] 0.06903f
C9795 _0643_/a_253_47# _0350_ 0
C9796 clknet_1_0__leaf__0458_ _0844_/a_79_21# 0
C9797 hold23/a_391_47# _0179_ 0
C9798 _0489_ _0976_/a_218_47# 0
C9799 _1022_/a_381_47# _1005_/a_1059_315# 0
C9800 net45 _0218_ 0.44067f
C9801 hold51/a_49_47# hold51/a_285_47# 0.22264f
C9802 net46 _0609_/a_109_297# 0.00245f
C9803 net58 acc0.A\[6\] 0.09687f
C9804 _0800_/a_240_47# _0668_/a_79_21# 0
C9805 hold12/a_285_47# clknet_1_0__leaf__0460_ 0.00166f
C9806 _0983_/a_381_47# clknet_1_0__leaf__0461_ 0
C9807 net11 _0523_/a_81_21# 0.01968f
C9808 comp0.B\[7\] net8 0.0333f
C9809 _0438_ _0253_ 0.00748f
C9810 net26 hold84/a_285_47# 0
C9811 _0512_/a_109_297# _0181_ 0.01052f
C9812 _0482_ control0.state\[2\] 0
C9813 _1008_/a_27_47# _1008_/a_634_159# 0.14145f
C9814 _0815_/a_199_47# _0084_ 0
C9815 _0466_ _1069_/a_466_413# 0
C9816 _0488_ _1069_/a_1059_315# 0
C9817 _1021_/a_381_47# clknet_1_1__leaf_clk 0
C9818 _1054_/a_1017_47# clknet_1_1__leaf__0458_ 0
C9819 hold16/a_285_47# _0129_ 0.00763f
C9820 pp[27] _0707_/a_208_47# 0
C9821 clknet_1_0__leaf__0463_ input30/a_75_212# 0.01854f
C9822 net40 _0279_ 0
C9823 _1002_/a_592_47# net88 0.00107f
C9824 _1020_/a_466_413# _1020_/a_381_47# 0.03733f
C9825 _1020_/a_193_47# _1020_/a_975_413# 0
C9826 _1020_/a_1059_315# _1020_/a_891_413# 0.31086f
C9827 _1002_/a_975_413# _0100_ 0
C9828 hold18/a_285_47# hold18/a_391_47# 0.41909f
C9829 _0243_ _0459_ 0.01674f
C9830 _0400_ acc0.A\[15\] 0.0256f
C9831 _1035_/a_193_47# comp0.B\[3\] 0
C9832 _0180_ _0447_ 0.00234f
C9833 _0343_ _0581_/a_27_297# 0
C9834 _0564_/a_68_297# _0173_ 0
C9835 clkbuf_1_0__f__0464_/a_110_47# _1049_/a_466_413# 0.0107f
C9836 _0343_ acc0.A\[14\] 0.0282f
C9837 _0305_ _0326_ 0
C9838 _0747_/a_79_21# clknet_0__0460_ 0.00173f
C9839 hold28/a_49_47# _0147_ 0.00446f
C9840 _0298_ _0346_ 0
C9841 _0983_/a_561_413# net47 0.00247f
C9842 acc0.A\[22\] _0350_ 0
C9843 _0217_ _0380_ 0
C9844 _0515_/a_81_21# _0515_/a_299_297# 0.08213f
C9845 clknet_1_1__leaf_clk _0173_ 0
C9846 control0.sh _0561_/a_240_47# 0
C9847 _0747_/a_510_47# _0250_ 0.00457f
C9848 _0188_ _0512_/a_27_297# 0.11374f
C9849 _0199_ _1048_/a_1059_315# 0.00143f
C9850 acc0.A\[20\] _0713_/a_27_47# 0
C9851 _1013_/a_634_159# net99 0
C9852 _1001_/a_592_47# net46 0
C9853 _0346_ _0296_ 0.25536f
C9854 _0554_/a_68_297# clknet_1_1__leaf__0463_ 0
C9855 _1041_/a_27_47# _0172_ 0.03156f
C9856 _1041_/a_193_47# net30 0
C9857 _0404_ _0997_/a_27_47# 0
C9858 _0222_ _0383_ 0
C9859 _0349_ hold95/a_391_47# 0.05f
C9860 _0388_ _0768_/a_27_47# 0.0517f
C9861 clkload4/Y clknet_1_0__leaf__0459_ 0.33696f
C9862 net227 hold80/a_285_47# 0.01139f
C9863 hold7/a_285_47# _0523_/a_299_297# 0
C9864 _0992_/a_27_47# _0345_ 0
C9865 _0533_/a_27_297# clkbuf_1_1__f__0457_/a_110_47# 0
C9866 _0645_/a_377_297# net41 0.00646f
C9867 _0285_ VPWR 1.36994f
C9868 _0390_ clknet_1_0__leaf__0461_ 0.00295f
C9869 _0472_ control0.sh 0.02862f
C9870 hold94/a_285_47# _0754_/a_149_47# 0
C9871 hold94/a_49_47# _0754_/a_240_47# 0
C9872 _0570_/a_27_297# _0347_ 0
C9873 _0826_/a_219_297# _0826_/a_301_297# 0.00516f
C9874 _0587_/a_27_47# _0218_ 0.26161f
C9875 pp[17] _0336_ 0
C9876 _0990_/a_27_47# net62 0.03811f
C9877 comp0.B\[2\] _0208_ 0.10271f
C9878 VPWR net133 0.51215f
C9879 _0982_/a_193_47# _0855_/a_81_21# 0.00297f
C9880 _1072_/a_466_413# _0468_ 0
C9881 net190 _0687_/a_59_75# 0.00133f
C9882 _0229_ _0249_ 0
C9883 hold42/a_49_47# _1058_/a_27_47# 0.01327f
C9884 _0275_ _0824_/a_59_75# 0
C9885 _0176_ _0138_ 0.001f
C9886 _0211_ _0176_ 0
C9887 _1058_/a_27_47# _1057_/a_466_413# 0
C9888 _1058_/a_193_47# _1057_/a_634_159# 0
C9889 _1058_/a_634_159# _1057_/a_193_47# 0
C9890 _1058_/a_466_413# _1057_/a_27_47# 0
C9891 _0413_ _0411_ 0.06974f
C9892 _0464_ _1061_/a_891_413# 0.00681f
C9893 clk VPWR 1.16227f
C9894 _0476_ control0.state\[2\] 0.17925f
C9895 B[9] hold5/a_49_47# 0.00849f
C9896 _0476_ net120 0
C9897 input20/a_75_212# net196 0
C9898 _0258_ _0399_ 0
C9899 _1000_/a_891_413# _0347_ 0
C9900 _1000_/a_634_159# _0352_ 0.03689f
C9901 VPWR _1063_/a_891_413# 0.19506f
C9902 _0996_/a_27_47# _1060_/a_1059_315# 0
C9903 _0285_ _0654_/a_27_413# 0.09474f
C9904 _1052_/a_1017_47# net73 0
C9905 _0369_ net91 0
C9906 _0098_ _0245_ 0.02208f
C9907 _0195_ net57 0.06953f
C9908 net210 _0195_ 0.09585f
C9909 VPWR _0959_/a_217_297# 0.18604f
C9910 hold60/a_49_47# _0345_ 0.00289f
C9911 VPWR _0585_/a_27_297# 0.22938f
C9912 _0328_ clkbuf_0__0462_/a_110_47# 0.13753f
C9913 _0453_ _0263_ 0
C9914 net190 hold9/a_391_47# 0.04694f
C9915 pp[8] pp[4] 0
C9916 _0272_ _0269_ 0.36653f
C9917 _1056_/a_27_47# net62 0
C9918 _0347_ hold50/a_49_47# 0.0027f
C9919 net211 _0461_ 0.03492f
C9920 _0111_ net42 0
C9921 _0236_ _0235_ 0.06367f
C9922 VPWR _1060_/a_891_413# 0.19978f
C9923 _0548_/a_51_297# _0548_/a_245_297# 0.01218f
C9924 _1019_/a_891_413# acc0.A\[19\] 0.00325f
C9925 pp[28] _0707_/a_544_297# 0.00121f
C9926 net220 _0383_ 0
C9927 _0856_/a_215_47# _0856_/a_510_47# 0.00529f
C9928 net208 net116 0.01014f
C9929 hold84/a_49_47# hold84/a_391_47# 0.00188f
C9930 VPWR _0988_/a_1017_47# 0
C9931 _0855_/a_299_297# _0446_ 0
C9932 _0659_/a_68_297# _0181_ 0
C9933 _0172_ hold7/a_285_47# 0
C9934 _1054_/a_381_47# _0186_ 0
C9935 VPWR comp0.B\[10\] 1.89883f
C9936 _0402_ _0655_/a_215_53# 0
C9937 _1000_/a_193_47# _0774_/a_68_297# 0
C9938 net157 _1047_/a_381_47# 0.01626f
C9939 clknet_0_clk _0974_/a_222_93# 0.00266f
C9940 clknet_1_0__leaf__0459_ clknet_1_0__leaf__0461_ 0.06993f
C9941 _0472_ net157 0
C9942 hold89/a_49_47# _0486_ 0.00768f
C9943 hold89/a_285_47# control0.state\[2\] 0.0937f
C9944 _0135_ _0175_ 0
C9945 _0619_/a_68_297# _0989_/a_634_159# 0
C9946 hold45/a_391_47# _0511_/a_299_297# 0
C9947 _0643_/a_103_199# _0443_ 0
C9948 net56 clknet_1_1__leaf__0462_ 0.90073f
C9949 pp[28] pp[29] 0.21044f
C9950 net219 _0242_ 0.09334f
C9951 net206 acc0.A\[19\] 0.06715f
C9952 _0369_ _0288_ 0
C9953 _0348_ _1011_/a_193_47# 0
C9954 _0094_ _0185_ 0
C9955 net55 _0361_ 0
C9956 _0704_/a_68_297# acc0.A\[30\] 0.21384f
C9957 _0766_/a_109_297# _0392_ 0.0033f
C9958 _1044_/a_975_413# net20 0
C9959 _0682_/a_68_297# _1025_/a_27_47# 0
C9960 pp[27] _1010_/a_634_159# 0
C9961 clknet_1_1__leaf__0458_ _0523_/a_81_21# 0.0151f
C9962 hold59/a_391_47# _0853_/a_68_297# 0
C9963 pp[27] acc0.A\[30\] 0.00508f
C9964 _0195_ _0125_ 0.02722f
C9965 _0183_ hold71/a_391_47# 0
C9966 clknet_1_0__leaf__0465_ _0441_ 0
C9967 _0457_ _1015_/a_561_413# 0
C9968 net21 _0172_ 0.42349f
C9969 _0329_ _1008_/a_891_413# 0
C9970 _0753_/a_297_297# hold30/a_49_47# 0
C9971 _0327_ _0686_/a_301_297# 0
C9972 _0349_ net209 0
C9973 net36 _0346_ 0.02111f
C9974 _0350_ _0379_ 0.28313f
C9975 _1001_/a_1017_47# VPWR 0
C9976 _0372_ _0350_ 0.02687f
C9977 _0964_/a_109_297# _0478_ 0
C9978 net45 _1017_/a_975_413# 0
C9979 VPWR _1062_/a_592_47# 0
C9980 _0247_ _0240_ 0.01067f
C9981 _0157_ net229 0.09981f
C9982 _1018_/a_634_159# _0347_ 0
C9983 _0849_/a_510_47# acc0.A\[15\] 0.00118f
C9984 _1039_/a_381_47# _0137_ 0.12469f
C9985 _1021_/a_561_413# VPWR 0.00321f
C9986 _0369_ _0247_ 0
C9987 _1038_/a_1059_315# _0135_ 0
C9988 hold58/a_49_47# _0557_/a_149_47# 0
C9989 _0762_/a_510_47# _0369_ 0.00199f
C9990 _0279_ _0647_/a_285_47# 0.07414f
C9991 _0343_ _0758_/a_510_47# 0
C9992 clkbuf_0__0458_/a_110_47# _0841_/a_215_47# 0
C9993 clkbuf_1_0__f__0457_/a_110_47# _0369_ 0.00352f
C9994 _0453_ clknet_1_0__leaf__0461_ 0
C9995 _1000_/a_27_47# _0773_/a_35_297# 0
C9996 clkbuf_1_0__f__0457_/a_110_47# clknet_0__0457_ 0.42929f
C9997 _0984_/a_891_413# clkbuf_1_0__f__0458_/a_110_47# 0.01653f
C9998 _0346_ _0811_/a_81_21# 0.1744f
C9999 net36 _0935_/a_27_47# 0
C10000 _1011_/a_193_47# _0332_ 0
C10001 _0308_ _0306_ 0.31115f
C10002 net36 _1061_/a_193_47# 0
C10003 _0234_ net49 0.00172f
C10004 acc0.A\[23\] net52 0.00644f
C10005 net105 _0181_ 0.00176f
C10006 net69 _0635_/a_109_297# 0
C10007 net238 clkbuf_1_1__f__0459_/a_110_47# 0
C10008 _0642_/a_27_413# VPWR 0.20448f
C10009 _1065_/a_1059_315# _1065_/a_1017_47# 0
C10010 hold18/a_49_47# _0844_/a_79_21# 0
C10011 _0677_/a_47_47# _0352_ 0
C10012 _0677_/a_285_47# _0347_ 0.00406f
C10013 net232 clknet_1_1__leaf_clk 0.03688f
C10014 _0629_/a_59_75# net36 0
C10015 _0999_/a_891_413# net41 0
C10016 _0967_/a_215_297# _1066_/a_466_413# 0
C10017 hold69/a_391_47# _0460_ 0.004f
C10018 _0508_/a_299_297# _0185_ 0.00863f
C10019 hold28/a_391_47# VPWR 0.16494f
C10020 net228 acc0.A\[13\] 0.09558f
C10021 hold66/a_285_47# _1005_/a_466_413# 0
C10022 _0998_/a_1017_47# _0218_ 0
C10023 _0343_ net216 0
C10024 _0428_ _0190_ 0.00248f
C10025 _0467_ hold89/a_391_47# 0
C10026 _0186_ _0522_/a_27_297# 0.12527f
C10027 net168 acc0.A\[6\] 0.07741f
C10028 _0520_/a_373_47# net13 0
C10029 _1036_/a_466_413# B[15] 0
C10030 _1068_/a_1059_315# _0487_ 0.00181f
C10031 _0723_/a_207_413# _0333_ 0
C10032 _0856_/a_79_21# net247 0.0018f
C10033 _0707_/a_75_199# _0338_ 0.07184f
C10034 _0707_/a_201_297# _0335_ 0.00594f
C10035 comp0.B\[11\] _1042_/a_381_47# 0.01857f
C10036 comp0.B\[12\] _1042_/a_891_413# 0
C10037 _1014_/a_466_413# _1014_/a_561_413# 0.00772f
C10038 _1014_/a_634_159# _1014_/a_975_413# 0
C10039 _1071_/a_27_47# _1071_/a_1059_315# 0.04875f
C10040 _1071_/a_193_47# _1071_/a_466_413# 0.0802f
C10041 net152 net20 0
C10042 acc0.A\[15\] hold71/a_391_47# 0.05085f
C10043 net4 net143 0
C10044 _0996_/a_193_47# _0796_/a_215_47# 0
C10045 B[4] control0.sh 0
C10046 _1015_/a_193_47# _0208_ 0.48307f
C10047 _1015_/a_1059_315# _0173_ 0
C10048 input21/a_75_212# input19/a_75_212# 0
C10049 net56 net242 0.46034f
C10050 _0816_/a_150_297# _0347_ 0.00135f
C10051 clkbuf_1_1__f__0463_/a_110_47# _0496_/a_27_47# 0.0151f
C10052 _0985_/a_891_413# _0458_ 0.01561f
C10053 _0183_ clkbuf_0__0459_/a_110_47# 0.00598f
C10054 _0798_/a_113_297# net5 0
C10055 hold56/a_391_47# _0163_ 0
C10056 VPWR _0105_ 0.45269f
C10057 _0137_ net174 0
C10058 _0179_ net137 0
C10059 _0343_ _0230_ 0.03246f
C10060 _0499_/a_59_75# _0175_ 0
C10061 _0217_ _0386_ 0
C10062 _0617_/a_150_297# _0460_ 0
C10063 _0572_/a_27_297# _1026_/a_193_47# 0
C10064 _0836_/a_68_297# _0989_/a_27_47# 0
C10065 VPWR _0536_/a_149_47# 0
C10066 hold33/a_49_47# net10 0
C10067 _0717_/a_303_47# _0334_ 0
C10068 _1055_/a_1017_47# net16 0
C10069 hold13/a_391_47# _0175_ 0
C10070 net212 _0989_/a_27_47# 0.01242f
C10071 hold25/a_49_47# hold25/a_285_47# 0.22264f
C10072 _0305_ _1059_/a_634_159# 0.0201f
C10073 clkbuf_1_0__f__0459_/a_110_47# _1017_/a_381_47# 0
C10074 comp0.B\[15\] comp0.B\[0\] 0.04937f
C10075 net86 net219 0.03788f
C10076 net45 _0581_/a_109_47# 0.00179f
C10077 clknet_1_1__leaf__0465_ net74 0
C10078 hold63/a_391_47# net111 0.02262f
C10079 _1015_/a_27_47# net17 0
C10080 VPWR _0848_/a_27_47# 0.00602f
C10081 _0285_ _0283_ 0.00965f
C10082 _0340_ pp[31] 0
C10083 net2 _0510_/a_109_47# 0.00191f
C10084 _0514_/a_27_297# _0187_ 0
C10085 net168 _0523_/a_384_47# 0
C10086 _1026_/a_381_47# acc0.A\[25\] 0.03171f
C10087 _0454_ _0852_/a_285_297# 0.07195f
C10088 net36 _1039_/a_193_47# 0.07392f
C10089 net88 _1067_/a_193_47# 0
C10090 _0195_ _1048_/a_27_47# 0
C10091 _0243_ _0772_/a_79_21# 0
C10092 _0770_/a_79_21# net223 0.00127f
C10093 _1042_/a_27_47# _0542_/a_51_297# 0
C10094 hold78/a_391_47# _0344_ 0
C10095 _1012_/a_27_47# _0352_ 0.03877f
C10096 _1012_/a_466_413# _0347_ 0.00764f
C10097 output54/a_27_47# hold9/a_391_47# 0
C10098 hold67/a_391_47# acc0.A\[8\] 0
C10099 _1056_/a_1017_47# _0186_ 0
C10100 _0210_ _0176_ 0.01753f
C10101 VPWR _0218_ 6.56461f
C10102 net149 control0.sh 0
C10103 clknet_1_1__leaf__0462_ _0345_ 0.30852f
C10104 _0343_ _1016_/a_634_159# 0.0053f
C10105 clknet_1_0__leaf__0462_ _0231_ 0
C10106 clknet_1_0__leaf__0462_ _0575_/a_109_47# 0
C10107 _0582_/a_27_297# acc0.A\[18\] 0
C10108 _0831_/a_285_297# acc0.A\[6\] 0.03793f
C10109 clknet_1_0__leaf__0465_ hold83/a_49_47# 0
C10110 _0216_ _1010_/a_634_159# 0
C10111 hold15/a_285_47# _0340_ 0
C10112 hold15/a_391_47# _0341_ 0
C10113 output48/a_27_47# pp[23] 0
C10114 _0981_/a_109_297# net167 0.01111f
C10115 _0981_/a_109_47# _0490_ 0.00149f
C10116 clknet_1_0__leaf__0459_ _1060_/a_891_413# 0
C10117 _0216_ acc0.A\[30\] 0.30665f
C10118 _1052_/a_634_159# _0180_ 0.01185f
C10119 _1042_/a_466_413# net20 0
C10120 hold49/a_49_47# net196 0
C10121 _0222_ _1022_/a_1017_47# 0.00189f
C10122 _0963_/a_35_297# control0.count\[1\] 0.1201f
C10123 _0500_/a_27_47# _0180_ 0.04645f
C10124 net59 pp[30] 0.01395f
C10125 clkbuf_0__0459_/a_110_47# acc0.A\[15\] 0.07495f
C10126 _0500_/a_27_47# net218 0
C10127 _0179_ hold71/a_391_47# 0
C10128 _0571_/a_109_297# _1026_/a_891_413# 0
C10129 hold42/a_285_47# output37/a_27_47# 0
C10130 _0553_/a_149_47# net29 0.00108f
C10131 _0223_ _0315_ 0
C10132 _0424_ _0423_ 0.06687f
C10133 net144 A[12] 0.0053f
C10134 _0278_ clkbuf_1_1__f__0459_/a_110_47# 0
C10135 _0253_ _0829_/a_27_47# 0
C10136 _0459_ _0612_/a_145_75# 0
C10137 _0352_ _0242_ 0.02113f
C10138 _0344_ net163 0
C10139 _1013_/a_381_47# pp[31] 0
C10140 _0498_/a_51_297# _0159_ 0.10284f
C10141 _0498_/a_240_47# net247 0.04108f
C10142 net22 _0546_/a_149_47# 0
C10143 _0498_/a_149_47# net7 0.00351f
C10144 _0220_ _0567_/a_109_47# 0
C10145 _0084_ _0986_/a_27_47# 0.09151f
C10146 _0445_ _0986_/a_634_159# 0
C10147 _0113_ clknet_1_0__leaf__0461_ 0.03048f
C10148 _0399_ _0988_/a_193_47# 0.00517f
C10149 _1038_/a_634_159# _0136_ 0
C10150 comp0.B\[2\] _1033_/a_561_413# 0.00284f
C10151 _0557_/a_512_297# _0134_ 0
C10152 acc0.A\[22\] _1005_/a_1059_315# 0
C10153 net150 _1005_/a_381_47# 0.00735f
C10154 clkload1/a_268_47# _0257_ 0.00105f
C10155 _0126_ _1028_/a_1059_315# 0
C10156 _0189_ _0181_ 0.02429f
C10157 clknet_1_0__leaf__0465_ input13/a_75_212# 0.05281f
C10158 _1032_/a_193_47# _0565_/a_51_297# 0
C10159 _0350_ net244 0.08871f
C10160 hold36/a_285_47# _0174_ 0
C10161 _1022_/a_27_47# _1022_/a_634_159# 0.14145f
C10162 acc0.A\[31\] _1013_/a_634_159# 0
C10163 net162 _1013_/a_27_47# 0
C10164 _0178_ _0584_/a_27_297# 0
C10165 _0576_/a_109_47# acc0.A\[23\] 0.00137f
C10166 _0442_ clknet_0__0465_ 0
C10167 _1003_/a_381_47# clknet_1_0__leaf__0460_ 0.01002f
C10168 _1021_/a_634_159# _0462_ 0
C10169 _1059_/a_381_47# acc0.A\[15\] 0.00233f
C10170 _0717_/a_209_47# pp[27] 0
C10171 VPWR _0775_/a_215_47# 0.01183f
C10172 hold20/a_285_47# VPWR 0.30016f
C10173 net98 _0347_ 0.00909f
C10174 _1018_/a_891_413# _0116_ 0.0334f
C10175 net149 net157 0.30422f
C10176 _0957_/a_32_297# comp0.B\[5\] 0
C10177 _0579_/a_109_47# _1001_/a_27_47# 0
C10178 output65/a_27_47# output63/a_27_47# 0.00151f
C10179 _1008_/a_891_413# _1008_/a_975_413# 0.00851f
C10180 _1008_/a_27_47# net94 0.23041f
C10181 _1008_/a_381_47# _1008_/a_561_413# 0.00123f
C10182 _1055_/a_634_159# _1055_/a_1059_315# 0
C10183 _1055_/a_27_47# _1055_/a_381_47# 0.06222f
C10184 _1055_/a_193_47# _1055_/a_891_413# 0.19685f
C10185 _0466_ _0167_ 0.00133f
C10186 clkbuf_1_0__f__0459_/a_110_47# acc0.A\[14\] 0.00391f
C10187 net203 comp0.B\[0\] 0.00459f
C10188 pp[16] _0995_/a_1059_315# 0
C10189 _0337_ _1011_/a_1059_315# 0
C10190 _1020_/a_381_47# _0118_ 0.13417f
C10191 net53 _1025_/a_561_413# 0
C10192 pp[25] _1025_/a_891_413# 0
C10193 _0305_ clknet_0__0461_ 0.03343f
C10194 net242 _0345_ 0
C10195 clkbuf_0__0461_/a_110_47# _0775_/a_79_21# 0.00905f
C10196 _0343_ _0116_ 0.00117f
C10197 _0559_/a_512_297# _0173_ 0
C10198 _1035_/a_1017_47# comp0.B\[5\] 0
C10199 _1003_/a_193_47# _1003_/a_466_413# 0.07482f
C10200 _1003_/a_27_47# _1003_/a_1059_315# 0.04875f
C10201 _0399_ net72 0.0032f
C10202 clkbuf_1_0__f__0464_/a_110_47# _0147_ 0.00143f
C10203 net23 comp0.B\[5\] 0
C10204 _1055_/a_466_413# net181 0
C10205 _1016_/a_891_413# _0114_ 0
C10206 _0750_/a_181_47# net48 0
C10207 _0230_ _0376_ 0.04455f
C10208 _1001_/a_193_47# _0399_ 0
C10209 _0390_ _0218_ 0.09767f
C10210 _0289_ _0508_/a_299_297# 0
C10211 clknet_0__0458_ _0986_/a_592_47# 0
C10212 _0954_/a_32_297# clknet_1_1__leaf__0464_ 0.0017f
C10213 net114 hold50/a_391_47# 0.03868f
C10214 clknet_0__0457_ _1014_/a_592_47# 0
C10215 hold58/a_49_47# hold58/a_391_47# 0.00188f
C10216 _0343_ _0236_ 0
C10217 net84 _1017_/a_891_413# 0
C10218 _0525_/a_81_21# net148 0
C10219 hold67/a_285_47# _0290_ 0
C10220 _0275_ _0425_ 0.00127f
C10221 VPWR _0690_/a_150_297# 0.00115f
C10222 _0833_/a_215_47# _0439_ 0.00549f
C10223 _0997_/a_466_413# _0219_ 0.00792f
C10224 _0997_/a_561_413# _0345_ 0.00124f
C10225 _0216_ _0779_/a_79_21# 0
C10226 _1004_/a_1059_315# _0758_/a_215_47# 0
C10227 _1004_/a_27_47# _0347_ 0.00609f
C10228 net54 _0324_ 0
C10229 acc0.A\[1\] clknet_1_1__leaf__0457_ 0.30014f
C10230 _0199_ clkbuf_1_1__f__0457_/a_110_47# 0.01228f
C10231 VPWR _0833_/a_215_47# 0
C10232 hold75/a_391_47# net47 0
C10233 net17 _0215_ 0.09916f
C10234 hold87/a_49_47# _0181_ 0.05754f
C10235 _0307_ hold72/a_391_47# 0
C10236 _0126_ _0347_ 0
C10237 net190 _0352_ 0
C10238 clknet_0__0459_ _0094_ 0.08945f
C10239 _1054_/a_27_47# _1053_/a_466_413# 0.00105f
C10240 _0559_/a_149_47# _0212_ 0.00154f
C10241 _0982_/a_1059_315# _0456_ 0.00401f
C10242 _0982_/a_561_413# net234 0
C10243 _0144_ net135 0.00766f
C10244 comp0.B\[4\] net24 0.05589f
C10245 net200 net199 0.00122f
C10246 _0191_ _0433_ 0
C10247 _1058_/a_27_47# net189 0.03719f
C10248 net187 _0183_ 0.13186f
C10249 net247 _0846_/a_51_297# 0
C10250 _0280_ _0287_ 0.0161f
C10251 VPWR _0177_ 0.50599f
C10252 _0951_/a_209_311# _0468_ 0
C10253 _0179_ _1059_/a_381_47# 0
C10254 _0409_ hold91/a_285_47# 0
C10255 _0180_ A[8] 0
C10256 net86 _0352_ 0.00296f
C10257 _0985_/a_1059_315# _0268_ 0
C10258 pp[30] _0335_ 0
C10259 _0398_ net221 0
C10260 net59 _0339_ 0.00248f
C10261 _0462_ _0586_/a_27_47# 0
C10262 net46 _0606_/a_215_297# 0.0057f
C10263 _0387_ _0780_/a_117_297# 0
C10264 net208 _0220_ 0.00537f
C10265 _0982_/a_27_47# _0452_ 0
C10266 VPWR _0112_ 0.34626f
C10267 _0257_ _0836_/a_68_297# 0
C10268 clknet_1_0__leaf_clk _1064_/a_634_159# 0
C10269 _1048_/a_27_47# _1048_/a_193_47# 0.96639f
C10270 net214 net142 0
C10271 VPWR _1017_/a_975_413# 0.00418f
C10272 _0717_/a_209_297# pp[28] 0.003f
C10273 _0106_ hold50/a_49_47# 0
C10274 _0365_ hold50/a_391_47# 0.05397f
C10275 clknet_0__0458_ _0449_ 0
C10276 clknet_1_0__leaf__0459_ _0218_ 0.35591f
C10277 _0833_/a_215_47# output62/a_27_47# 0
C10278 VPWR input25/a_75_212# 0.21833f
C10279 _0223_ _0742_/a_81_21# 0
C10280 net70 net229 0
C10281 _0563_/a_149_47# _0563_/a_240_47# 0.06872f
C10282 _0563_/a_51_297# _0214_ 0.116f
C10283 _0548_/a_149_47# net173 0.01268f
C10284 _0829_/a_27_47# output61/a_27_47# 0
C10285 _0179_ clkload2/a_110_47# 0
C10286 _0113_ _0585_/a_27_297# 0
C10287 _0096_ _0459_ 0
C10288 _1017_/a_381_47# clkbuf_0__0461_/a_110_47# 0
C10289 VPWR _1033_/a_891_413# 0.19128f
C10290 net61 _0438_ 0
C10291 clknet_1_0__leaf__0465_ _1049_/a_891_413# 0
C10292 _0343_ hold62/a_391_47# 0.00167f
C10293 _0783_/a_79_21# _0218_ 0
C10294 hold86/a_391_47# VPWR 0.1719f
C10295 net190 net115 0
C10296 VPWR _1050_/a_592_47# 0
C10297 _0217_ _0854_/a_79_21# 0
C10298 net36 _1041_/a_1059_315# 0
C10299 _0179_ _0519_/a_299_297# 0.05851f
C10300 _0151_ _1054_/a_27_47# 0.00295f
C10301 net61 _0636_/a_59_75# 0.20818f
C10302 hold33/a_391_47# net31 0
C10303 net45 _0792_/a_80_21# 0
C10304 _0275_ _0432_ 0.02219f
C10305 _1010_/a_1059_315# _1010_/a_891_413# 0.31086f
C10306 _1010_/a_193_47# _1010_/a_975_413# 0
C10307 _1010_/a_466_413# _1010_/a_381_47# 0.03733f
C10308 net178 acc0.A\[9\] 0
C10309 clknet_1_0__leaf__0462_ _1004_/a_381_47# 0.00253f
C10310 _1056_/a_193_47# _0514_/a_27_297# 0
C10311 _1056_/a_27_47# _0514_/a_109_297# 0
C10312 output40/a_27_47# net6 0
C10313 net60 net41 0.01419f
C10314 hold55/a_285_47# _1015_/a_27_47# 0.00123f
C10315 hold92/a_49_47# _0345_ 0.0064f
C10316 _0991_/a_381_47# _0181_ 0
C10317 _1040_/a_193_47# _1040_/a_891_413# 0.19226f
C10318 _1040_/a_27_47# _1040_/a_381_47# 0.05761f
C10319 _1040_/a_634_159# _1040_/a_1059_315# 0
C10320 hold36/a_49_47# net194 0.00229f
C10321 _0452_ _0446_ 0
C10322 hold79/a_285_47# _0976_/a_76_199# 0.0022f
C10323 _0475_ _0494_/a_27_47# 0
C10324 _0979_/a_27_297# _0979_/a_109_297# 0.17136f
C10325 net5 net41 0.13208f
C10326 _0229_ _0225_ 0
C10327 _0146_ _1048_/a_381_47# 0.13112f
C10328 net22 _0176_ 0.02763f
C10329 _0697_/a_472_297# _0328_ 0.00145f
C10330 _0432_ _0837_/a_585_47# 0
C10331 _0519_/a_81_21# net75 0
C10332 _0527_/a_27_297# _0527_/a_109_297# 0.17136f
C10333 _0195_ _1027_/a_634_159# 0
C10334 _0216_ _1027_/a_27_47# 0.08529f
C10335 VPWR net240 0.31745f
C10336 _0453_ _0218_ 0
C10337 _1002_/a_561_413# _0217_ 0
C10338 _1002_/a_891_413# _0183_ 0.01f
C10339 _0328_ _0695_/a_300_47# 0.00264f
C10340 _0550_/a_51_297# net153 0
C10341 _0222_ net110 0
C10342 VPWR _0099_ 0.27352f
C10343 _0375_ _0238_ 0
C10344 _1020_/a_1017_47# _0461_ 0
C10345 _0846_/a_245_297# _0846_/a_240_47# 0
C10346 acc0.A\[14\] _0996_/a_193_47# 0.01622f
C10347 net45 _1016_/a_1059_315# 0.00316f
C10348 _1067_/a_634_159# _1067_/a_1059_315# 0
C10349 _1067_/a_27_47# _1067_/a_381_47# 0.06222f
C10350 _1067_/a_193_47# _1067_/a_891_413# 0.19497f
C10351 net9 _0987_/a_466_413# 0.00844f
C10352 net104 _0347_ 0.00186f
C10353 _0968_/a_193_297# _0468_ 0
C10354 net156 acc0.A\[25\] 0
C10355 clknet_1_0__leaf__0459_ _0775_/a_215_47# 0
C10356 hold31/a_391_47# _0369_ 0.00462f
C10357 _1019_/a_193_47# _1015_/a_193_47# 0.00149f
C10358 _0805_/a_27_47# _0805_/a_109_47# 0.00517f
C10359 _0314_ _0682_/a_68_297# 0.1071f
C10360 clknet_1_0__leaf__0463_ _0176_ 0.2181f
C10361 _1071_/a_193_47# _0480_ 0
C10362 _1072_/a_634_159# _1071_/a_1059_315# 0
C10363 _0985_/a_27_47# _0529_/a_27_297# 0.01072f
C10364 _1000_/a_634_159# _0392_ 0
C10365 _0181_ clknet_0__0461_ 0.05221f
C10366 VPWR _0359_ 1.68384f
C10367 clknet_1_0__leaf__0462_ _0225_ 0.01411f
C10368 VPWR _0581_/a_109_47# 0
C10369 net70 clknet_0__0458_ 0
C10370 _0313_ _0368_ 0.04762f
C10371 _1009_/a_634_159# _1009_/a_592_47# 0
C10372 acc0.A\[22\] _0592_/a_68_297# 0.16714f
C10373 net65 _0989_/a_634_159# 0.03621f
C10374 acc0.A\[7\] _0989_/a_193_47# 0
C10375 _0195_ _0700_/a_113_47# 0
C10376 VPWR net15 0.20841f
C10377 _0989_/a_634_159# _0989_/a_466_413# 0.23992f
C10378 _0989_/a_193_47# _0989_/a_1059_315# 0.03405f
C10379 _0989_/a_27_47# _0989_/a_891_413# 0.03224f
C10380 net32 _0203_ 0
C10381 comp0.B\[13\] hold36/a_285_47# 0
C10382 control0.state\[1\] _0950_/a_75_212# 0
C10383 _0956_/a_220_297# net201 0
C10384 net7 _0540_/a_51_297# 0
C10385 _0316_ net54 0
C10386 _0717_/a_80_21# _0335_ 0.14542f
C10387 _0982_/a_975_413# VPWR 0.00468f
C10388 _0348_ _0707_/a_75_199# 0.11125f
C10389 _0476_ _1066_/a_561_413# 0
C10390 hold66/a_285_47# _0103_ 0
C10391 _0992_/a_634_159# _0992_/a_466_413# 0.23992f
C10392 _0992_/a_193_47# _0992_/a_1059_315# 0.03405f
C10393 _0992_/a_27_47# _0992_/a_891_413# 0.03224f
C10394 _1036_/a_1017_47# net121 0
C10395 _0695_/a_80_21# clkbuf_1_0__f__0462_/a_110_47# 0
C10396 net24 _0563_/a_245_297# 0
C10397 _0186_ _0193_ 0.51634f
C10398 net161 B[15] 0
C10399 _0606_/a_109_53# VPWR 0.10892f
C10400 _0428_ _0346_ 0.02619f
C10401 VPWR _1053_/a_1059_315# 0.40125f
C10402 _0607_/a_109_47# net43 0.00145f
C10403 _0718_/a_129_47# pp[27] 0
C10404 _0335_ _0339_ 0
C10405 _0125_ _1027_/a_466_413# 0.00493f
C10406 acc0.A\[27\] _1027_/a_381_47# 0
C10407 _1032_/a_381_47# net118 0
C10408 _0280_ _0655_/a_297_297# 0.00216f
C10409 net226 _0168_ 0.18605f
C10410 _0355_ _1029_/a_27_47# 0
C10411 _0354_ _1029_/a_193_47# 0
C10412 _1014_/a_1059_315# acc0.A\[0\] 0.13055f
C10413 _0272_ clkbuf_0__0458_/a_110_47# 0
C10414 _1014_/a_975_413# net100 0
C10415 _1071_/a_891_413# _1071_/a_1017_47# 0.00617f
C10416 hold55/a_391_47# _0566_/a_27_47# 0
C10417 net54 _0347_ 0.04507f
C10418 net48 net240 0.00157f
C10419 _0996_/a_561_413# net238 0.00178f
C10420 _1045_/a_1059_315# _1043_/a_27_47# 0
C10421 _0433_ clkbuf_1_0__f__0465_/a_110_47# 0.1109f
C10422 hold75/a_49_47# _0267_ 0.00265f
C10423 _1000_/a_466_413# clknet_0__0461_ 0.00518f
C10424 _0256_ acc0.A\[3\] 0
C10425 _0713_/a_27_47# _0208_ 0.22425f
C10426 _0263_ _0345_ 0.45624f
C10427 _0346_ hold60/a_391_47# 0.02259f
C10428 _0935_/a_27_47# _1061_/a_27_47# 0
C10429 _1061_/a_27_47# _1061_/a_193_47# 0.97453f
C10430 _0983_/a_27_47# net206 0
C10431 hold54/a_391_47# _0565_/a_51_297# 0
C10432 net187 hold40/a_285_47# 0.02157f
C10433 net200 VPWR 0.31561f
C10434 _0659_/a_68_297# _0990_/a_193_47# 0
C10435 hold39/a_391_47# net186 0.13298f
C10436 _0216_ _1026_/a_466_413# 0.0064f
C10437 net155 _1026_/a_1059_315# 0.00187f
C10438 _0195_ _1026_/a_891_413# 0.01895f
C10439 _0124_ _1026_/a_193_47# 0.201f
C10440 net157 _1046_/a_891_413# 0
C10441 _0736_/a_56_297# _0362_ 0.04484f
C10442 _0216_ _1024_/a_561_413# 0
C10443 _0817_/a_81_21# _0288_ 0.00133f
C10444 _0817_/a_368_297# acc0.A\[9\] 0.00165f
C10445 _0549_/a_68_297# _0207_ 0.10673f
C10446 _0437_ _0989_/a_1017_47# 0
C10447 _0549_/a_150_297# net171 0
C10448 _0305_ net145 0
C10449 acc0.A\[24\] _1006_/a_891_413# 0
C10450 _0179_ _0148_ 0.10516f
C10451 _0190_ _0988_/a_193_47# 0
C10452 _0172_ _0173_ 0
C10453 _0343_ acc0.A\[8\] 0.30206f
C10454 clkload1/a_268_47# clknet_1_1__leaf__0458_ 0
C10455 _1020_/a_891_413# acc0.A\[20\] 0.00591f
C10456 _0181_ _0082_ 0.00253f
C10457 clkbuf_1_0__f__0459_/a_110_47# _1016_/a_634_159# 0.00141f
C10458 _0243_ _1019_/a_27_47# 0
C10459 _0189_ _0187_ 0.00313f
C10460 acc0.A\[26\] acc0.A\[25\] 0.02701f
C10461 _0304_ _0420_ 0
C10462 _0217_ _1014_/a_193_47# 0.45465f
C10463 _0390_ _0099_ 0
C10464 clkbuf_1_1__f__0462_/a_110_47# _0350_ 0.01916f
C10465 _0555_/a_240_47# _0175_ 0
C10466 clknet_1_0__leaf__0459_ _0112_ 0
C10467 pp[7] A[8] 0
C10468 _1033_/a_975_413# _0215_ 0.00109f
C10469 _0715_/a_27_47# _0346_ 0.36464f
C10470 _0786_/a_300_47# _0345_ 0
C10471 _0984_/a_891_413# acc0.A\[15\] 0.00562f
C10472 _0115_ acc0.A\[18\] 0
C10473 _0343_ _0991_/a_193_47# 0.02732f
C10474 _0789_/a_75_199# _0218_ 0
C10475 _0569_/a_27_297# _1029_/a_27_47# 0
C10476 VPWR _1028_/a_466_413# 0.23896f
C10477 _1069_/a_193_47# _1069_/a_381_47# 0.10164f
C10478 _1069_/a_634_159# _1069_/a_891_413# 0.03684f
C10479 _1069_/a_27_47# _1069_/a_561_413# 0.0027f
C10480 hold4/a_285_47# net109 0.02967f
C10481 hold4/a_49_47# net177 0.0294f
C10482 net1 comp0.B\[15\] 0
C10483 A[11] acc0.A\[11\] 0.00213f
C10484 _0343_ _0773_/a_285_47# 0
C10485 _0535_/a_68_297# _0545_/a_68_297# 0
C10486 _0402_ _0672_/a_510_47# 0
C10487 net10 _0203_ 0.043f
C10488 output43/a_27_47# hold78/a_391_47# 0
C10489 net224 _0362_ 0.00628f
C10490 _1037_/a_466_413# comp0.B\[4\] 0
C10491 _1041_/a_27_47# _1040_/a_193_47# 0.00305f
C10492 _1041_/a_193_47# _1040_/a_27_47# 0.00367f
C10493 _1031_/a_193_47# _0220_ 0.11744f
C10494 _1031_/a_27_47# _0336_ 0
C10495 _0536_/a_512_297# _0172_ 0.00116f
C10496 input31/a_75_212# B[14] 0.00433f
C10497 B[8] input22/a_75_212# 0.00207f
C10498 net69 _0450_ 0
C10499 _0997_/a_1059_315# _0799_/a_80_21# 0
C10500 _0398_ _1017_/a_27_47# 0
C10501 _0571_/a_27_297# acc0.A\[26\] 0
C10502 _1059_/a_634_159# hold82/a_391_47# 0.00982f
C10503 _1059_/a_466_413# hold82/a_285_47# 0.01371f
C10504 _1059_/a_1059_315# hold82/a_49_47# 0.00923f
C10505 _0964_/a_109_297# VPWR 0.00794f
C10506 net81 net6 0
C10507 _0685_/a_68_297# _0321_ 0
C10508 input24/a_75_212# B[1] 0.19876f
C10509 _1030_/a_193_47# net209 0.24522f
C10510 _0596_/a_59_75# net150 0.00511f
C10511 clknet_1_0__leaf__0461_ _0345_ 0.04033f
C10512 VPWR net228 0.80199f
C10513 _0556_/a_68_297# _0554_/a_68_297# 0.01285f
C10514 _1051_/a_27_47# net9 0
C10515 _0305_ net67 0
C10516 _1018_/a_466_413# clkbuf_1_0__f__0461_/a_110_47# 0
C10517 _1018_/a_27_47# clknet_0__0461_ 0.00107f
C10518 _0733_/a_222_93# acc0.A\[25\] 0
C10519 _0718_/a_377_297# pp[28] 0.00331f
C10520 _1002_/a_193_47# _0181_ 0.0139f
C10521 _0592_/a_68_297# _0379_ 0
C10522 _0183_ _0103_ 0
C10523 control0.count\[3\] _0487_ 0.00772f
C10524 _0483_ _0484_ 0.16531f
C10525 _0343_ _0380_ 0
C10526 _0538_/a_245_297# _0538_/a_240_47# 0
C10527 _0833_/a_79_21# acc0.A\[6\] 0
C10528 clknet_1_1__leaf__0462_ _1008_/a_592_47# 0
C10529 comp0.B\[5\] _0213_ 0.05354f
C10530 _0474_ _0561_/a_240_47# 0.0028f
C10531 _0216_ _0315_ 0
C10532 hold43/a_285_47# clknet_1_1__leaf__0462_ 0.00204f
C10533 _0183_ hold18/a_285_47# 0.00622f
C10534 _1022_/a_381_47# _1022_/a_561_413# 0.00123f
C10535 _1022_/a_891_413# _1022_/a_975_413# 0.00851f
C10536 hold75/a_285_47# _0218_ 0.02043f
C10537 _0645_/a_47_47# _0276_ 0
C10538 _1065_/a_27_47# _1062_/a_634_159# 0
C10539 _0174_ _0545_/a_68_297# 0.04886f
C10540 hold2/a_49_47# clknet_1_0__leaf__0461_ 0
C10541 net55 VPWR 1.13523f
C10542 clknet_1_0__leaf__0459_ _0099_ 0
C10543 _0994_/a_634_159# _0994_/a_1059_315# 0
C10544 _0994_/a_27_47# _0994_/a_381_47# 0.06222f
C10545 _0994_/a_193_47# _0994_/a_891_413# 0.19497f
C10546 _1020_/a_634_159# clknet_1_0__leaf__0457_ 0.00168f
C10547 _0285_ _0808_/a_266_47# 0.00567f
C10548 _0284_ _0808_/a_368_297# 0
C10549 _0275_ _0986_/a_381_47# 0.01143f
C10550 _0779_/a_215_47# _0779_/a_510_47# 0.00529f
C10551 _0472_ _0474_ 0.20345f
C10552 net211 _1001_/a_561_413# 0
C10553 net44 _0352_ 0.21281f
C10554 _0328_ _1008_/a_27_47# 0
C10555 B[9] net152 0
C10556 _0179_ _0525_/a_384_47# 0
C10557 _1055_/a_466_413# net179 0.03309f
C10558 _1055_/a_1059_315# net141 0
C10559 VPWR hold3/a_285_47# 0.31597f
C10560 _1023_/a_634_159# output51/a_27_47# 0.00866f
C10561 _0422_ hold81/a_285_47# 0
C10562 hold5/a_285_47# _1043_/a_891_413# 0
C10563 hold5/a_391_47# _1043_/a_1059_315# 0
C10564 hold22/a_49_47# _1053_/a_27_47# 0
C10565 net64 _0343_ 0.42314f
C10566 _0984_/a_891_413# _0179_ 0
C10567 _1003_/a_634_159# net89 0
C10568 net23 hold84/a_49_47# 0
C10569 _1003_/a_193_47# _0101_ 0.57059f
C10570 _1003_/a_891_413# _1003_/a_1017_47# 0.00617f
C10571 _0343_ _0621_/a_117_297# 0.00482f
C10572 net36 _1047_/a_466_413# 0.01594f
C10573 _0984_/a_193_47# _0181_ 0
C10574 hold26/a_49_47# _0174_ 0.01811f
C10575 _1036_/a_1059_315# net27 0
C10576 _0207_ _1040_/a_891_413# 0
C10577 _0751_/a_29_53# _0374_ 0.08637f
C10578 hold2/a_285_47# net47 0
C10579 comp0.B\[1\] _0584_/a_27_297# 0.02149f
C10580 _1039_/a_27_47# _1039_/a_193_47# 0.95936f
C10581 _0258_ _0346_ 0.23506f
C10582 _0967_/a_403_297# VPWR 0.00569f
C10583 control0.count\[1\] _0484_ 0
C10584 _0836_/a_68_297# clknet_1_1__leaf__0458_ 0.00612f
C10585 _1020_/a_27_47# _0457_ 0.01236f
C10586 _0197_ _0529_/a_27_297# 0.1095f
C10587 _0343_ _0423_ 0
C10588 _0212_ comp0.B\[5\] 0.43519f
C10589 net185 comp0.B\[6\] 0.0451f
C10590 clknet_0__0458_ _0260_ 0.01362f
C10591 hold46/a_391_47# _0172_ 0.00116f
C10592 _0663_/a_27_413# _0661_/a_27_297# 0.01902f
C10593 _1054_/a_975_413# _0191_ 0.00114f
C10594 _0211_ net28 0.03219f
C10595 net212 clknet_1_1__leaf__0458_ 0.00444f
C10596 _0183_ _0856_/a_215_47# 0.0098f
C10597 _0258_ net65 0.00695f
C10598 _0257_ _0989_/a_891_413# 0
C10599 _0844_/a_79_21# _0448_ 0.10612f
C10600 _1004_/a_975_413# _0352_ 0
C10601 _0518_/a_27_297# _0399_ 0
C10602 _0111_ net60 0
C10603 _0126_ _0106_ 0.00132f
C10604 net33 _1062_/a_193_47# 0
C10605 _0534_/a_299_297# net175 0
C10606 _0983_/a_891_413# _0347_ 0
C10607 hold15/a_391_47# acc0.A\[30\] 0.00336f
C10608 net23 _1065_/a_381_47# 0.01603f
C10609 _0399_ _0208_ 0.02615f
C10610 hold18/a_285_47# acc0.A\[15\] 0.00954f
C10611 clknet_1_1__leaf__0459_ _0400_ 0
C10612 net140 _1053_/a_193_47# 0.03673f
C10613 net169 _1053_/a_27_47# 0
C10614 _0222_ _0618_/a_79_21# 0.12295f
C10615 _0992_/a_193_47# _0809_/a_81_21# 0
C10616 _0285_ _0345_ 0.0219f
C10617 _0392_ _0242_ 0
C10618 VPWR _0792_/a_80_21# 0.15748f
C10619 VPWR _0987_/a_592_47# 0
C10620 _1024_/a_634_159# _1024_/a_381_47# 0
C10621 hold30/a_391_47# _0225_ 0
C10622 net86 hold72/a_285_47# 0
C10623 _0220_ _0395_ 0.0016f
C10624 hold65/a_49_47# _0432_ 0
C10625 _0811_/a_384_47# _0420_ 0
C10626 _0217_ _0369_ 0.02662f
C10627 net16 _0186_ 0.02994f
C10628 net48 hold3/a_285_47# 0.01168f
C10629 _0718_/a_47_47# _0335_ 0
C10630 clknet_0__0457_ _0217_ 0.90309f
C10631 hold56/a_285_47# clkbuf_1_1__f_clk/a_110_47# 0
C10632 hold30/a_49_47# hold29/a_49_47# 0.00442f
C10633 _0797_/a_207_413# net6 0
C10634 _1011_/a_1059_315# _0333_ 0
C10635 _0985_/a_466_413# _0180_ 0.00439f
C10636 _1036_/a_27_47# input25/a_75_212# 0
C10637 net66 acc0.A\[11\] 0.00481f
C10638 _0738_/a_68_297# _0321_ 0
C10639 _0807_/a_68_297# _0281_ 0
C10640 net145 _0181_ 0
C10641 VPWR _1029_/a_592_47# 0
C10642 net61 _0829_/a_27_47# 0.00359f
C10643 _0514_/a_27_297# clknet_1_1__leaf__0465_ 0.05342f
C10644 _0180_ _1049_/a_27_47# 0
C10645 _0644_/a_47_47# acc0.A\[13\] 0.04438f
C10646 comp0.B\[2\] _1032_/a_466_413# 0
C10647 _0231_ _0591_/a_109_297# 0.00314f
C10648 _0540_/a_51_297# _0202_ 0.1238f
C10649 _0540_/a_149_47# _0540_/a_240_47# 0.06872f
C10650 net36 _0782_/a_27_47# 0
C10651 clk _1064_/a_466_413# 0.00461f
C10652 hold96/a_285_47# _0217_ 0.07127f
C10653 _1048_/a_466_413# _1048_/a_592_47# 0.00553f
C10654 _1048_/a_634_159# _1048_/a_1017_47# 0
C10655 net53 _0737_/a_285_297# 0
C10656 _0712_/a_297_297# _0220_ 0.04707f
C10657 _1034_/a_381_47# clknet_1_1__leaf__0463_ 0.00552f
C10658 output64/a_27_47# VPWR 0.38638f
C10659 _0195_ net42 0.00332f
C10660 acc0.A\[14\] _0794_/a_326_47# 0
C10661 hold34/a_285_47# acc0.A\[9\] 0.00575f
C10662 VPWR _0956_/a_32_297# 0.27393f
C10663 VPWR _1016_/a_1059_315# 0.37591f
C10664 _0458_ _0630_/a_109_297# 0
C10665 _0924_/a_27_47# _0178_ 0
C10666 acc0.A\[16\] _0780_/a_117_297# 0
C10667 _0232_ _0368_ 0
C10668 _1035_/a_193_47# net24 0
C10669 _0846_/a_240_47# _0448_ 0.01485f
C10670 _0856_/a_215_47# acc0.A\[15\] 0
C10671 _0312_ _1007_/a_592_47# 0
C10672 _0640_/a_465_297# _0434_ 0
C10673 _0460_ _0219_ 0.14488f
C10674 hold11/a_391_47# net158 0.1316f
C10675 _1016_/a_634_159# clkbuf_0__0461_/a_110_47# 0
C10676 _1060_/a_193_47# _0219_ 0
C10677 _0232_ _0618_/a_215_47# 0.00761f
C10678 hold23/a_285_47# acc0.A\[3\] 0.02168f
C10679 hold27/a_285_47# VPWR 0.27477f
C10680 hold33/a_391_47# net7 0.04394f
C10681 _0216_ control0.add 0
C10682 _0569_/a_27_297# _1028_/a_891_413# 0
C10683 _0569_/a_109_297# _1028_/a_1059_315# 0
C10684 _0216_ _0742_/a_81_21# 0.00296f
C10685 net230 net140 0.00336f
C10686 clknet_0__0465_ _0832_/a_113_47# 0
C10687 clknet_1_1__leaf__0460_ _0731_/a_81_21# 0
C10688 _0179_ hold18/a_285_47# 0
C10689 clknet_0__0461_ clknet_1_1__leaf__0461_ 0.00993f
C10690 _1056_/a_193_47# _0189_ 0.00433f
C10691 hold6/a_49_47# net32 0.02267f
C10692 hold6/a_285_47# net152 0
C10693 _0130_ _1015_/a_561_413# 0
C10694 net67 _0181_ 0.00673f
C10695 _1040_/a_466_413# net174 0.03099f
C10696 _1053_/a_634_159# acc0.A\[6\] 0.00223f
C10697 clknet_1_0__leaf__0465_ _1054_/a_466_413# 0
C10698 _0410_ _0300_ 0
C10699 output64/a_27_47# output62/a_27_47# 0.00151f
C10700 hold79/a_285_47# _0488_ 0.00889f
C10701 hold79/a_49_47# _0466_ 0
C10702 _0357_ _0728_/a_145_75# 0
C10703 _0979_/a_109_297# _0169_ 0.00169f
C10704 _0249_ _1006_/a_27_47# 0.00363f
C10705 _1072_/a_634_159# _1072_/a_381_47# 0
C10706 _0527_/a_373_47# net11 0.00173f
C10707 _0830_/a_510_47# _0186_ 0
C10708 _0751_/a_29_53# _0249_ 0.01478f
C10709 _0183_ _0505_/a_109_47# 0.00217f
C10710 net9 A[4] 0.00184f
C10711 clknet_1_0__leaf__0458_ net165 0.06398f
C10712 _0172_ net153 0.2408f
C10713 _0821_/a_113_47# _0429_ 0.00973f
C10714 acc0.A\[20\] _0346_ 0.01784f
C10715 _0198_ clknet_1_1__leaf__0457_ 0.04418f
C10716 _0372_ net92 0.02788f
C10717 VPWR _0325_ 0.31178f
C10718 net1 _0382_ 0
C10719 net237 hold90/a_285_47# 0.01019f
C10720 _0477_ clknet_0_clk 0
C10721 _1037_/a_1059_315# _0549_/a_68_297# 0
C10722 _0221_ hold80/a_285_47# 0
C10723 _1067_/a_27_47# control0.add 0.00385f
C10724 net9 _0085_ 0.03268f
C10725 _0283_ net228 0.04047f
C10726 net217 _0281_ 0
C10727 comp0.B\[4\] _0561_/a_149_47# 0.00119f
C10728 _0429_ _0989_/a_891_413# 0.01089f
C10729 _0251_ _0989_/a_561_413# 0
C10730 hold31/a_49_47# net178 0
C10731 net105 _1015_/a_27_47# 0
C10732 _0342_ _0999_/a_1059_315# 0
C10733 _0713_/a_27_47# _1019_/a_193_47# 0
C10734 _1003_/a_193_47# net35 0
C10735 net86 _0392_ 0
C10736 clknet_1_1__leaf__0460_ _1006_/a_193_47# 0
C10737 _0985_/a_634_159# net10 0.01108f
C10738 _0476_ _0175_ 0.03291f
C10739 _0343_ _0386_ 0.0272f
C10740 _0217_ _1024_/a_27_47# 0.00223f
C10741 _1004_/a_466_413# _0380_ 0
C10742 _1004_/a_1059_315# _0350_ 0.06106f
C10743 _0313_ clknet_0__0460_ 0
C10744 _0997_/a_634_159# _0997_/a_381_47# 0
C10745 _0640_/a_215_297# _0465_ 0.0142f
C10746 hold56/a_285_47# VPWR 0.30213f
C10747 net78 _0289_ 0
C10748 _0181_ _0986_/a_975_413# 0
C10749 net198 _1042_/a_27_47# 0.02572f
C10750 hold36/a_49_47# net132 0.00464f
C10751 _0248_ _0240_ 0
C10752 _0348_ _0338_ 0.15739f
C10753 acc0.A\[16\] net165 0
C10754 VPWR _1051_/a_381_47# 0.07636f
C10755 _0248_ _0369_ 0.2322f
C10756 _0349_ _1010_/a_27_47# 0.00396f
C10757 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0462_/a_110_47# 0
C10758 net39 _0993_/a_27_47# 0
C10759 _0279_ _0399_ 0.21258f
C10760 _0337_ acc0.A\[30\] 0.05523f
C10761 _0238_ VPWR 0.73418f
C10762 _0434_ _0988_/a_27_47# 0
C10763 hold6/a_49_47# _1042_/a_1059_315# 0
C10764 hold6/a_285_47# _1042_/a_466_413# 0
C10765 hold6/a_391_47# _1042_/a_634_159# 0
C10766 VPWR _1045_/a_975_413# 0.00468f
C10767 _0125_ net156 0.00396f
C10768 net54 _0106_ 0.22169f
C10769 clkbuf_1_0__f__0458_/a_110_47# _0445_ 0
C10770 _0218_ _0808_/a_266_47# 0
C10771 hold63/a_391_47# VPWR 0.18917f
C10772 _0793_/a_512_297# _0400_ 0
C10773 _0407_ _0792_/a_209_297# 0
C10774 _0793_/a_149_47# _0405_ 0
C10775 net243 _0756_/a_129_47# 0
C10776 _0098_ clknet_0__0461_ 0
C10777 net45 clkbuf_1_0__f__0461_/a_110_47# 0.0188f
C10778 _1027_/a_634_159# _1027_/a_466_413# 0.23992f
C10779 _1027_/a_193_47# _1027_/a_1059_315# 0.03405f
C10780 _1027_/a_27_47# _1027_/a_891_413# 0.03224f
C10781 _1055_/a_193_47# net47 0.00138f
C10782 _0626_/a_68_297# _0261_ 0
C10783 comp0.B\[13\] hold26/a_49_47# 0.01227f
C10784 acc0.A\[15\] _0505_/a_109_47# 0
C10785 _0996_/a_634_159# net41 0
C10786 VPWR _1032_/a_193_47# 0.30413f
C10787 _1061_/a_466_413# _1061_/a_592_47# 0.00553f
C10788 _1061_/a_634_159# _1061_/a_1017_47# 0
C10789 _0753_/a_297_297# _0222_ 0.04558f
C10790 _0305_ _1009_/a_193_47# 0.00298f
C10791 acc0.A\[8\] _0990_/a_381_47# 0
C10792 _0210_ net28 0.01176f
C10793 hold6/a_49_47# net10 0.04804f
C10794 _0224_ _0380_ 0
C10795 clkbuf_0__0460_/a_110_47# _0368_ 0
C10796 acc0.A\[2\] _0465_ 0.00379f
C10797 clkbuf_1_0__f__0457_/a_110_47# hold40/a_391_47# 0.00259f
C10798 hold101/a_49_47# _0441_ 0
C10799 _1007_/a_1017_47# _0219_ 0
C10800 _0105_ _0345_ 0.00832f
C10801 _0984_/a_1059_315# net165 0
C10802 _0746_/a_81_21# _0460_ 0
C10803 hold29/a_391_47# _0757_/a_68_297# 0
C10804 _1032_/a_27_47# _1015_/a_1059_315# 0
C10805 _1035_/a_193_47# _1035_/a_381_47# 0.09503f
C10806 _1035_/a_634_159# _1035_/a_891_413# 0.03684f
C10807 _1035_/a_27_47# _1035_/a_561_413# 0.0027f
C10808 _0298_ net238 0
C10809 _0404_ _0410_ 0.00112f
C10810 _0730_/a_79_21# _0729_/a_68_297# 0
C10811 _0278_ _0277_ 0.10965f
C10812 _0770_/a_79_21# _0350_ 0.01973f
C10813 net185 net26 0.0053f
C10814 _1053_/a_193_47# input14/a_75_212# 0
C10815 clknet_1_0__leaf__0462_ hold68/a_391_47# 0.01409f
C10816 _1000_/a_27_47# _0247_ 0.03563f
C10817 _0092_ _0414_ 0.11561f
C10818 _0489_ _1069_/a_561_413# 0.00121f
C10819 acc0.A\[31\] _0338_ 0
C10820 clknet_1_0__leaf__0462_ _0462_ 0
C10821 _0983_/a_27_47# _0849_/a_215_47# 0
C10822 _0287_ _0815_/a_113_297# 0
C10823 _0661_/a_277_297# _0425_ 0
C10824 _1013_/a_466_413# clknet_1_1__leaf__0461_ 0
C10825 _1048_/a_27_47# acc0.A\[15\] 0
C10826 _0848_/a_27_47# _0345_ 0.00127f
C10827 VPWR _0268_ 0.57136f
C10828 VPWR _0767_/a_145_75# 0
C10829 _1010_/a_193_47# _0701_/a_80_21# 0
C10830 _1010_/a_27_47# _0701_/a_209_297# 0
C10831 _0764_/a_81_21# _0764_/a_299_297# 0.08213f
C10832 net169 A[5] 0
C10833 _0216_ clknet_1_1__leaf__0457_ 0.0019f
C10834 VPWR _0721_/a_27_47# 0.37312f
C10835 comp0.B\[15\] control0.sh 0.04206f
C10836 _1054_/a_193_47# acc0.A\[8\] 0
C10837 acc0.A\[15\] _0506_/a_384_47# 0
C10838 _0127_ _1029_/a_27_47# 0
C10839 acc0.A\[29\] _1029_/a_466_413# 0.00196f
C10840 _0218_ _0345_ 0.3521f
C10841 output55/a_27_47# _0333_ 0.02781f
C10842 _0814_/a_27_47# _0218_ 0
C10843 clknet_1_0__leaf__0459_ _1016_/a_1059_315# 0.01139f
C10844 _1069_/a_1059_315# _0167_ 0
C10845 _1069_/a_891_413# clknet_1_0__leaf_clk 0
C10846 _1069_/a_193_47# control0.count\[0\] 0.00568f
C10847 _0461_ _0582_/a_27_297# 0
C10848 VPWR _0090_ 0.32947f
C10849 _0349_ pp[30] 0.00153f
C10850 _1059_/a_1017_47# acc0.A\[13\] 0.00109f
C10851 _0696_/a_109_297# _0320_ 0
C10852 _0231_ _0600_/a_253_47# 0.02014f
C10853 _0135_ comp0.B\[4\] 0
C10854 _0144_ _0172_ 0.02251f
C10855 _0835_/a_78_199# clkbuf_1_0__f__0465_/a_110_47# 0
C10856 hold10/a_391_47# net125 0
C10857 clkload3/a_268_47# acc0.A\[16\] 0.00119f
C10858 net45 _0710_/a_109_297# 0
C10859 _0125_ acc0.A\[26\] 0
C10860 net58 net141 0
C10861 _0157_ hold82/a_285_47# 0
C10862 hold64/a_49_47# _0217_ 0
C10863 _0488_ _0970_/a_285_47# 0
C10864 _0577_/a_27_297# net150 0.05921f
C10865 _0346_ net72 0
C10866 _0953_/a_114_297# _1061_/a_27_47# 0
C10867 _0846_/a_512_297# acc0.A\[15\] 0
C10868 _0533_/a_373_47# _0171_ 0
C10869 _1001_/a_193_47# _0346_ 0
C10870 net90 _0379_ 0
C10871 VPWR net3 0.25899f
C10872 _0416_ _0399_ 0.10059f
C10873 _0568_/a_109_297# hold62/a_285_47# 0
C10874 _0568_/a_27_297# hold62/a_391_47# 0.01653f
C10875 net243 net110 0.01457f
C10876 _0311_ _0679_/a_150_297# 0
C10877 acc0.A\[22\] _1022_/a_561_413# 0
C10878 _0120_ _1022_/a_1059_315# 0
C10879 _0221_ _0220_ 0
C10880 clknet_1_1__leaf__0458_ _0989_/a_891_413# 0
C10881 _0545_/a_68_297# comp0.B\[9\] 0.17482f
C10882 _0538_/a_149_47# _0143_ 0
C10883 _0201_ net183 0
C10884 _0233_ _0751_/a_111_297# 0
C10885 _0231_ _0751_/a_29_53# 0.0015f
C10886 VPWR _0760_/a_285_47# 0.00163f
C10887 _0524_/a_109_297# net148 0.01104f
C10888 clkbuf_0__0463_/a_110_47# _0175_ 0.00652f
C10889 clknet_1_1__leaf__0463_ net201 0
C10890 net53 _0195_ 0
C10891 _0343_ _0986_/a_466_413# 0
C10892 clknet_1_0__leaf__0459_ _1019_/a_1017_47# 0
C10893 _0299_ A[13] 0
C10894 _0472_ _0563_/a_51_297# 0
C10895 _0326_ _0693_/a_68_297# 0
C10896 _0550_/a_240_47# input30/a_75_212# 0
C10897 _0550_/a_245_297# B[7] 0
C10898 _0259_ _0428_ 0.27725f
C10899 _0982_/a_27_47# net36 0.03372f
C10900 net211 net223 0
C10901 _0259_ _0660_/a_113_47# 0
C10902 net45 _1013_/a_27_47# 0.03323f
C10903 hold26/a_49_47# comp0.B\[9\] 0.32375f
C10904 _0174_ hold51/a_285_47# 0
C10905 _0179_ _1048_/a_27_47# 0.04511f
C10906 _0705_/a_59_75# hold61/a_49_47# 0.00102f
C10907 _0972_/a_250_297# _0972_/a_584_47# 0
C10908 _0401_ _0990_/a_1059_315# 0
C10909 _0290_ _0990_/a_891_413# 0
C10910 _0255_ _0270_ 0
C10911 comp0.B\[15\] net157 0.05044f
C10912 net45 _0607_/a_27_297# 0.01046f
C10913 net36 _0145_ 0.24786f
C10914 hold37/a_391_47# _0172_ 0.00133f
C10915 comp0.B\[12\] net20 0.0475f
C10916 _0278_ _0298_ 0.03245f
C10917 _0993_/a_634_159# _0993_/a_381_47# 0
C10918 A[11] A[12] 0.90888f
C10919 _1058_/a_891_413# _0156_ 0
C10920 net144 _0511_/a_81_21# 0
C10921 net8 net201 0
C10922 hold48/a_285_47# comp0.B\[12\] 0.05901f
C10923 acc0.A\[31\] net99 0.0014f
C10924 _0710_/a_109_297# _0587_/a_27_47# 0
C10925 net102 net219 0
C10926 _1039_/a_466_413# _1039_/a_592_47# 0.00553f
C10927 _1039_/a_634_159# _1039_/a_1017_47# 0
C10928 net185 hold84/a_285_47# 0
C10929 hold67/a_391_47# _0369_ 0.05499f
C10930 _0182_ _0531_/a_373_47# 0
C10931 net203 control0.sh 0
C10932 hold32/a_391_47# acc0.A\[9\] 0.00104f
C10933 _0785_/a_384_47# clknet_0__0465_ 0
C10934 _1039_/a_193_47# _0953_/a_32_297# 0.00129f
C10935 _1038_/a_193_47# _0463_ 0
C10936 _1038_/a_1059_315# clkbuf_0__0463_/a_110_47# 0
C10937 _0483_ hold89/a_391_47# 0
C10938 _0663_/a_207_413# _0287_ 0.06965f
C10939 _0663_/a_27_413# _0293_ 0
C10940 _1056_/a_381_47# net64 0
C10941 input4/a_75_212# net3 0.03317f
C10942 net211 _0982_/a_891_413# 0
C10943 _0172_ _1046_/a_592_47# 0.00147f
C10944 net247 clknet_1_1__leaf__0457_ 1.42196f
C10945 _1032_/a_1059_315# _0215_ 0.01157f
C10946 _0316_ net224 0
C10947 clknet_0__0462_ _0686_/a_27_53# 0.06764f
C10948 _1049_/a_975_413# _0196_ 0
C10949 net135 _0528_/a_81_21# 0
C10950 pp[9] _1055_/a_1059_315# 0
C10951 _1026_/a_634_159# _1026_/a_592_47# 0
C10952 _0985_/a_27_47# _0449_ 0
C10953 clknet_0__0462_ _1008_/a_891_413# 0
C10954 _0985_/a_592_47# clknet_1_0__leaf__0458_ 0
C10955 _0752_/a_27_413# _0103_ 0
C10956 net36 _0446_ 0
C10957 _0343_ _0342_ 0
C10958 net23 control0.reset 0.03981f
C10959 net4 net37 0.04375f
C10960 _0715_/a_27_47# _0259_ 0.00608f
C10961 _0181_ _1009_/a_193_47# 0.02134f
C10962 _0992_/a_1059_315# _0420_ 0
C10963 net224 _0347_ 0
C10964 _0695_/a_80_21# _0324_ 0.06291f
C10965 _1024_/a_891_413# _0122_ 0.00118f
C10966 _1024_/a_381_47# net110 0
C10967 _1024_/a_634_159# acc0.A\[24\] 0
C10968 _0354_ acc0.A\[28\] 0
C10969 _0227_ _0228_ 0.13321f
C10970 _0349_ _0339_ 0.02123f
C10971 hold66/a_49_47# hold66/a_285_47# 0.22264f
C10972 _1014_/a_381_47# _0181_ 0
C10973 _0119_ _1020_/a_27_47# 0
C10974 clknet_1_1__leaf__0464_ net19 0
C10975 _0234_ _0232_ 0.0067f
C10976 _0343_ _0854_/a_79_21# 0.00179f
C10977 net67 _0187_ 0.02172f
C10978 _0105_ net52 0
C10979 _0354_ net209 0
C10980 _1057_/a_1059_315# net143 0
C10981 _0343_ _0334_ 0.01759f
C10982 _1037_/a_27_47# _1037_/a_193_47# 0.96639f
C10983 pp[16] _0997_/a_466_413# 0
C10984 hold89/a_391_47# control0.count\[1\] 0
C10985 hold21/a_285_47# _1054_/a_891_413# 0
C10986 hold21/a_391_47# _1054_/a_1059_315# 0
C10987 _0189_ clknet_1_1__leaf__0465_ 0.09795f
C10988 comp0.B\[2\] net202 0
C10989 VPWR B[13] 0.37776f
C10990 comp0.B\[10\] _1040_/a_27_47# 0.01215f
C10991 acc0.A\[3\] hold71/a_285_47# 0
C10992 _0235_ _0369_ 0
C10993 net189 A[10] 0
C10994 comp0.B\[2\] clknet_1_1__leaf__0463_ 0.08899f
C10995 _0344_ _0220_ 0
C10996 net14 acc0.A\[7\] 0
C10997 _0186_ _0989_/a_193_47# 0
C10998 hold1/a_285_47# _0186_ 0
C10999 clknet_0__0464_ net154 0
C11000 _0957_/a_220_297# net24 0.00189f
C11001 control0.state\[1\] _1067_/a_27_47# 0
C11002 _1020_/a_891_413# _0208_ 0
C11003 clknet_1_0__leaf__0460_ net51 0.15907f
C11004 _0790_/a_35_297# _0790_/a_285_297# 0.02504f
C11005 _0112_ _0345_ 0
C11006 _1068_/a_592_47# _0468_ 0
C11007 _0538_/a_245_297# _0473_ 0.00318f
C11008 _1041_/a_193_47# _1041_/a_381_47# 0.09799f
C11009 _1041_/a_634_159# _1041_/a_891_413# 0.03684f
C11010 _1041_/a_27_47# _1041_/a_561_413# 0.00163f
C11011 _1048_/a_466_413# clknet_1_1__leaf__0457_ 0
C11012 net121 B[1] 0.00328f
C11013 VPWR _0991_/a_466_413# 0.26087f
C11014 hold99/a_285_47# _0993_/a_1059_315# 0.0054f
C11015 clknet_1_0__leaf__0458_ _0426_ 0
C11016 _1017_/a_1059_315# _0219_ 0
C11017 clknet_1_0__leaf__0459_ _0721_/a_27_47# 0.00994f
C11018 _0157_ _0661_/a_27_297# 0
C11019 _0770_/a_79_21# _0244_ 0
C11020 acc0.A\[27\] _0330_ 0.02437f
C11021 net31 _0204_ 0
C11022 _0113_ _0956_/a_32_297# 0
C11023 net33 net17 0
C11024 _0092_ _0404_ 0
C11025 _1002_/a_1059_315# net1 0.00689f
C11026 _0176_ _1043_/a_193_47# 0.00377f
C11027 _0853_/a_68_297# net47 0.10907f
C11028 hold76/a_391_47# _1001_/a_1059_315# 0.01554f
C11029 net234 acc0.A\[1\] 0.26256f
C11030 comp0.B\[2\] net8 0
C11031 net31 hold6/a_391_47# 0
C11032 acc0.A\[12\] _0650_/a_150_297# 0
C11033 _0569_/a_373_47# net114 0
C11034 hold54/a_391_47# VPWR 0.17635f
C11035 _0139_ _0140_ 0.00106f
C11036 net167 net159 0
C11037 acc0.A\[29\] _0723_/a_207_413# 0.08075f
C11038 _0836_/a_68_297# _0218_ 0.17794f
C11039 _1051_/a_193_47# net13 0
C11040 hold86/a_391_47# _0345_ 0.00597f
C11041 _0247_ acc0.A\[19\] 0
C11042 _0305_ net6 0.02077f
C11043 _0707_/a_208_47# _0333_ 0.00506f
C11044 hold12/a_391_47# net17 0
C11045 acc0.A\[16\] clkbuf_1_1__f__0461_/a_110_47# 0.02438f
C11046 net212 _0218_ 0
C11047 comp0.B\[4\] _0160_ 0
C11048 clknet_1_0__leaf__0465_ net169 0
C11049 _0644_/a_285_47# clkbuf_1_1__f__0459_/a_110_47# 0.00305f
C11050 clkbuf_1_0__f__0457_/a_110_47# acc0.A\[19\] 0.00229f
C11051 _0090_ _0283_ 0
C11052 _0195_ _0530_/a_299_297# 0.057f
C11053 _0251_ _0831_/a_35_297# 0.08603f
C11054 hold54/a_49_47# _1015_/a_891_413# 0.00132f
C11055 net53 net90 0.00182f
C11056 VPWR clkbuf_1_0__f__0461_/a_110_47# 1.22781f
C11057 clknet_1_0__leaf__0463_ net28 0
C11058 _0476_ _0955_/a_114_297# 0.00137f
C11059 _0444_ _0084_ 0.00126f
C11060 _0963_/a_35_297# _1069_/a_27_47# 0
C11061 _0259_ _0258_ 0
C11062 _0782_/a_27_47# hold60/a_391_47# 0
C11063 A[12] net66 0.00107f
C11064 _0452_ _0269_ 0
C11065 _0640_/a_215_297# _0254_ 0.19459f
C11066 _0455_ net165 0
C11067 _1013_/a_975_413# net60 0
C11068 VPWR _1025_/a_1017_47# 0.00103f
C11069 input2/a_75_212# _0515_/a_81_21# 0
C11070 _0661_/a_109_297# net67 0.00105f
C11071 _0099_ _0345_ 0.09068f
C11072 _0624_/a_145_75# acc0.A\[4\] 0
C11073 hold69/a_49_47# _0370_ 0.00167f
C11074 _0743_/a_149_47# _0359_ 0.00664f
C11075 _0182_ _0584_/a_109_297# 0.00147f
C11076 _1012_/a_27_47# _0110_ 0.08136f
C11077 _1012_/a_634_159# _0351_ 0
C11078 clknet_1_1__leaf__0460_ net57 0
C11079 _0143_ clkbuf_0__0464_/a_110_47# 0.00497f
C11080 acc0.A\[16\] _0185_ 0.00227f
C11081 hold27/a_49_47# _0172_ 0.05283f
C11082 _0800_/a_240_47# pp[14] 0
C11083 _0472_ _1040_/a_891_413# 0
C11084 _0430_ VPWR 0.50639f
C11085 _1051_/a_891_413# _0523_/a_299_297# 0
C11086 hold66/a_49_47# _0183_ 0
C11087 acc0.A\[18\] clkbuf_0__0457_/a_110_47# 0
C11088 _0216_ _0570_/a_109_47# 0.003f
C11089 _0644_/a_47_47# VPWR 0.30503f
C11090 _0567_/a_27_297# net209 0
C11091 _0254_ _0465_ 0.14045f
C11092 net58 _0831_/a_35_297# 0
C11093 _0421_ _0420_ 0.18659f
C11094 _0359_ _0345_ 0.0503f
C11095 hold99/a_49_47# hold99/a_391_47# 0.00188f
C11096 net18 _1042_/a_1017_47# 0
C11097 _0140_ _1042_/a_561_413# 0.00146f
C11098 VPWR _1044_/a_561_413# 0.00302f
C11099 VPWR _0784_/a_113_47# 0
C11100 _0399_ clkbuf_1_0__f__0465_/a_110_47# 0.00106f
C11101 _0569_/a_109_297# _0106_ 0
C11102 _0519_/a_81_21# _0436_ 0
C11103 VPWR _0401_ 1.51886f
C11104 VPWR acc0.A\[5\] 0.77524f
C11105 _0153_ acc0.A\[9\] 0.38193f
C11106 _0161_ hold84/a_49_47# 0
C11107 _0650_/a_68_297# _0650_/a_150_297# 0.00477f
C11108 clknet_0__0459_ _1059_/a_891_413# 0.0013f
C11109 _0225_ _0600_/a_253_47# 0.00383f
C11110 _1044_/a_27_47# net196 0
C11111 hold35/a_285_47# net2 0
C11112 _0631_/a_109_297# _0261_ 0.00174f
C11113 clkload4/a_110_47# clkload4/Y 0.00568f
C11114 _0470_ hold84/a_391_47# 0.01752f
C11115 _0096_ _0347_ 0.00524f
C11116 _0982_/a_975_413# _0345_ 0
C11117 _1020_/a_1059_315# acc0.A\[21\] 0
C11118 output65/a_27_47# _0435_ 0.00997f
C11119 _0661_/a_27_297# acc0.A\[9\] 0.00239f
C11120 net55 net56 0.02142f
C11121 _0756_/a_129_47# _0378_ 0.00208f
C11122 _0095_ _0400_ 0
C11123 _1001_/a_561_413# _0461_ 0
C11124 _1035_/a_27_47# _0561_/a_240_47# 0
C11125 _1035_/a_1059_315# _0561_/a_51_297# 0.00944f
C11126 _0402_ _0810_/a_113_47# 0
C11127 _0983_/a_193_47# _0264_ 0
C11128 _1027_/a_634_159# net156 0
C11129 _0606_/a_109_53# _0345_ 0.00752f
C11130 _0181_ _1067_/a_1059_315# 0.02301f
C11131 hold8/a_391_47# net113 0
C11132 VPWR _0528_/a_299_297# 0.28363f
C11133 VPWR net222 0.32157f
C11134 net101 _1019_/a_466_413# 0
C11135 _0710_/a_109_297# VPWR 0.12768f
C11136 output47/a_27_47# pp[1] 0.33776f
C11137 clknet_1_0__leaf__0462_ _1023_/a_891_413# 0.00358f
C11138 clknet_0__0460_ _0321_ 0
C11139 clknet_1_1__leaf__0460_ _0125_ 0.00163f
C11140 _0751_/a_29_53# _0225_ 0.30546f
C11141 _0197_ _0449_ 0.0018f
C11142 clknet_1_0__leaf__0464_ _1061_/a_891_413# 0.00217f
C11143 net119 comp0.B\[6\] 0
C11144 _0757_/a_68_297# net50 0.05254f
C11145 clkbuf_0__0460_/a_110_47# clknet_0__0460_ 1.8786f
C11146 _0634_/a_113_47# clknet_1_0__leaf__0461_ 0
C11147 net176 _0350_ 0
C11148 _1052_/a_27_47# _1052_/a_634_159# 0.13832f
C11149 _1032_/a_193_47# _0113_ 0
C11150 net202 _1015_/a_193_47# 0
C11151 _0478_ _1071_/a_27_47# 0.08919f
C11152 control0.reset _1063_/a_466_413# 0
C11153 acc0.A\[12\] acc0.A\[15\] 0.06465f
C11154 acc0.A\[27\] net190 0.02873f
C11155 _1035_/a_1059_315# _0133_ 0.06563f
C11156 _1035_/a_891_413# net121 0
C11157 _0390_ clkbuf_1_0__f__0461_/a_110_47# 0.00158f
C11158 _0248_ _0764_/a_384_47# 0
C11159 _1058_/a_193_47# _1058_/a_466_413# 0.07482f
C11160 _1058_/a_27_47# _1058_/a_1059_315# 0.04861f
C11161 _0450_ _0843_/a_150_297# 0
C11162 _0891_/a_27_47# _0208_ 0.05485f
C11163 _0186_ net142 0.02818f
C11164 hold69/a_285_47# _0350_ 0.0418f
C11165 hold10/a_285_47# _0499_/a_59_75# 0
C11166 _0195_ clkbuf_1_1__f__0462_/a_110_47# 0
C11167 _1051_/a_891_413# _0172_ 0.05567f
C11168 _0809_/a_81_21# _0420_ 0.11301f
C11169 _0172_ _1045_/a_561_413# 0
C11170 VPWR _0182_ 1.56234f
C11171 _0983_/a_466_413# _0082_ 0
C11172 net69 _0849_/a_79_21# 0
C11173 _0211_ clknet_0__0463_ 0
C11174 _0558_/a_68_297# _1035_/a_1059_315# 0.00179f
C11175 _0451_ _0219_ 0.00165f
C11176 _1050_/a_27_47# _0527_/a_109_297# 0
C11177 _1050_/a_193_47# _0527_/a_27_297# 0.00104f
C11178 _0680_/a_80_21# _0680_/a_300_47# 0.00997f
C11179 _0680_/a_217_297# _0680_/a_472_297# 0.00517f
C11180 _0310_ _0780_/a_285_297# 0.05413f
C11181 acc0.A\[30\] _0333_ 0
C11182 _0718_/a_47_47# _0349_ 0.14379f
C11183 _0718_/a_129_47# _0337_ 0.0031f
C11184 _0725_/a_209_297# hold62/a_285_47# 0
C11185 _0725_/a_80_21# hold62/a_391_47# 0
C11186 acc0.A\[29\] net191 0.07475f
C11187 _1011_/a_193_47# _0355_ 0.04107f
C11188 _1011_/a_27_47# net227 0.00207f
C11189 _1011_/a_634_159# _0354_ 0.00537f
C11190 _0462_ _0773_/a_35_297# 0
C11191 VPWR _1013_/a_27_47# 0.68612f
C11192 _0983_/a_27_47# clknet_1_0__leaf__0458_ 0.01121f
C11193 net32 _1043_/a_891_413# 0
C11194 _0139_ _1043_/a_634_159# 0
C11195 _0598_/a_79_21# clknet_1_0__leaf__0460_ 0
C11196 _0607_/a_27_297# VPWR 0.2152f
C11197 _1052_/a_1059_315# net148 0.00218f
C11198 _1052_/a_193_47# net12 0.03386f
C11199 net190 _0364_ 0
C11200 _0642_/a_215_297# _0434_ 0.01391f
C11201 control0.sh _0176_ 0.58924f
C11202 _0617_/a_68_297# _0350_ 0
C11203 _0174_ _0935_/a_27_47# 0
C11204 _0113_ _0721_/a_27_47# 0
C11205 _0174_ _1061_/a_193_47# 0.00173f
C11206 _0477_ _1065_/a_27_47# 0
C11207 net125 _1061_/a_1017_47# 0
C11208 _0443_ VPWR 0.71727f
C11209 acc0.A\[9\] _0990_/a_27_47# 0
C11210 acc0.A\[22\] _0183_ 0.74082f
C11211 net150 _0120_ 0
C11212 comp0.B\[10\] _1061_/a_466_413# 0
C11213 _0195_ _1018_/a_381_47# 0.01273f
C11214 _1027_/a_634_159# acc0.A\[26\] 0
C11215 net156 _1026_/a_891_413# 0
C11216 hold68/a_49_47# _0350_ 0
C11217 net58 _0988_/a_381_47# 0.00437f
C11218 hold77/a_391_47# _0347_ 0
C11219 _0467_ _1067_/a_561_413# 0
C11220 _0297_ _0405_ 0.12928f
C11221 _0128_ hold62/a_391_47# 0.05487f
C11222 hold97/a_391_47# _0319_ 0
C11223 _0195_ _1049_/a_1059_315# 0.00405f
C11224 _0181_ net6 0.10948f
C11225 comp0.B\[10\] net171 0
C11226 _1038_/a_466_413# _0176_ 0.01696f
C11227 net89 clkbuf_0_clk/a_110_47# 0
C11228 _0563_/a_240_47# _0208_ 0.02679f
C11229 _0214_ _0173_ 0.18032f
C11230 net228 _0345_ 0.04554f
C11231 clknet_1_0__leaf__0465_ _0464_ 0.01584f
C11232 net211 clkbuf_0__0457_/a_110_47# 0.00661f
C11233 output45/a_27_47# _0340_ 0
C11234 hold59/a_391_47# net206 0.18737f
C11235 _0530_/a_299_297# _1048_/a_193_47# 0
C11236 net205 _1034_/a_27_47# 0
C11237 _0996_/a_466_413# clkbuf_0__0459_/a_110_47# 0
C11238 clknet_1_0__leaf__0462_ _0312_ 0.00202f
C11239 _0985_/a_27_47# _0260_ 0
C11240 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0461_/a_110_47# 0.05608f
C11241 acc0.A\[12\] _0179_ 0.0349f
C11242 net9 net170 0.01562f
C11243 _0994_/a_27_47# _0218_ 0.03959f
C11244 net59 _1012_/a_466_413# 0
C11245 _0403_ _0993_/a_634_159# 0
C11246 _0195_ acc0.A\[17\] 0.15644f
C11247 _0948_/a_109_297# clkbuf_0_clk/a_110_47# 0
C11248 _0239_ _0307_ 0
C11249 clknet_0__0462_ _0320_ 0.00121f
C11250 comp0.B\[11\] net195 0
C11251 net73 _0193_ 0.00125f
C11252 _0995_/a_466_413# pp[14] 0.00194f
C11253 _0579_/a_27_297# net105 0
C11254 _0412_ _0405_ 0.01725f
C11255 net46 _0223_ 0.00231f
C11256 _0520_/a_109_297# net14 0.01461f
C11257 _0538_/a_149_47# _0174_ 0.02166f
C11258 _0346_ _0208_ 0
C11259 VPWR _1042_/a_634_159# 0.17966f
C11260 _1056_/a_27_47# acc0.A\[9\] 0.04071f
C11261 _1018_/a_975_413# _0247_ 0
C11262 _0397_ _0240_ 0
C11263 _1028_/a_193_47# _1008_/a_27_47# 0
C11264 net55 _0345_ 0
C11265 _0154_ net66 0.00101f
C11266 _0518_/a_27_297# net65 0
C11267 _0397_ _0369_ 0
C11268 _0395_ _0347_ 0.29766f
C11269 _0998_/a_27_47# net83 0
C11270 _0463_ net29 0
C11271 clknet_0__0460_ _1009_/a_27_47# 0
C11272 _0343_ _0240_ 0.03366f
C11273 acc0.A\[8\] acc0.A\[6\] 0.15644f
C11274 _0255_ _0085_ 0
C11275 _0426_ _0288_ 0.00432f
C11276 pp[27] _1030_/a_891_413# 0.00118f
C11277 _0373_ _0219_ 0.02903f
C11278 _0988_/a_27_47# _0988_/a_466_413# 0.27314f
C11279 _0988_/a_193_47# _0988_/a_634_159# 0.11897f
C11280 _0343_ _0369_ 0.30563f
C11281 control0.reset _0213_ 0
C11282 _1039_/a_193_47# _0174_ 0
C11283 _0984_/a_1059_315# _0983_/a_27_47# 0
C11284 _0671_/a_113_297# _0670_/a_79_21# 0
C11285 net157 _0176_ 0
C11286 _0998_/a_27_47# _0781_/a_68_297# 0
C11287 _0730_/a_79_21# _0357_ 0.05894f
C11288 _0369_ net95 0
C11289 _0580_/a_27_297# _0117_ 0.13492f
C11290 _0304_ _0347_ 0.68536f
C11291 _0359_ net52 0
C11292 _0195_ net60 0
C11293 net10 _1043_/a_891_413# 0.01961f
C11294 clkbuf_1_0__f__0457_/a_110_47# net1 0
C11295 hold20/a_285_47# _0490_ 0
C11296 hold20/a_49_47# net167 0
C11297 _0953_/a_32_297# _0953_/a_114_297# 0.01439f
C11298 _0315_ _0319_ 0
C11299 hold21/a_391_47# hold22/a_285_47# 0.00676f
C11300 _0343_ hold96/a_285_47# 0
C11301 _0542_/a_51_297# _0542_/a_149_47# 0.02487f
C11302 _0967_/a_215_297# _1064_/a_891_413# 0.00229f
C11303 hold96/a_49_47# _0575_/a_27_297# 0
C11304 _0162_ _1064_/a_1059_315# 0.00202f
C11305 _0485_ _1064_/a_561_413# 0
C11306 hold52/a_285_47# net200 0
C11307 _0207_ _0173_ 0
C11308 _1026_/a_891_413# acc0.A\[26\] 0.00352f
C11309 hold94/a_285_47# net51 0.00258f
C11310 _0465_ _1047_/a_975_413# 0
C11311 _0224_ _0592_/a_150_297# 0
C11312 _0999_/a_27_47# _0396_ 0
C11313 _0880_/a_27_47# _1062_/a_193_47# 0
C11314 _0329_ _0324_ 0.00825f
C11315 _0356_ _0725_/a_303_47# 0
C11316 VPWR _0562_/a_150_297# 0.002f
C11317 _0817_/a_81_21# _0424_ 0.08848f
C11318 _0416_ _0091_ 0
C11319 clknet_1_1__leaf__0460_ _1009_/a_891_413# 0.01556f
C11320 _0242_ _0771_/a_298_297# 0
C11321 clknet_1_0__leaf__0458_ acc0.A\[3\] 0
C11322 clknet_1_1__leaf__0458_ _0988_/a_1059_315# 0
C11323 _0324_ clknet_1_0__leaf__0460_ 0.0034f
C11324 A[2] net10 0
C11325 net110 acc0.A\[24\] 0
C11326 net195 _0202_ 0
C11327 _0141_ _0540_/a_149_47# 0
C11328 input6/a_75_212# output40/a_27_47# 0.00124f
C11329 _0401_ _0283_ 0.02819f
C11330 _0982_/a_634_159# hold60/a_49_47# 0
C11331 _0982_/a_27_47# hold60/a_391_47# 0
C11332 _0982_/a_193_47# hold60/a_285_47# 0
C11333 pp[26] _0571_/a_373_47# 0
C11334 output54/a_27_47# acc0.A\[27\] 0.04902f
C11335 net153 _1040_/a_193_47# 0.00104f
C11336 net59 net98 0
C11337 _0787_/a_80_21# _0787_/a_209_47# 0.01013f
C11338 hold47/a_285_47# net154 0.00331f
C11339 acc0.A\[0\] _0181_ 0.02304f
C11340 _0461_ _0614_/a_111_297# 0
C11341 _0230_ _0377_ 0.04305f
C11342 _0273_ _0087_ 0
C11343 _0792_/a_80_21# _0345_ 0.00858f
C11344 _0471_ _0161_ 0
C11345 net9 _0525_/a_81_21# 0
C11346 _0174_ _1040_/a_592_47# 0
C11347 _1037_/a_466_413# _1037_/a_592_47# 0.00553f
C11348 _1037_/a_634_159# _1037_/a_1017_47# 0
C11349 net101 _0352_ 0.00251f
C11350 net200 net52 0
C11351 output36/a_27_47# input30/a_75_212# 0
C11352 _0997_/a_193_47# _0218_ 0.00195f
C11353 VPWR hold70/a_49_47# 0.26228f
C11354 _0195_ _0998_/a_634_159# 0.0111f
C11355 _0183_ _0379_ 0
C11356 _0387_ _0462_ 0
C11357 _0557_/a_240_47# _0209_ 0
C11358 pp[30] _1030_/a_193_47# 0.03667f
C11359 A[4] A[7] 0
C11360 clknet_0__0459_ acc0.A\[16\] 0
C11361 VPWR _1005_/a_561_413# 0.00579f
C11362 net42 acc0.A\[15\] 2.0559f
C11363 _1039_/a_1059_315# _0173_ 0
C11364 _0427_ net62 0
C11365 VPWR _0089_ 0.35105f
C11366 _0985_/a_193_47# _0447_ 0
C11367 _0985_/a_1059_315# _0844_/a_297_47# 0
C11368 net234 _0854_/a_297_297# 0
C11369 net54 _0360_ 0
C11370 _0228_ _0352_ 0
C11371 clkbuf_1_1__f__0462_/a_110_47# _1010_/a_891_413# 0
C11372 _1054_/a_592_47# _0180_ 0.00274f
C11373 _1016_/a_27_47# _0219_ 0
C11374 output66/a_27_47# _0186_ 0
C11375 _1001_/a_193_47# _1001_/a_634_159# 0.12126f
C11376 _1001_/a_27_47# _1001_/a_466_413# 0.27314f
C11377 net64 acc0.A\[6\] 0.85565f
C11378 _0621_/a_117_297# acc0.A\[6\] 0
C11379 _0607_/a_27_297# clknet_1_0__leaf__0459_ 0
C11380 net23 _0460_ 0
C11381 net233 _0843_/a_68_297# 0
C11382 _1062_/a_27_47# _1062_/a_193_47# 0.9705f
C11383 _0217_ hold40/a_391_47# 0.00569f
C11384 _0183_ hold40/a_49_47# 0
C11385 _0717_/a_209_47# _0333_ 0.00408f
C11386 VPWR _0765_/a_510_47# 0
C11387 _1039_/a_1017_47# _0473_ 0
C11388 hold9/a_391_47# _1008_/a_891_413# 0
C11389 clknet_1_0__leaf__0458_ _0851_/a_113_47# 0
C11390 _0831_/a_35_297# _0831_/a_285_297# 0.02504f
C11391 _0963_/a_35_297# _0489_ 0.04398f
C11392 _0275_ _0817_/a_266_47# 0
C11393 _0146_ _0531_/a_109_297# 0.00222f
C11394 _1049_/a_1059_315# _1048_/a_193_47# 0
C11395 _1049_/a_891_413# _1048_/a_27_47# 0.0012f
C11396 hold8/a_285_47# hold8/a_391_47# 0.41909f
C11397 hold14/a_285_47# _1037_/a_27_47# 0
C11398 _0287_ net37 0
C11399 _0376_ _0369_ 0
C11400 hold54/a_391_47# _0113_ 0
C11401 _0967_/a_215_297# hold84/a_49_47# 0
C11402 _0967_/a_109_93# hold84/a_285_47# 0
C11403 VPWR _1006_/a_891_413# 0.21201f
C11404 _0457_ net23 0.0401f
C11405 _0222_ hold29/a_49_47# 0.00374f
C11406 _0279_ _0346_ 0
C11407 _1000_/a_27_47# _0217_ 0
C11408 _0326_ _0743_/a_51_297# 0
C11409 clkload1/Y _0256_ 0
C11410 _1055_/a_891_413# A[10] 0
C11411 net45 _0781_/a_150_297# 0
C11412 _0195_ _1030_/a_561_413# 0.00175f
C11413 net48 _1005_/a_561_413# 0
C11414 pp[8] net47 0.00174f
C11415 net35 _0460_ 0
C11416 _0328_ _0460_ 0
C11417 VPWR _0986_/a_891_413# 0.20841f
C11418 _1046_/a_634_159# _1061_/a_27_47# 0
C11419 _0550_/a_240_47# _0176_ 0.00698f
C11420 _0714_/a_245_297# _0219_ 0.00156f
C11421 _1019_/a_1017_47# _0345_ 0.00139f
C11422 pp[9] _1058_/a_466_413# 0
C11423 _0260_ _0197_ 0
C11424 VPWR _0495_/a_68_297# 0.16955f
C11425 clknet_1_0__leaf__0465_ _0830_/a_79_21# 0
C11426 _0951_/a_209_311# _0951_/a_368_53# 0.0026f
C11427 _1013_/a_466_413# _0567_/a_27_297# 0
C11428 _0701_/a_209_47# _0332_ 0
C11429 _0186_ _0988_/a_27_47# 0
C11430 _1004_/a_634_159# _0216_ 0.01695f
C11431 _0161_ hold93/a_391_47# 0
C11432 clknet_1_0__leaf__0457_ clknet_1_0__leaf__0461_ 0.05041f
C11433 acc0.A\[5\] _0523_/a_81_21# 0
C11434 _0561_/a_51_297# _0561_/a_245_297# 0.01218f
C11435 VPWR _0616_/a_78_199# 0.27372f
C11436 net145 clknet_1_1__leaf__0465_ 0.27823f
C11437 _0218_ _0411_ 0.03806f
C11438 _1072_/a_634_159# _1068_/a_193_47# 0
C11439 _1072_/a_193_47# _1068_/a_634_159# 0
C11440 _1072_/a_466_413# _1068_/a_27_47# 0
C11441 _1072_/a_27_47# _1068_/a_466_413# 0
C11442 _0180_ _0522_/a_373_47# 0.00139f
C11443 _0515_/a_81_21# _0514_/a_27_297# 0
C11444 _0689_/a_150_297# _0319_ 0
C11445 _0339_ clknet_1_1__leaf__0461_ 0
C11446 _0174_ clkbuf_0__0464_/a_110_47# 0.00257f
C11447 acc0.A\[18\] _0350_ 0
C11448 comp0.B\[13\] _0538_/a_149_47# 0.00629f
C11449 _0502_/a_27_47# _0551_/a_27_47# 0
C11450 _0316_ _0329_ 0.02525f
C11451 _0289_ _0288_ 0.82697f
C11452 _0293_ acc0.A\[9\] 0.19429f
C11453 net165 _0448_ 0
C11454 _0538_/a_51_297# _1046_/a_1059_315# 0
C11455 _0461_ net223 0.00838f
C11456 _1035_/a_634_159# _0132_ 0
C11457 _1035_/a_1059_315# _0208_ 0.00126f
C11458 _0133_ _0561_/a_245_297# 0
C11459 _0272_ _0275_ 0.19042f
C11460 _0236_ _0377_ 0
C11461 _0238_ _0345_ 0.00284f
C11462 net47 _1060_/a_27_47# 0
C11463 _1047_/a_634_159# _1047_/a_466_413# 0.23992f
C11464 _1047_/a_193_47# _1047_/a_1059_315# 0.03405f
C11465 _1047_/a_27_47# _1047_/a_891_413# 0.03224f
C11466 _0985_/a_1059_315# clknet_0__0458_ 0
C11467 _1030_/a_193_47# _0339_ 0.01837f
C11468 _0206_ _1040_/a_381_47# 0.01651f
C11469 hold1/a_391_47# _0987_/a_193_47# 0.00644f
C11470 acc0.A\[13\] net229 0.00393f
C11471 _0185_ _0506_/a_299_297# 0.00323f
C11472 _0329_ _0347_ 0.02206f
C11473 _0957_/a_32_297# _0475_ 0.14247f
C11474 _0957_/a_114_297# _0472_ 0.0045f
C11475 _0957_/a_304_297# _0473_ 0
C11476 _0464_ net137 0
C11477 _0714_/a_51_297# _0129_ 0
C11478 net101 net207 0.00123f
C11479 _0137_ _0463_ 0.02132f
C11480 net47 _0988_/a_891_413# 0.00445f
C11481 clknet_1_0__leaf__0460_ hold3/a_391_47# 0
C11482 net62 net142 0
C11483 clknet_1_0__leaf__0460_ _0347_ 0.06501f
C11484 _1041_/a_1059_315# _0174_ 0.06782f
C11485 _0323_ _0352_ 0
C11486 pp[28] _0726_/a_51_297# 0
C11487 _0582_/a_27_297# _0115_ 0.1119f
C11488 net234 _1014_/a_634_159# 0
C11489 _0797_/a_27_413# acc0.A\[13\] 0
C11490 net178 _0517_/a_299_297# 0.06479f
C11491 _1052_/a_891_413# _1052_/a_975_413# 0.00851f
C11492 _1052_/a_381_47# _1052_/a_561_413# 0.00123f
C11493 _1007_/a_634_159# _1007_/a_592_47# 0
C11494 _1001_/a_1059_315# clknet_1_0__leaf__0461_ 0
C11495 control0.reset _0161_ 0
C11496 net67 clknet_1_1__leaf__0465_ 0.96718f
C11497 hold96/a_391_47# _1004_/a_634_159# 0
C11498 hold96/a_285_47# _1004_/a_466_413# 0.00148f
C11499 VPWR _0854_/a_215_47# 0.00236f
C11500 _0177_ _1061_/a_466_413# 0.00175f
C11501 _0195_ net175 0.43392f
C11502 net240 hold93/a_49_47# 0
C11503 _1058_/a_891_413# _1058_/a_1017_47# 0.00617f
C11504 _1058_/a_634_159# net144 0
C11505 _0172_ _1044_/a_381_47# 0.02194f
C11506 hold69/a_391_47# _1006_/a_193_47# 0
C11507 _0416_ _0346_ 0
C11508 _0179_ _1052_/a_381_47# 0.01665f
C11509 _0502_/a_27_47# _0533_/a_27_297# 0
C11510 _1020_/a_466_413# _0352_ 0.00135f
C11511 net197 _1027_/a_193_47# 0
C11512 _1021_/a_193_47# clknet_1_0__leaf__0461_ 0
C11513 _0104_ clknet_1_0__leaf__0460_ 0.00347f
C11514 net63 _0434_ 0
C11515 net44 _0110_ 0
C11516 VPWR net31 0.23033f
C11517 _0557_/a_51_297# VPWR 0.44621f
C11518 clknet_1_1__leaf__0461_ net6 0
C11519 _0635_/a_109_297# _0265_ 0.01031f
C11520 _1050_/a_466_413# net11 0.00306f
C11521 _0258_ _0446_ 0
C11522 _0500_/a_27_47# _0181_ 0.0052f
C11523 net185 B[15] 0
C11524 hold32/a_285_47# output47/a_27_47# 0
C11525 _0305_ _0311_ 0.09554f
C11526 _1003_/a_634_159# _0487_ 0
C11527 control0.state\[0\] _0951_/a_109_93# 0
C11528 _0669_/a_29_53# net41 0
C11529 _0971_/a_299_297# _0971_/a_384_47# 0
C11530 _0954_/a_32_297# _0140_ 0
C11531 comp0.B\[11\] _0204_ 0
C11532 _0568_/a_27_297# _0334_ 0
C11533 _0353_ net209 0
C11534 net97 _0354_ 0.00103f
C11535 _1011_/a_975_413# _0109_ 0
C11536 net57 _0726_/a_240_47# 0
C11537 clk control0.count\[0\] 0.00194f
C11538 _0216_ _0726_/a_245_297# 0.00101f
C11539 _1018_/a_193_47# _0580_/a_27_297# 0
C11540 _1033_/a_466_413# control0.reset 0.00699f
C11541 _0268_ _0345_ 0.04597f
C11542 _1002_/a_592_47# VPWR 0
C11543 _0309_ _0307_ 0
C11544 _0558_/a_68_297# _0558_/a_150_297# 0.00477f
C11545 hold21/a_285_47# A[7] 0
C11546 _1061_/a_193_47# comp0.B\[9\] 0
C11547 _0182_ _0113_ 0
C11548 _0469_ clknet_0_clk 0.03153f
C11549 clkbuf_0_clk/a_110_47# _1063_/a_634_159# 0
C11550 net61 _0989_/a_634_159# 0.00157f
C11551 hold46/a_49_47# net174 0
C11552 hold59/a_49_47# _0350_ 0
C11553 _0924_/a_27_47# _0180_ 0.00204f
C11554 clkbuf_1_0__f__0462_/a_110_47# hold90/a_285_47# 0.01986f
C11555 hold75/a_285_47# net222 0.00997f
C11556 hold40/a_49_47# hold40/a_285_47# 0.22264f
C11557 _0983_/a_193_47# _0454_ 0.00529f
C11558 _0983_/a_27_47# _0455_ 0.08914f
C11559 _0617_/a_150_297# _1006_/a_193_47# 0
C11560 _0761_/a_113_47# _0219_ 0
C11561 _0283_ hold70/a_49_47# 0
C11562 net169 _0519_/a_299_297# 0
C11563 _1063_/a_27_47# _1063_/a_1059_315# 0.04875f
C11564 _1063_/a_193_47# _1063_/a_466_413# 0.07482f
C11565 _0090_ _0345_ 0.00144f
C11566 _1058_/a_381_47# _0186_ 0
C11567 _0645_/a_377_297# acc0.A\[15\] 0
C11568 _0770_/a_297_47# clkbuf_1_0__f__0457_/a_110_47# 0
C11569 _0975_/a_59_75# control0.state\[2\] 0.09951f
C11570 _0463_ comp0.B\[6\] 0.0014f
C11571 _1019_/a_193_47# _0346_ 0.0343f
C11572 _1037_/a_193_47# _0208_ 0
C11573 _1037_/a_1059_315# _0173_ 0
C11574 net159 _1063_/a_27_47# 0
C11575 _0788_/a_150_297# _0403_ 0.00178f
C11576 _0786_/a_217_297# _0402_ 0.00271f
C11577 _1063_/a_891_413# clknet_1_0__leaf__0457_ 0.00172f
C11578 _0462_ _1006_/a_27_47# 0.00513f
C11579 net172 _0176_ 0.04905f
C11580 net203 _0474_ 0
C11581 _0974_/a_448_47# net159 0.05738f
C11582 _1039_/a_466_413# _0177_ 0
C11583 hold58/a_285_47# comp0.B\[2\] 0
C11584 hold52/a_49_47# _1025_/a_27_47# 0
C11585 hold85/a_49_47# _1062_/a_27_47# 0.01003f
C11586 _0536_/a_51_297# clknet_0__0464_ 0
C11587 control0.state\[2\] net231 0
C11588 net63 acc0.A\[7\] 0.06253f
C11589 _0984_/a_592_47# VPWR 0
C11590 _0172_ _0205_ 0.09064f
C11591 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# 1.67709f
C11592 _0820_/a_79_21# net66 0.00218f
C11593 net211 _0350_ 0.00566f
C11594 hold19/a_49_47# _0459_ 0.00359f
C11595 _1004_/a_1059_315# net90 0
C11596 _0354_ _0707_/a_201_297# 0
C11597 _0355_ _0707_/a_75_199# 0
C11598 _1011_/a_1059_315# acc0.A\[29\] 0.02752f
C11599 net14 _0186_ 0.00224f
C11600 _1004_/a_634_159# _1024_/a_193_47# 0
C11601 net197 _1026_/a_1059_315# 0
C11602 _1004_/a_466_413# _1024_/a_27_47# 0
C11603 _1004_/a_27_47# _1024_/a_466_413# 0
C11604 _1004_/a_193_47# _1024_/a_634_159# 0
C11605 _0369_ _0990_/a_381_47# 0
C11606 _0732_/a_80_21# _0315_ 0.00527f
C11607 _0732_/a_209_297# _0366_ 0.01823f
C11608 _0217_ net165 0.16938f
C11609 VPWR net128 0.34032f
C11610 _0476_ comp0.B\[4\] 0.37476f
C11611 VPWR _0704_/a_150_297# 0.00161f
C11612 _0343_ _0409_ 0
C11613 _1060_/a_27_47# _1060_/a_1059_315# 0.04875f
C11614 _1060_/a_193_47# _1060_/a_466_413# 0.07482f
C11615 _0204_ _0202_ 0.00407f
C11616 _0191_ net65 0
C11617 clkbuf_1_0__f__0459_/a_110_47# _0369_ 0.16231f
C11618 pp[26] _0216_ 0.23429f
C11619 _1039_/a_193_47# comp0.B\[9\] 0
C11620 VPWR _0384_ 0.48559f
C11621 _0143_ _1050_/a_193_47# 0
C11622 _0325_ net52 0.01244f
C11623 _1012_/a_27_47# _0097_ 0
C11624 hold47/a_285_47# clknet_0__0464_ 0
C11625 _0805_/a_27_47# clknet_1_1__leaf__0459_ 0.03197f
C11626 hold56/a_49_47# _1065_/a_891_413# 0
C11627 hold56/a_285_47# _1065_/a_1059_315# 0
C11628 _0988_/a_193_47# net74 0.01355f
C11629 _0988_/a_1059_315# _0988_/a_1017_47# 0
C11630 _0467_ _0971_/a_81_21# 0.18057f
C11631 _0856_/a_215_47# _0456_ 0.00837f
C11632 _0787_/a_209_47# _0402_ 0
C11633 _1067_/a_27_47# clknet_1_1__leaf_clk 0.24765f
C11634 net46 _0216_ 0.03564f
C11635 _0968_/a_109_297# control0.state\[0\] 0
C11636 _1053_/a_891_413# acc0.A\[7\] 0.00297f
C11637 clk _1062_/a_466_413# 0
C11638 _0358_ _0108_ 0.0012f
C11639 comp0.B\[14\] net174 0
C11640 _0315_ clkbuf_1_0__f__0460_/a_110_47# 0
C11641 _0320_ _0687_/a_59_75# 0.01331f
C11642 _0217_ acc0.A\[19\] 0.2151f
C11643 _1041_/a_193_47# _0206_ 0
C11644 _1041_/a_634_159# comp0.B\[8\] 0
C11645 _0982_/a_891_413# _0465_ 0.00269f
C11646 _0953_/a_304_297# comp0.B\[10\] 0.00326f
C11647 _0753_/a_297_297# _0378_ 0
C11648 clknet_1_0__leaf__0463_ clknet_0__0463_ 0.01439f
C11649 _0606_/a_109_53# hold94/a_391_47# 0
C11650 VPWR _1014_/a_466_413# 0.2512f
C11651 _1071_/a_27_47# VPWR 0.66399f
C11652 _0542_/a_240_47# net19 0.0663f
C11653 _0109_ _0334_ 0
C11654 _0315_ _0250_ 0
C11655 _0998_/a_891_413# _0779_/a_79_21# 0
C11656 clknet_1_0__leaf__0465_ _0826_/a_301_297# 0
C11657 _1001_/a_1017_47# clknet_1_0__leaf__0457_ 0
C11658 clkbuf_1_0__f__0463_/a_110_47# net29 0.00153f
C11659 _0172_ _1042_/a_193_47# 0
C11660 _0467_ _0164_ 0
C11661 _0820_/a_79_21# _0350_ 0
C11662 hold14/a_391_47# net121 0.061f
C11663 _0238_ net52 0.0053f
C11664 _0216_ _0584_/a_109_47# 0.00145f
C11665 _1035_/a_1017_47# net27 0
C11666 _1021_/a_561_413# clknet_1_0__leaf__0457_ 0
C11667 _1021_/a_891_413# _0460_ 0.00638f
C11668 _0327_ hold95/a_285_47# 0
C11669 _0343_ pp[31] 0.00109f
C11670 _0701_/a_209_297# _0701_/a_303_47# 0
C11671 hold46/a_49_47# clknet_0__0464_ 0
C11672 comp0.B\[13\] clkbuf_0__0464_/a_110_47# 0
C11673 _0244_ acc0.A\[18\] 0.23607f
C11674 net133 _1047_/a_891_413# 0
C11675 net23 net27 0.00164f
C11676 clknet_1_1__leaf__0462_ _0687_/a_145_75# 0
C11677 _1001_/a_27_47# _0241_ 0
C11678 net36 _0269_ 0
C11679 _1067_/a_193_47# clkbuf_1_1__f_clk/a_110_47# 0.01336f
C11680 _0257_ _0270_ 0.0049f
C11681 _0992_/a_27_47# net143 0
C11682 clkbuf_0__0464_/a_110_47# _1046_/a_193_47# 0.02274f
C11683 hold73/a_49_47# hold73/a_391_47# 0.00188f
C11684 net48 _0384_ 0
C11685 _1050_/a_466_413# clknet_1_1__leaf__0458_ 0
C11686 hold79/a_285_47# _0167_ 0
C11687 hold79/a_391_47# clknet_1_0__leaf_clk 0.06721f
C11688 _0275_ _0181_ 0.10199f
C11689 _1008_/a_891_413# _0739_/a_215_47# 0
C11690 _0959_/a_80_21# _0561_/a_240_47# 0
C11691 _0400_ _0219_ 0.17514f
C11692 A[11] _0511_/a_81_21# 0
C11693 _0144_ _1061_/a_1059_315# 0
C11694 _0536_/a_240_47# net147 0
C11695 _0228_ _0237_ 0.15399f
C11696 _0999_/a_27_47# net43 0
C11697 _1037_/a_592_47# _0135_ 0.00164f
C11698 net175 _1048_/a_193_47# 0.00386f
C11699 _0996_/a_1059_315# hold91/a_285_47# 0.0054f
C11700 _0195_ net84 0.02418f
C11701 _0179_ _0440_ 0
C11702 _0596_/a_145_75# VPWR 0
C11703 hold25/a_391_47# _1038_/a_27_47# 0.01134f
C11704 hold25/a_285_47# _1038_/a_193_47# 0.01156f
C11705 hold25/a_49_47# _1038_/a_634_159# 0
C11706 VPWR _0781_/a_150_297# 0.00191f
C11707 _0221_ hold95/a_49_47# 0
C11708 _0538_/a_51_297# _1045_/a_634_159# 0
C11709 _0635_/a_109_297# _0267_ 0
C11710 clknet_1_1__leaf__0459_ _0779_/a_215_47# 0
C11711 _0467_ hold38/a_391_47# 0
C11712 clkbuf_1_0__f__0462_/a_110_47# clknet_0__0462_ 0.32336f
C11713 output59/a_27_47# _0568_/a_27_297# 0
C11714 clknet_1_1__leaf__0460_ _0680_/a_217_297# 0
C11715 _0311_ _0181_ 0
C11716 hold45/a_49_47# net3 0
C11717 _0728_/a_145_75# _0356_ 0.00145f
C11718 hold9/a_285_47# net113 0
C11719 _0188_ acc0.A\[10\] 0.00222f
C11720 net58 _0451_ 0.00367f
C11721 _0993_/a_27_47# net38 0.00455f
C11722 pp[28] VPWR 0.5114f
C11723 hold13/a_49_47# _0133_ 0
C11724 _0470_ net23 0.02685f
C11725 _0172_ _0562_/a_68_297# 0
C11726 hold30/a_285_47# acc0.A\[23\] 0
C11727 VPWR _0679_/a_68_297# 0.19909f
C11728 _1001_/a_466_413# _0772_/a_79_21# 0
C11729 _1001_/a_193_47# _0772_/a_215_47# 0
C11730 _1001_/a_1059_315# _1001_/a_1017_47# 0
C11731 acc0.A\[21\] acc0.A\[20\] 0.10739f
C11732 net234 net247 0
C11733 _0991_/a_466_413# _0345_ 0
C11734 hold47/a_49_47# clknet_1_0__leaf__0464_ 0.00987f
C11735 _1035_/a_634_159# net25 0
C11736 _0136_ _0957_/a_32_297# 0
C11737 _1062_/a_466_413# _1062_/a_592_47# 0.00553f
C11738 _1062_/a_634_159# _1062_/a_1017_47# 0
C11739 net17 _0880_/a_27_47# 0.00775f
C11740 _0302_ clkbuf_1_1__f__0459_/a_110_47# 0.03866f
C11741 net132 _0527_/a_27_297# 0
C11742 _1011_/a_634_159# _0353_ 0
C11743 net130 net13 0
C11744 _0992_/a_891_413# net228 0
C11745 hold38/a_391_47# comp0.B\[0\] 0
C11746 _1021_/a_634_159# _1021_/a_381_47# 0
C11747 _1033_/a_193_47# net23 0
C11748 _1003_/a_975_413# net49 0
C11749 net61 _0258_ 0.25665f
C11750 net199 _1024_/a_634_159# 0.00787f
C11751 hold41/a_285_47# net188 0.00833f
C11752 _0091_ net246 0.00482f
C11753 _0854_/a_215_47# _0453_ 0
C11754 _1056_/a_975_413# _0186_ 0
C11755 _1017_/a_193_47# _0459_ 0.00495f
C11756 _0147_ _1048_/a_634_159# 0
C11757 _1049_/a_466_413# net134 0.00631f
C11758 _0576_/a_27_297# _0757_/a_68_297# 0.00183f
C11759 net53 acc0.A\[26\] 0.0217f
C11760 _0102_ acc0.A\[23\] 0
C11761 _0607_/a_109_47# _0399_ 0
C11762 _0346_ clkbuf_1_0__f__0465_/a_110_47# 0
C11763 _0732_/a_80_21# _0742_/a_81_21# 0.00201f
C11764 _0645_/a_47_47# _0645_/a_285_47# 0.01755f
C11765 _0510_/a_27_297# _0510_/a_109_47# 0.00393f
C11766 _0996_/a_1059_315# _0670_/a_215_47# 0
C11767 acc0.A\[31\] _0708_/a_68_297# 0.17862f
C11768 comp0.B\[14\] clknet_0__0464_ 0.03911f
C11769 hold59/a_49_47# _0244_ 0
C11770 hold15/a_49_47# net60 0.00161f
C11771 hold64/a_391_47# net45 0
C11772 _0667_/a_113_47# net5 0
C11773 _0733_/a_79_199# _0733_/a_222_93# 0.22112f
C11774 _0218_ clknet_1_0__leaf__0457_ 0.02134f
C11775 _0481_ clknet_1_0__leaf_clk 0.11926f
C11776 _0857_/a_27_47# net17 0.00584f
C11777 net62 _0988_/a_27_47# 0.00576f
C11778 net194 _0143_ 0.16191f
C11779 VPWR _0548_/a_240_47# 0.00764f
C11780 hold98/a_49_47# net42 0
C11781 _0181_ _0583_/a_27_297# 0
C11782 _0241_ _0459_ 0.01818f
C11783 net65 clkbuf_1_0__f__0465_/a_110_47# 0
C11784 hold87/a_49_47# net36 0.32415f
C11785 clkbuf_1_0__f__0465_/a_110_47# _0989_/a_466_413# 0
C11786 _0294_ _1060_/a_27_47# 0.01074f
C11787 _1031_/a_634_159# _1013_/a_27_47# 0
C11788 _1031_/a_27_47# _1013_/a_634_159# 0
C11789 control0.state\[0\] _0486_ 0.24423f
C11790 control0.state\[1\] control0.state\[2\] 0.2886f
C11791 clkbuf_1_0__f__0461_/a_110_47# _0345_ 0
C11792 clknet_1_1__leaf__0464_ _1043_/a_975_413# 0
C11793 _0376_ _0756_/a_47_47# 0
C11794 _0195_ _0568_/a_109_297# 0.05373f
C11795 _1046_/a_27_47# net147 0
C11796 _0195_ _1015_/a_381_47# 0
C11797 _0248_ acc0.A\[19\] 0.08241f
C11798 _0996_/a_193_47# _0369_ 0
C11799 net118 control0.add 0.00134f
C11800 _1034_/a_634_159# clknet_0__0463_ 0
C11801 _0799_/a_80_21# net41 0
C11802 hold26/a_285_47# net152 0
C11803 _0742_/a_81_21# clkbuf_1_0__f__0460_/a_110_47# 0
C11804 _0343_ _0084_ 0.00234f
C11805 hold38/a_391_47# _1034_/a_634_159# 0
C11806 hold38/a_285_47# _1034_/a_466_413# 0
C11807 _0657_/a_109_297# _0181_ 0
C11808 _0225_ _1022_/a_891_413# 0
C11809 hold17/a_49_47# _1071_/a_193_47# 0.00284f
C11810 hold17/a_285_47# _1071_/a_27_47# 0
C11811 _0984_/a_27_47# _0399_ 0
C11812 hold78/a_49_47# net225 0
C11813 net46 _1024_/a_193_47# 0
C11814 _0750_/a_27_47# _0460_ 0.00274f
C11815 _0561_/a_240_47# _0173_ 0.01301f
C11816 _0717_/a_209_297# net44 0
C11817 VPWR _1067_/a_193_47# 0.32684f
C11818 hold100/a_391_47# _0261_ 0.03393f
C11819 hold100/a_285_47# _0263_ 0.0468f
C11820 _1072_/a_27_47# _0166_ 0
C11821 hold90/a_391_47# _0105_ 0
C11822 VPWR _0383_ 0.53558f
C11823 _0461_ clkbuf_0__0457_/a_110_47# 0.00414f
C11824 _0488_ _0468_ 0
C11825 net17 _1062_/a_27_47# 0
C11826 net53 _0733_/a_222_93# 0
C11827 _0119_ net23 0
C11828 _0515_/a_81_21# _0189_ 0.17213f
C11829 _0515_/a_384_47# net2 0
C11830 _0228_ _1005_/a_27_47# 0.00136f
C11831 VPWR input18/a_75_212# 0.28627f
C11832 pp[17] _0338_ 0
C11833 A[11] net181 0
C11834 _0982_/a_466_413# _0261_ 0
C11835 _0982_/a_634_159# _0263_ 0
C11836 output55/a_27_47# acc0.A\[29\] 0.01716f
C11837 _0640_/a_109_53# _0271_ 0.11686f
C11838 clkbuf_0__0461_/a_110_47# _0240_ 0.00339f
C11839 _1020_/a_466_413# net106 0
C11840 net149 net47 0
C11841 _0869_/a_27_47# _0391_ 0
C11842 _0180_ net71 0
C11843 _0475_ _0213_ 0.02891f
C11844 _0472_ _0173_ 0.04531f
C11845 _0369_ clkbuf_0__0461_/a_110_47# 0.02256f
C11846 hold39/a_391_47# _0175_ 0.03028f
C11847 _1036_/a_592_47# clknet_1_1__leaf__0463_ 0
C11848 hold14/a_49_47# hold14/a_285_47# 0.22264f
C11849 _0346_ _0792_/a_209_47# 0
C11850 _0389_ _0771_/a_27_413# 0.00144f
C11851 _0510_/a_109_47# _0181_ 0
C11852 _0461_ _1019_/a_561_413# 0
C11853 _0538_/a_512_297# net132 0
C11854 _0401_ _0345_ 0.0555f
C11855 _0401_ _0814_/a_27_47# 0.23524f
C11856 VPWR _0852_/a_285_47# 0
C11857 _0423_ _0814_/a_181_47# 0
C11858 _0644_/a_285_47# _0296_ 0
C11859 _1001_/a_1059_315# _0218_ 0.01459f
C11860 _0248_ _0249_ 0.05591f
C11861 comp0.B\[15\] _0563_/a_51_297# 0
C11862 net121 _0132_ 0
C11863 _1041_/a_1059_315# comp0.B\[9\] 0.08396f
C11864 _1041_/a_561_413# net153 0
C11865 _0350_ _1008_/a_193_47# 0.00126f
C11866 _1047_/a_634_159# _0145_ 0.02004f
C11867 _0329_ _0106_ 0
C11868 hold12/a_285_47# _0237_ 0
C11869 hold12/a_391_47# _0381_ 0
C11870 hold1/a_49_47# _0085_ 0
C11871 hold1/a_285_47# net73 0
C11872 net186 clknet_1_1__leaf_clk 0
C11873 net225 _0129_ 0
C11874 net181 _0744_/a_27_47# 0
C11875 clkbuf_1_1__f__0459_/a_110_47# net6 0
C11876 net222 _0345_ 0
C11877 net125 _1046_/a_27_47# 0
C11878 _0973_/a_27_297# net107 0
C11879 _0725_/a_80_21# _0334_ 0.00251f
C11880 _0710_/a_109_297# _0345_ 0
C11881 _0474_ _0176_ 0.14383f
C11882 net188 _0513_/a_384_47# 0.01006f
C11883 hold41/a_285_47# _0155_ 0
C11884 _0217_ _1018_/a_975_413# 0
C11885 _0109_ _0724_/a_113_297# 0
C11886 B[5] _0175_ 0
C11887 _1004_/a_27_47# _0756_/a_285_47# 0
C11888 net190 _0689_/a_68_297# 0
C11889 net58 _0271_ 0
C11890 _0464_ _0148_ 0
C11891 _0536_/a_240_47# _0473_ 0.00605f
C11892 net10 _0545_/a_68_297# 0
C11893 net243 _1004_/a_975_413# 0
C11894 clknet_1_1__leaf__0460_ _0372_ 0.0197f
C11895 _0101_ _0373_ 0
C11896 _0440_ _0441_ 0.14193f
C11897 _0805_/a_109_47# _0281_ 0
C11898 _0118_ _0352_ 0.35458f
C11899 _0502_/a_27_47# _0199_ 0
C11900 _0305_ _0677_/a_285_47# 0.00492f
C11901 net48 _0383_ 0.04732f
C11902 B[11] net19 0.00886f
C11903 _0217_ _0575_/a_109_47# 0.00282f
C11904 VPWR net7 1.49726f
C11905 hold42/a_285_47# net37 0.02944f
C11906 _0350_ _0611_/a_150_297# 0
C11907 control0.sh net28 0.07375f
C11908 _0535_/a_68_297# _0535_/a_150_297# 0.00477f
C11909 _1057_/a_1059_315# net37 0.01511f
C11910 _0732_/a_209_297# acc0.A\[24\] 0.00235f
C11911 clknet_1_0__leaf__0459_ _0781_/a_150_297# 0.00145f
C11912 _0734_/a_377_297# _0362_ 0.00514f
C11913 _0137_ clkbuf_1_0__f__0463_/a_110_47# 0.04782f
C11914 _0217_ net1 0.06463f
C11915 acc0.A\[4\] net154 0.02449f
C11916 _1034_/a_27_47# _1034_/a_193_47# 0.96968f
C11917 net89 _0487_ 0.18808f
C11918 _0183_ acc0.A\[17\] 0
C11919 _0796_/a_79_21# _0796_/a_215_47# 0.04584f
C11920 hold26/a_49_47# net10 0
C11921 net162 _1030_/a_27_47# 0
C11922 _0181_ _0163_ 0.00606f
C11923 _0128_ _0334_ 0
C11924 net168 _1053_/a_27_47# 0
C11925 hold10/a_49_47# comp0.B\[15\] 0.29448f
C11926 _0131_ control0.reset 0
C11927 _0782_/a_27_47# _0208_ 0.21954f
C11928 _0993_/a_27_47# _0282_ 0
C11929 net64 _0826_/a_219_297# 0.01008f
C11930 _0608_/a_27_47# VPWR 0.00489f
C11931 _0380_ net109 0
C11932 _1057_/a_381_47# net67 0.004f
C11933 _0819_/a_384_47# acc0.A\[8\] 0
C11934 _0428_ _0659_/a_68_297# 0
C11935 hold25/a_49_47# _0550_/a_149_47# 0
C11936 _0982_/a_634_159# clknet_1_0__leaf__0461_ 0.00118f
C11937 hold64/a_285_47# net234 0
C11938 _1038_/a_466_413# net28 0
C11939 _1013_/a_27_47# _0345_ 0.00877f
C11940 _0983_/a_592_47# _0081_ 0
C11941 _0617_/a_68_297# net92 0.00936f
C11942 _0755_/a_109_297# _0374_ 0.00239f
C11943 VPWR _0825_/a_150_297# 0.0014f
C11944 acc0.A\[12\] clknet_1_1__leaf__0459_ 0.2989f
C11945 _0517_/a_81_21# _0181_ 0
C11946 net45 _0678_/a_68_297# 0
C11947 _1063_/a_891_413# _1063_/a_1017_47# 0.00617f
C11948 _1063_/a_193_47# _0161_ 0.64539f
C11949 _0224_ _0756_/a_47_47# 0
C11950 hold69/a_49_47# _0369_ 0
C11951 VPWR _0844_/a_297_47# 0.00354f
C11952 _0968_/a_193_297# _1068_/a_27_47# 0
C11953 net204 _0207_ 0
C11954 hold64/a_285_47# net46 0
C11955 hold74/a_391_47# _0507_/a_109_297# 0
C11956 hold100/a_49_47# _0265_ 0.00106f
C11957 hold100/a_391_47# net47 0
C11958 acc0.A\[1\] hold2/a_285_47# 0.07865f
C11959 VPWR _1024_/a_634_159# 0.18285f
C11960 _0443_ _0345_ 0.01836f
C11961 _0161_ _0460_ 0.00532f
C11962 net203 _0563_/a_51_297# 0.1227f
C11963 _0982_/a_193_47# _0265_ 0
C11964 _0956_/a_32_297# net24 0
C11965 clknet_1_0__leaf__0464_ _1050_/a_891_413# 0
C11966 _0172_ B[8] 0
C11967 _0748_/a_384_47# _0294_ 0.01011f
C11968 _0235_ _0374_ 0
C11969 _0349_ _1012_/a_466_413# 0.00544f
C11970 net17 net107 0
C11971 VPWR _1048_/a_1059_315# 0.40797f
C11972 pp[30] _0567_/a_27_297# 0
C11973 _0183_ net5 0.06388f
C11974 net158 net135 0
C11975 _1028_/a_381_47# net113 0
C11976 _0434_ _0824_/a_59_75# 0
C11977 _1055_/a_634_159# acc0.A\[8\] 0
C11978 _0305_ _0114_ 0
C11979 VPWR net229 0.151f
C11980 _0601_/a_68_297# _0223_ 0
C11981 _0642_/a_298_297# _0253_ 0.00464f
C11982 hold47/a_49_47# hold47/a_391_47# 0.00188f
C11983 _0809_/a_299_297# net228 0.01362f
C11984 hold13/a_49_47# _0174_ 0
C11985 net181 net66 0.09993f
C11986 _0473_ _1046_/a_27_47# 0.00629f
C11987 comp0.B\[6\] clkbuf_1_0__f__0463_/a_110_47# 0
C11988 _0354_ _0339_ 0.04437f
C11989 net235 clknet_1_1__leaf__0458_ 0
C11990 _0216_ _0569_/a_373_47# 0.00287f
C11991 _0500_/a_27_47# _0531_/a_27_297# 0.00901f
C11992 net190 net112 0
C11993 _1004_/a_27_47# _0122_ 0
C11994 VPWR _1010_/a_975_413# 0.00489f
C11995 _1000_/a_634_159# _1000_/a_381_47# 0
C11996 _1033_/a_891_413# clknet_1_0__leaf__0457_ 0
C11997 _0715_/a_27_47# _0659_/a_68_297# 0
C11998 _1060_/a_891_413# _1060_/a_1017_47# 0.00617f
C11999 _1060_/a_193_47# _0158_ 0.17294f
C12000 _1060_/a_634_159# net146 0
C12001 VPWR _0797_/a_27_413# 0.24467f
C12002 _1051_/a_466_413# net154 0.01166f
C12003 _1051_/a_27_47# net11 0.0015f
C12004 _0168_ _0979_/a_109_47# 0
C12005 _0192_ net168 0
C12006 _0462_ _0247_ 0.00131f
C12007 _1072_/a_634_159# VPWR 0.18621f
C12008 VPWR _0841_/a_297_297# 0.00738f
C12009 _0362_ clknet_0__0462_ 0
C12010 _1039_/a_1059_315# net204 0
C12011 clkbuf_1_0__f__0457_/a_110_47# _0462_ 0.01227f
C12012 _0953_/a_114_297# comp0.B\[9\] 0.00116f
C12013 clkbuf_0__0459_/a_110_47# _0219_ 0.08809f
C12014 _0329_ _1011_/a_27_47# 0
C12015 _0553_/a_240_47# _0136_ 0.04658f
C12016 _0399_ _0986_/a_561_413# 0
C12017 _0352_ _0320_ 0.16372f
C12018 net207 hold60/a_285_47# 0.01976f
C12019 _0252_ clkbuf_1_1__f__0458_/a_110_47# 0.00609f
C12020 net105 hold60/a_391_47# 0.02986f
C12021 hold8/a_49_47# hold9/a_391_47# 0
C12022 _0698_/a_113_297# _0330_ 0.09722f
C12023 clknet_1_1__leaf__0459_ _0650_/a_68_297# 0.01257f
C12024 hold14/a_285_47# _0208_ 0.00129f
C12025 VPWR _1009_/a_592_47# 0
C12026 clknet_0__0457_ net87 0.03123f
C12027 _0312_ _1006_/a_27_47# 0
C12028 clknet_1_0__leaf__0458_ hold59/a_391_47# 0
C12029 _0457_ _1033_/a_466_413# 0
C12030 _0346_ _0824_/a_145_75# 0.00165f
C12031 _0537_/a_68_297# comp0.B\[12\] 0.0157f
C12032 _0233_ _0379_ 0
C12033 _0161_ _1062_/a_891_413# 0.00264f
C12034 _0979_/a_27_297# clkbuf_1_0__f_clk/a_110_47# 0
C12035 clknet_1_0__leaf__0462_ hold4/a_391_47# 0.02294f
C12036 net240 clknet_1_0__leaf__0457_ 0.00127f
C12037 _1050_/a_27_47# _1050_/a_193_47# 0.97021f
C12038 net81 _0407_ 0
C12039 _0719_/a_27_47# _0391_ 0
C12040 _0959_/a_217_297# _0160_ 0.05148f
C12041 net58 pp[2] 0.01515f
C12042 clknet_1_0__leaf__0457_ _0099_ 0.0015f
C12043 acc0.A\[15\] net5 0.03412f
C12044 clknet_1_1__leaf__0462_ _0739_/a_510_47# 0
C12045 clkload1/a_110_47# _0432_ 0
C12046 hold74/a_49_47# clknet_1_1__leaf__0461_ 0.02233f
C12047 acc0.A\[21\] net107 0
C12048 _0221_ _1011_/a_27_47# 0.38841f
C12049 net67 _0808_/a_81_21# 0
C12050 _0256_ _0261_ 0
C12051 _1018_/a_634_159# _0181_ 0
C12052 _0179_ _1049_/a_1059_315# 0.05692f
C12053 _0819_/a_81_21# _0401_ 0.05696f
C12054 clknet_0__0458_ _0439_ 0
C12055 _0778_/a_150_297# _0347_ 0
C12056 _0181_ _1049_/a_27_47# 0
C12057 _0999_/a_634_159# _1012_/a_27_47# 0
C12058 hold86/a_391_47# _0635_/a_27_47# 0
C12059 B[4] input17/a_75_212# 0
C12060 clknet_0__0458_ VPWR 2.562f
C12061 _0458_ _0631_/a_109_297# 0
C12062 _0858_/a_27_47# _0263_ 0
C12063 hold25/a_285_47# net29 0
C12064 _0578_/a_27_297# clknet_1_0__leaf__0460_ 0.00956f
C12065 _0222_ _0754_/a_149_47# 0.0193f
C12066 clknet_1_1__leaf__0460_ net244 0.13246f
C12067 _0997_/a_1059_315# net41 0.04469f
C12068 _0997_/a_634_159# pp[14] 0
C12069 _0836_/a_68_297# acc0.A\[5\] 0.0424f
C12070 _1071_/a_1059_315# clknet_0_clk 0.00198f
C12071 _1008_/a_975_413# _0106_ 0.00175f
C12072 net54 _1027_/a_561_413# 0.00137f
C12073 _0313_ _0322_ 0.06078f
C12074 clknet_1_1__leaf__0465_ net6 0.28276f
C12075 VPWR comp0.B\[11\] 0.78178f
C12076 _0257_ _0085_ 0
C12077 hold13/a_49_47# _0208_ 0
C12078 _0212_ net27 0.01562f
C12079 _0305_ clkload3/Y 0.00246f
C12080 _0585_/a_373_47# _0208_ 0
C12081 net1 _0971_/a_81_21# 0
C12082 acc0.A\[5\] net212 0
C12083 hold64/a_391_47# VPWR 0.16154f
C12084 _0337_ _1030_/a_891_413# 0
C12085 _0349_ _1030_/a_466_413# 0
C12086 _0258_ _0431_ 0.66216f
C12087 _0538_/a_51_297# _1044_/a_193_47# 0
C12088 net9 _1048_/a_592_47# 0.00112f
C12089 _0314_ clknet_1_0__leaf__0460_ 0
C12090 _0313_ _0327_ 0
C12091 _0577_/a_109_297# VPWR 0.19343f
C12092 net46 _0756_/a_377_297# 0.00148f
C12093 control0.state\[2\] _1066_/a_634_159# 0
C12094 acc0.A\[14\] _1060_/a_193_47# 0.00385f
C12095 _1020_/a_27_47# net187 0
C12096 _1000_/a_27_47# _1018_/a_891_413# 0
C12097 _1000_/a_193_47# _1018_/a_1059_315# 0
C12098 control0.state\[2\] _1068_/a_634_159# 0
C12099 _0486_ _1068_/a_193_47# 0.06158f
C12100 _0143_ _1045_/a_27_47# 0.00177f
C12101 net21 _1045_/a_466_413# 0.01387f
C12102 net44 _0097_ 0.15594f
C12103 net149 _1047_/a_1017_47# 0
C12104 net3 _0156_ 0
C12105 hold70/a_49_47# _0345_ 0.00489f
C12106 clkload4/Y net103 0.07202f
C12107 VPWR _1022_/a_1017_47# 0
C12108 net59 net208 0
C12109 _0251_ clknet_1_0__leaf__0465_ 0
C12110 net123 _0552_/a_68_297# 0
C12111 _0343_ _1000_/a_27_47# 0.03053f
C12112 _0246_ clknet_1_0__leaf__0461_ 0
C12113 _1033_/a_27_47# _0173_ 0.00514f
C12114 output39/a_27_47# _0218_ 0.00252f
C12115 _0235_ _0249_ 0
C12116 _0852_/a_285_47# _0453_ 0
C12117 _0610_/a_59_75# _0242_ 0.11257f
C12118 _0978_/a_27_297# _0976_/a_505_21# 0
C12119 _0537_/a_150_297# _0202_ 0
C12120 _0999_/a_634_159# _0999_/a_592_47# 0
C12121 net17 _1063_/a_561_413# 0
C12122 _0339_ _0567_/a_27_297# 0.01737f
C12123 _0720_/a_68_297# _0352_ 0.01721f
C12124 _1001_/a_466_413# _1019_/a_27_47# 0
C12125 _1001_/a_193_47# _1019_/a_634_159# 0
C12126 _1001_/a_27_47# _1019_/a_466_413# 0
C12127 _1017_/a_891_413# _0115_ 0
C12128 _0772_/a_297_297# _0772_/a_215_47# 0
C12129 _0772_/a_79_21# _0772_/a_510_47# 0.00844f
C12130 _0754_/a_51_297# _0103_ 0.10355f
C12131 _0731_/a_81_21# _0219_ 0.00173f
C12132 _0583_/a_27_297# clknet_1_1__leaf__0461_ 0
C12133 _1001_/a_1059_315# _0099_ 0
C12134 VPWR _0993_/a_634_159# 0.18703f
C12135 _1054_/a_27_47# net148 0
C12136 _1016_/a_27_47# _0582_/a_109_297# 0
C12137 _0478_ _0486_ 0
C12138 _0089_ _0345_ 0.18229f
C12139 clknet_1_0__leaf__0462_ _1007_/a_634_159# 0.0134f
C12140 net1 _0164_ 0
C12141 net121 net25 0
C12142 net233 _0263_ 0
C12143 _0534_/a_299_297# _0465_ 0.00651f
C12144 _0369_ acc0.A\[6\] 0.08772f
C12145 _0983_/a_27_47# _0217_ 0
C12146 hold47/a_285_47# comp0.B\[14\] 0.00397f
C12147 _1020_/a_891_413# net202 0
C12148 _0695_/a_80_21# _0360_ 0
C12149 net191 clknet_1_1__leaf__0462_ 0.0032f
C12150 _1043_/a_193_47# _0542_/a_51_297# 0
C12151 hold100/a_49_47# _0267_ 0
C12152 _0311_ _0098_ 0
C12153 _1021_/a_891_413# _0119_ 0.00117f
C12154 _0094_ _1060_/a_1059_315# 0
C12155 net199 net110 0
C12156 _0558_/a_68_297# B[2] 0
C12157 clknet_0__0461_ _0308_ 0
C12158 _0147_ net134 0.09712f
C12159 _0130_ net23 0.00804f
C12160 net188 net4 0.02567f
C12161 _0999_/a_193_47# clknet_1_1__leaf__0461_ 0
C12162 _0732_/a_303_47# _0368_ 0.00306f
C12163 net168 A[5] 0
C12164 clknet_1_1__leaf__0459_ net42 0.15099f
C12165 _0577_/a_109_297# net48 0
C12166 _0324_ hold90/a_285_47# 0
C12167 _0359_ hold90/a_391_47# 0.0562f
C12168 VPWR _0202_ 0.72448f
C12169 _0510_/a_109_47# _0187_ 0
C12170 control0.count\[2\] _0979_/a_27_297# 0.03138f
C12171 clknet_1_0__leaf__0465_ hold7/a_49_47# 0.01662f
C12172 _1017_/a_634_159# _0218_ 0
C12173 _1051_/a_27_47# clknet_1_1__leaf__0458_ 0.0014f
C12174 _1043_/a_1059_315# net20 0
C12175 _0181_ _0114_ 0
C12176 _0181_ _0615_/a_109_297# 0
C12177 _0222_ _0228_ 0
C12178 _1011_/a_381_47# _0219_ 0.00611f
C12179 hold88/a_285_47# _0254_ 0
C12180 _0375_ _0618_/a_79_21# 0.04514f
C12181 _1006_/a_193_47# _0219_ 0
C12182 _0656_/a_145_75# _0345_ 0
C12183 hold12/a_391_47# _0468_ 0
C12184 clknet_1_0__leaf__0459_ net229 0
C12185 _0804_/a_79_21# _0218_ 0
C12186 acc0.A\[12\] _0655_/a_215_53# 0
C12187 _0751_/a_111_297# _0219_ 0
C12188 _0467_ _1068_/a_466_413# 0
C12189 _0518_/a_27_297# _0518_/a_109_297# 0.17136f
C12190 _0217_ _0225_ 0
C12191 _0614_/a_29_53# _0614_/a_183_297# 0.00868f
C12192 _0461_ _0773_/a_285_297# 0.00132f
C12193 comp0.B\[10\] _0206_ 0.30822f
C12194 _0424_ _0426_ 0.07313f
C12195 _0985_/a_193_47# _0985_/a_466_413# 0.07855f
C12196 _0985_/a_27_47# _0985_/a_1059_315# 0.04875f
C12197 net194 _0174_ 0
C12198 hold46/a_49_47# comp0.B\[14\] 0.12277f
C12199 _0368_ clknet_0__0460_ 0
C12200 acc0.A\[25\] _0219_ 0.00297f
C12201 _0780_/a_117_297# _0397_ 0
C12202 _1018_/a_27_47# _1018_/a_634_159# 0.13601f
C12203 clknet_1_0__leaf__0465_ net183 0.00412f
C12204 _0985_/a_27_47# _1049_/a_193_47# 0
C12205 _0985_/a_193_47# _1049_/a_27_47# 0
C12206 _0404_ _0670_/a_79_21# 0
C12207 net178 _0439_ 0
C12208 net50 _1022_/a_193_47# 0
C12209 _0642_/a_298_297# _0642_/a_382_47# 0
C12210 net194 _1050_/a_27_47# 0
C12211 hold47/a_391_47# _1050_/a_891_413# 0
C12212 _0280_ _0285_ 0
C12213 hold29/a_49_47# net151 0
C12214 net178 VPWR 0.40382f
C12215 _0275_ _0990_/a_193_47# 0
C12216 A[4] net11 0.00735f
C12217 net62 _0267_ 0
C12218 acc0.A\[29\] acc0.A\[30\] 0
C12219 _0254_ _0086_ 0.00633f
C12220 _0195_ acc0.A\[18\] 0.08764f
C12221 _0267_ _0450_ 1.06476f
C12222 _0080_ _0261_ 0.00278f
C12223 _0524_/a_27_297# _0522_/a_27_297# 0
C12224 _0582_/a_109_47# net206 0
C12225 _1019_/a_466_413# _0459_ 0
C12226 _0145_ _0208_ 0
C12227 _0118_ net106 0.00136f
C12228 net11 _0085_ 0.00319f
C12229 net68 _1047_/a_27_47# 0
C12230 _0461_ _0350_ 0.03576f
C12231 _0530_/a_299_297# _0530_/a_384_47# 0
C12232 hold44/a_49_47# _0195_ 0
C12233 _0780_/a_35_297# acc0.A\[17\] 0.00308f
C12234 acc0.A\[4\] clknet_0__0464_ 0
C12235 VPWR _0756_/a_129_47# 0
C12236 _0172_ clknet_1_1__leaf__0464_ 1.15995f
C12237 _0734_/a_129_47# _0359_ 0
C12238 _0172_ _0548_/a_149_47# 0.00272f
C12239 VPWR _1027_/a_381_47# 0.07652f
C12240 _0143_ net132 0.01771f
C12241 net204 _1037_/a_1059_315# 0
C12242 _0350_ _0318_ 0
C12243 hold79/a_49_47# hold79/a_285_47# 0.22264f
C12244 VPWR _0749_/a_81_21# 0.20435f
C12245 net170 _0843_/a_68_297# 0
C12246 acc0.A\[14\] _0796_/a_79_21# 0
C12247 net89 _0760_/a_47_47# 0
C12248 net17 _0208_ 0.08466f
C12249 _0997_/a_634_159# _0408_ 0
C12250 VPWR _0678_/a_68_297# 0.17288f
C12251 _0179_ acc0.A\[11\] 0.11975f
C12252 _1056_/a_634_159# acc0.A\[10\] 0.02851f
C12253 _0459_ net219 0.03142f
C12254 clkbuf_0_clk/a_110_47# _0487_ 0.0426f
C12255 VPWR _0766_/a_109_297# 0.00502f
C12256 net63 _0186_ 0.11792f
C12257 net109 _1005_/a_891_413# 0
C12258 _1042_/a_466_413# hold51/a_391_47# 0
C12259 _0176_ _0563_/a_51_297# 0
C12260 _0165_ net107 0.00876f
C12261 net45 _0675_/a_68_297# 0.00902f
C12262 net116 _0352_ 0
C12263 _0399_ _1014_/a_891_413# 0
C12264 _0487_ _1063_/a_634_159# 0
C12265 _0205_ _1040_/a_193_47# 0
C12266 _1019_/a_1059_315# clknet_1_0__leaf__0461_ 0
C12267 clkbuf_1_1__f_clk/a_110_47# _0951_/a_109_93# 0
C12268 comp0.B\[10\] _1046_/a_1059_315# 0
C12269 net178 output62/a_27_47# 0
C12270 _0584_/a_109_297# clkbuf_1_1__f__0457_/a_110_47# 0
C12271 _1004_/a_891_413# _0379_ 0.00912f
C12272 _0731_/a_81_21# _0746_/a_81_21# 0.00143f
C12273 _0155_ net4 0.01894f
C12274 _0343_ _0374_ 0
C12275 hold54/a_285_47# _0214_ 0
C12276 net44 net162 0
C12277 pp[17] acc0.A\[31\] 0.31558f
C12278 _0346_ _0991_/a_891_413# 0
C12279 clkload3/Y _0181_ 0
C12280 _0994_/a_466_413# net80 0
C12281 _0176_ _0541_/a_68_297# 0.14292f
C12282 hold78/a_49_47# _0340_ 0.00883f
C12283 hold78/a_285_47# _0341_ 0.06162f
C12284 _0544_/a_245_297# net198 0.00153f
C12285 _0544_/a_149_47# _0204_ 0.00154f
C12286 _0544_/a_51_297# net18 0.10616f
C12287 net175 acc0.A\[15\] 0
C12288 hold64/a_391_47# clknet_1_0__leaf__0459_ 0
C12289 _0274_ _0433_ 0.04796f
C12290 net10 hold51/a_285_47# 0.03793f
C12291 _0217_ control0.sh 0
C12292 B[0] net17 0.00369f
C12293 net216 _0460_ 0.1457f
C12294 _1058_/a_891_413# net143 0
C12295 _0637_/a_311_297# _0263_ 0
C12296 _1034_/a_466_413# _1034_/a_592_47# 0.00553f
C12297 _1034_/a_634_159# _1034_/a_1017_47# 0
C12298 _0536_/a_240_47# _0200_ 0
C12299 hold6/a_285_47# _0544_/a_240_47# 0.0014f
C12300 _0513_/a_81_21# acc0.A\[11\] 0.00349f
C12301 _0452_ acc0.A\[0\] 0
C12302 _0343_ _0507_/a_27_297# 0.0032f
C12303 _0497_/a_150_297# _0177_ 0
C12304 _0607_/a_27_297# _0394_ 0
C12305 _1021_/a_592_47# acc0.A\[21\] 0
C12306 _0559_/a_240_47# net205 0.04211f
C12307 net67 _0811_/a_81_21# 0
C12308 _0258_ _0269_ 0.00634f
C12309 _0891_/a_27_47# net202 0.11211f
C12310 net48 _0749_/a_81_21# 0
C12311 hold59/a_49_47# _0195_ 0
C12312 net68 clknet_1_0__leaf__0461_ 0.09244f
C12313 hold25/a_285_47# _0137_ 0
C12314 _0640_/a_297_297# clknet_0__0465_ 0
C12315 net172 net28 0
C12316 _0627_/a_109_93# VPWR 0.09829f
C12317 net16 acc0.A\[9\] 0.15767f
C12318 _1013_/a_561_413# _0219_ 0
C12319 hold36/a_391_47# comp0.B\[12\] 0
C12320 _0570_/a_109_297# net190 0.01052f
C12321 _0343_ net165 0.03873f
C12322 _0230_ _0460_ 0
C12323 hold10/a_49_47# _0176_ 0
C12324 _0842_/a_59_75# _0084_ 0
C12325 _0129_ _0340_ 0.30135f
C12326 VPWR _1026_/a_592_47# 0
C12327 _0324_ clknet_0__0462_ 0.36109f
C12328 net34 net1 0
C12329 _0483_ _1072_/a_975_413# 0
C12330 control0.count\[3\] _1072_/a_1017_47# 0
C12331 net206 net47 0.18694f
C12332 _0470_ _0161_ 0.01364f
C12333 hold78/a_285_47# _1013_/a_891_413# 0.01623f
C12334 hold78/a_391_47# _1013_/a_1059_315# 0.00277f
C12335 _0344_ _1013_/a_193_47# 0
C12336 hold29/a_49_47# _0378_ 0
C12337 VPWR _0817_/a_368_297# 0.00183f
C12338 _0549_/a_68_297# _0176_ 0.13763f
C12339 acc0.A\[20\] net105 0
C12340 comp0.B\[14\] _0543_/a_68_297# 0.00195f
C12341 _1001_/a_27_47# _0352_ 0.00444f
C12342 _0793_/a_512_297# net42 0
C12343 VPWR net110 0.62326f
C12344 hold27/a_391_47# net147 0.00523f
C12345 _0172_ net247 0.00254f
C12346 net30 net7 0
C12347 _0517_/a_299_297# _0153_ 0.05025f
C12348 _1018_/a_466_413# _0242_ 0
C12349 _0559_/a_149_47# _0211_ 0
C12350 _1071_/a_466_413# _0488_ 0
C12351 _1071_/a_634_159# _0466_ 0.00552f
C12352 _0080_ net47 0
C12353 net58 net76 0
C12354 hold8/a_49_47# _0739_/a_215_47# 0
C12355 _0770_/a_297_47# _0248_ 0.00135f
C12356 net81 _0995_/a_193_47# 0.00436f
C12357 _0993_/a_193_47# _0286_ 0
C12358 _0227_ net51 0.41364f
C12359 hold77/a_49_47# _1009_/a_193_47# 0
C12360 hold77/a_285_47# _1009_/a_27_47# 0
C12361 net18 _0141_ 0
C12362 clknet_1_0__leaf__0460_ _1005_/a_975_413# 0
C12363 _1050_/a_27_47# _0987_/a_193_47# 0
C12364 _1050_/a_193_47# _0987_/a_27_47# 0
C12365 _0343_ acc0.A\[19\] 0
C12366 _1017_/a_466_413# _1017_/a_561_413# 0.00772f
C12367 _1017_/a_634_159# _1017_/a_975_413# 0
C12368 net141 acc0.A\[8\] 0
C12369 _0487_ _1062_/a_381_47# 0
C12370 net211 _0195_ 0
C12371 pp[28] net56 0.00857f
C12372 hold13/a_285_47# _0555_/a_51_297# 0.00175f
C12373 _0465_ _0350_ 0.07214f
C12374 _0343_ _0752_/a_300_297# 0
C12375 _0723_/a_27_413# hold80/a_285_47# 0.00182f
C12376 _0753_/a_297_297# _0375_ 0.04488f
C12377 _1052_/a_1059_315# net9 0.04781f
C12378 VPWR clkbuf_1_1__f__0457_/a_110_47# 1.2786f
C12379 output58/a_27_47# _0253_ 0.00389f
C12380 hold24/a_49_47# _0137_ 0.00179f
C12381 net103 _1060_/a_891_413# 0
C12382 _0984_/a_891_413# _0219_ 0.01037f
C12383 _0217_ net157 0.05311f
C12384 _0179_ net175 0.22618f
C12385 net190 hold50/a_285_47# 0
C12386 _0507_/a_109_47# acc0.A\[13\] 0
C12387 _1006_/a_891_413# net52 0.01608f
C12388 _1000_/a_381_47# net86 0
C12389 _1000_/a_634_159# net45 0.01903f
C12390 _1000_/a_891_413# _0098_ 0
C12391 acc0.A\[2\] _0350_ 0
C12392 _0464_ _1048_/a_27_47# 0
C12393 _0958_/a_303_47# _0161_ 0
C12394 _0149_ net154 0
C12395 _0621_/a_285_297# _0252_ 0.00139f
C12396 _0303_ acc0.A\[15\] 0.14882f
C12397 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0462_/a_110_47# 0.04845f
C12398 _0959_/a_472_297# _0477_ 0
C12399 _0463_ _0465_ 0
C12400 clknet_1_1__leaf__0463_ _0563_/a_240_47# 0
C12401 hold82/a_285_47# acc0.A\[13\] 0.00706f
C12402 clknet_1_1__leaf__0458_ _0085_ 0
C12403 _0704_/a_150_297# _0345_ 0
C12404 _0216_ _0601_/a_68_297# 0.00723f
C12405 _0521_/a_81_21# _0521_/a_299_297# 0.08213f
C12406 _0200_ _1046_/a_27_47# 0
C12407 _0536_/a_240_47# _1046_/a_466_413# 0
C12408 _1033_/a_27_47# _1033_/a_1059_315# 0.04875f
C12409 _1033_/a_193_47# _1033_/a_466_413# 0.08301f
C12410 net168 clknet_1_0__leaf__0465_ 0.00394f
C12411 _0662_/a_81_21# net66 0
C12412 net72 _0431_ 0
C12413 VPWR _0951_/a_109_93# 0.16143f
C12414 _0384_ _0345_ 0.03379f
C12415 VPWR input15/a_75_212# 0.19725f
C12416 _1012_/a_27_47# _1012_/a_1059_315# 0.04875f
C12417 _1012_/a_193_47# _1012_/a_466_413# 0.08301f
C12418 _0715_/a_27_47# _0991_/a_381_47# 0
C12419 _0289_ _0424_ 0
C12420 _0197_ _1049_/a_193_47# 0
C12421 _0352_ _1007_/a_1059_315# 0
C12422 _0758_/a_79_21# net93 0
C12423 _0107_ _1009_/a_27_47# 0.07555f
C12424 _0216_ _1031_/a_466_413# 0
C12425 _0195_ _1031_/a_891_413# 0
C12426 _0457_ _0131_ 0
C12427 _0363_ _1009_/a_466_413# 0
C12428 _0376_ _0374_ 0.04737f
C12429 _0399_ _0795_/a_81_21# 0.02794f
C12430 _0343_ _0249_ 0.07848f
C12431 control0.count\[3\] _0183_ 0
C12432 hold27/a_391_47# net125 0
C12433 _0343_ hold98/a_285_47# 0.01383f
C12434 hold21/a_285_47# net11 0
C12435 _0169_ clkbuf_1_0__f_clk/a_110_47# 0.00621f
C12436 comp0.B\[13\] net194 0
C12437 _1072_/a_381_47# clknet_0_clk 0.00739f
C12438 _1050_/a_466_413# _1050_/a_592_47# 0.00553f
C12439 _1050_/a_634_159# _1050_/a_1017_47# 0
C12440 pp[6] clknet_1_1__leaf__0458_ 0.00212f
C12441 _0518_/a_109_297# _0987_/a_27_47# 0
C12442 _0264_ hold60/a_49_47# 0
C12443 _0343_ clkload3/a_268_47# 0
C12444 _0990_/a_466_413# _0181_ 0
C12445 _0432_ _0434_ 0
C12446 _1041_/a_466_413# _0546_/a_51_297# 0.00884f
C12447 _0294_ _0393_ 0.02314f
C12448 _1024_/a_1059_315# net50 0
C12449 _0459_ _0352_ 0.00203f
C12450 VPWR _0837_/a_266_297# 0.00816f
C12451 net157 _0142_ 0
C12452 _1036_/a_891_413# net28 0
C12453 _0280_ _0218_ 0
C12454 _0565_/a_149_47# _0565_/a_240_47# 0.06872f
C12455 hold24/a_49_47# comp0.B\[6\] 0
C12456 clkload3/a_110_47# acc0.A\[17\] 0
C12457 hold24/a_285_47# comp0.B\[5\] 0
C12458 _0180_ _0527_/a_109_47# 0.00332f
C12459 net85 _1012_/a_27_47# 0
C12460 control0.state\[0\] _0965_/a_47_47# 0
C12461 _0461_ _0244_ 0.05901f
C12462 hold16/a_285_47# _0704_/a_68_297# 0
C12463 _0218_ _0246_ 0
C12464 net120 _0564_/a_68_297# 0
C12465 pp[27] hold16/a_285_47# 0
C12466 _0302_ _0277_ 0.01617f
C12467 net224 _1009_/a_1017_47# 0
C12468 _0409_ _0794_/a_326_47# 0.00409f
C12469 _0802_/a_59_75# _0403_ 0.01303f
C12470 net59 _0395_ 0
C12471 _0176_ _1040_/a_891_413# 0.03495f
C12472 _1014_/a_634_159# hold2/a_285_47# 0
C12473 acc0.A\[7\] _0180_ 0
C12474 _1039_/a_381_47# _0463_ 0.01206f
C12475 net64 net141 0
C12476 _0179_ _1054_/a_634_159# 0.04088f
C12477 clknet_1_1__leaf__0457_ _0526_/a_27_47# 0
C12478 net21 _1044_/a_634_159# 0.01703f
C12479 net183 _1044_/a_466_413# 0
C12480 _0201_ _1044_/a_891_413# 0
C12481 net179 _0621_/a_35_297# 0
C12482 acc0.A\[27\] _0323_ 0
C12483 _0788_/a_150_297# VPWR 0.00147f
C12484 control0.state\[2\] clknet_1_1__leaf_clk 0
C12485 _0833_/a_510_47# net62 0
C12486 _0995_/a_634_159# _0797_/a_27_413# 0.00698f
C12487 _0995_/a_193_47# _0797_/a_207_413# 0
C12488 net120 clknet_1_1__leaf_clk 0
C12489 _1056_/a_466_413# _0181_ 0
C12490 net21 net184 0
C12491 net231 _0175_ 0
C12492 _0750_/a_27_47# _0373_ 0.25566f
C12493 net205 _1036_/a_466_413# 0
C12494 _0973_/a_109_47# net240 0.00155f
C12495 net9 clknet_1_1__leaf__0457_ 0
C12496 _0555_/a_512_297# _0208_ 0.00161f
C12497 _0236_ _0460_ 0.07269f
C12498 _1024_/a_193_47# _1023_/a_193_47# 0.00148f
C12499 comp0.B\[13\] _1046_/a_634_159# 0
C12500 net193 _1046_/a_27_47# 0
C12501 hold98/a_49_47# net60 0
C12502 _0592_/a_68_297# net177 0
C12503 _0781_/a_150_297# _0345_ 0
C12504 net8 _1061_/a_193_47# 0
C12505 _1012_/a_193_47# net98 0.00453f
C12506 _1012_/a_466_413# clknet_1_1__leaf__0461_ 0
C12507 _1046_/a_27_47# _1046_/a_466_413# 0.26005f
C12508 _1046_/a_193_47# _1046_/a_634_159# 0.12095f
C12509 _0978_/a_27_297# _0466_ 0.22348f
C12510 _0978_/a_109_297# _0488_ 0.00225f
C12511 _0999_/a_592_47# net85 0
C12512 _0481_ _0970_/a_27_297# 0
C12513 _0316_ clknet_0__0462_ 0.03263f
C12514 hold55/a_285_47# _0208_ 0.00535f
C12515 _0270_ _0218_ 0.4793f
C12516 _0219_ _0103_ 0.00311f
C12517 net61 _0642_/a_298_297# 0
C12518 _1056_/a_193_47# _0517_/a_81_21# 0
C12519 _1056_/a_27_47# _0517_/a_299_297# 0.04767f
C12520 _0114_ clknet_1_1__leaf__0461_ 0
C12521 _1032_/a_193_47# clknet_1_0__leaf__0457_ 0.00388f
C12522 _1016_/a_381_47# net221 0.01647f
C12523 _1016_/a_193_47# _0115_ 0.02064f
C12524 net204 _0472_ 0
C12525 _0968_/a_109_297# VPWR 0
C12526 _0752_/a_300_297# _0376_ 0.12664f
C12527 net215 _1024_/a_466_413# 0
C12528 clknet_1_0__leaf__0462_ net93 0.00331f
C12529 net45 _0677_/a_47_47# 0
C12530 pp[28] _0345_ 0.00521f
C12531 _0329_ _0360_ 0
C12532 _0322_ _0321_ 0.14958f
C12533 hold18/a_285_47# _0219_ 0
C12534 _0131_ _0475_ 0.43345f
C12535 _0278_ A[13] 0
C12536 _0207_ _0205_ 0
C12537 _0664_/a_382_297# _0422_ 0
C12538 _0179_ _0281_ 0
C12539 _0322_ clkbuf_0__0460_/a_110_47# 0
C12540 _1050_/a_27_47# _1045_/a_27_47# 0.00142f
C12541 _0775_/a_297_297# _0393_ 0.00787f
C12542 clknet_0__0462_ _0347_ 0
C12543 clkbuf_1_0__f__0462_/a_110_47# _0352_ 0
C12544 VPWR _0692_/a_113_47# 0
C12545 _0984_/a_27_47# _0346_ 0.04177f
C12546 acc0.A\[20\] _0381_ 0
C12547 _0327_ _0321_ 0
C12548 _0996_/a_634_159# acc0.A\[15\] 0.00426f
C12549 clkbuf_1_1__f__0463_/a_110_47# _0215_ 0.0071f
C12550 clknet_1_0__leaf__0463_ _1038_/a_27_47# 0.05772f
C12551 _0211_ _1036_/a_634_159# 0
C12552 _0531_/a_27_297# _1049_/a_27_47# 0
C12553 _0327_ clkbuf_0__0460_/a_110_47# 0.0016f
C12554 _0839_/a_109_297# _0465_ 0
C12555 hold38/a_285_47# _0175_ 0.05331f
C12556 acc0.A\[12\] _1057_/a_634_159# 0
C12557 VPWR _0701_/a_80_21# 0.17362f
C12558 output58/a_27_47# output61/a_27_47# 0.0033f
C12559 hold27/a_391_47# _0473_ 0.01397f
C12560 _0723_/a_27_413# _0220_ 0.00147f
C12561 _0463_ net174 0
C12562 clknet_1_0__leaf__0461_ _0774_/a_68_297# 0
C12563 _0479_ control0.state\[2\] 0.00647f
C12564 _1016_/a_975_413# _0459_ 0
C12565 clknet_1_0__leaf__0465_ clknet_1_0__leaf__0464_ 0.01772f
C12566 _0857_/a_27_47# _1032_/a_1059_315# 0
C12567 _0279_ _0278_ 0.18238f
C12568 _0539_/a_150_297# _0176_ 0
C12569 _0175_ clknet_1_1__leaf__0457_ 0
C12570 net44 _0999_/a_634_159# 0
C12571 _0246_ _0775_/a_215_47# 0
C12572 clknet_0__0463_ control0.sh 0.04084f
C12573 control0.count\[2\] _0169_ 0.20463f
C12574 net185 net119 0
C12575 net103 _0218_ 0
C12576 hold34/a_285_47# VPWR 0.2591f
C12577 hold23/a_391_47# clknet_1_0__leaf__0464_ 0.00169f
C12578 _0181_ _0584_/a_27_297# 0.14741f
C12579 _1000_/a_193_47# net46 0
C12580 net57 _0219_ 0.02957f
C12581 _1052_/a_634_159# _0522_/a_109_297# 0
C12582 _1052_/a_466_413# _0522_/a_27_297# 0.0017f
C12583 hold26/a_391_47# net7 0
C12584 _0482_ clk 0.00641f
C12585 clknet_0__0459_ _0645_/a_47_47# 0.03163f
C12586 _0721_/a_27_47# clknet_1_0__leaf__0457_ 0.01931f
C12587 _0093_ net81 0.14018f
C12588 _0598_/a_79_21# _0227_ 0.15215f
C12589 _0467_ _0166_ 0
C12590 _0518_/a_109_297# _0191_ 0.00344f
C12591 _0518_/a_373_47# net15 0.00181f
C12592 VPWR _0675_/a_68_297# 0.14621f
C12593 hold41/a_391_47# VPWR 0.1713f
C12594 _1039_/a_193_47# net8 0.0651f
C12595 _0985_/a_193_47# _0083_ 0.41008f
C12596 _0985_/a_891_413# _0985_/a_1017_47# 0.00617f
C12597 _0214_ _0562_/a_68_297# 0.10606f
C12598 _0183_ net176 0
C12599 hold10/a_285_47# _0501_/a_27_47# 0.02027f
C12600 net233 _0218_ 0
C12601 _1018_/a_891_413# _1018_/a_975_413# 0.00851f
C12602 _1018_/a_27_47# net104 0.22945f
C12603 _1018_/a_381_47# _1018_/a_561_413# 0.00123f
C12604 net178 net182 0
C12605 _0277_ net6 0.07149f
C12606 comp0.B\[7\] hold26/a_49_47# 0
C12607 _0275_ clknet_1_1__leaf__0465_ 0
C12608 clknet_1_1__leaf__0461_ net98 0.15767f
C12609 _0298_ _0795_/a_299_297# 0
C12610 _0404_ _0795_/a_384_47# 0
C12611 hold47/a_285_47# acc0.A\[4\] 0
C12612 _0716_/a_27_47# hold81/a_285_47# 0
C12613 _0982_/a_634_159# _0982_/a_975_413# 0
C12614 _0982_/a_466_413# _0982_/a_561_413# 0.00772f
C12615 net96 acc0.A\[29\] 0
C12616 _0353_ _0339_ 0.04691f
C12617 _1049_/a_1059_315# _1049_/a_891_413# 0.31086f
C12618 _1049_/a_193_47# _1049_/a_975_413# 0
C12619 _1049_/a_466_413# _1049_/a_381_47# 0.03733f
C12620 _0983_/a_592_47# acc0.A\[15\] 0
C12621 net82 net41 0
C12622 _0194_ _0522_/a_27_297# 0.00185f
C12623 _0524_/a_27_297# _0193_ 0
C12624 net12 _0522_/a_109_47# 0
C12625 net207 _0459_ 0
C12626 _0343_ _0231_ 0.39813f
C12627 clkbuf_0__0465_/a_110_47# _0186_ 0
C12628 _0747_/a_79_21# _0747_/a_297_297# 0.01735f
C12629 net39 _0297_ 0
C12630 _0666_/a_113_47# _0277_ 0
C12631 _0383_ _0345_ 0
C12632 _0552_/a_68_297# _0209_ 0.10716f
C12633 VPWR _0618_/a_79_21# 0.44395f
C12634 clkload3/Y clknet_1_1__leaf__0461_ 0.34003f
C12635 _1053_/a_27_47# _1053_/a_634_159# 0.14145f
C12636 _0575_/a_27_297# _0575_/a_109_297# 0.17136f
C12637 _0220_ _0352_ 0
C12638 _0760_/a_377_297# _0460_ 0
C12639 _0637_/a_56_297# _0267_ 0.04595f
C12640 _1019_/a_1059_315# _0218_ 0
C12641 net158 _0172_ 0.08653f
C12642 _0195_ _1008_/a_193_47# 0
C12643 hold39/a_285_47# _1065_/a_27_47# 0
C12644 hold16/a_285_47# _0216_ 0
C12645 _1066_/a_1059_315# _1066_/a_891_413# 0.31086f
C12646 _1066_/a_193_47# _1066_/a_975_413# 0
C12647 _1066_/a_466_413# _1066_/a_381_47# 0.03733f
C12648 _0269_ net72 0.0448f
C12649 _0831_/a_35_297# acc0.A\[8\] 0.00424f
C12650 output37/a_27_47# net3 0.03711f
C12651 clkbuf_1_1__f__0461_/a_110_47# _0397_ 0.00787f
C12652 net1 _1066_/a_466_413# 0
C12653 net45 _0242_ 0.03574f
C12654 net45 _0999_/a_592_47# 0
C12655 VPWR _1052_/a_1017_47# 0
C12656 net31 _1040_/a_27_47# 0
C12657 _0833_/a_215_47# net235 0.07174f
C12658 _0201_ _1042_/a_27_47# 0
C12659 _1023_/a_381_47# _1022_/a_1059_315# 0
C12660 _0680_/a_80_21# _0462_ 0.02207f
C12661 _0476_ clk 0.0068f
C12662 _0401_ _0809_/a_299_297# 0.05078f
C12663 _1068_/a_1059_315# _1068_/a_891_413# 0.31086f
C12664 _1068_/a_193_47# _1068_/a_975_413# 0
C12665 _1068_/a_466_413# _1068_/a_381_47# 0.03733f
C12666 _0343_ clkbuf_1_1__f__0461_/a_110_47# 0.00518f
C12667 _1030_/a_27_47# _1030_/a_1059_315# 0.04875f
C12668 _1030_/a_193_47# _1030_/a_466_413# 0.07855f
C12669 _1041_/a_27_47# _0176_ 0
C12670 _0257_ net170 0
C12671 acc0.A\[14\] _0451_ 0.06095f
C12672 acc0.A\[22\] hold68/a_285_47# 0
C12673 _0183_ hold68/a_49_47# 0
C12674 _0217_ hold68/a_391_47# 0.06181f
C12675 _0402_ _0807_/a_150_297# 0
C12676 _1017_/a_193_47# _0347_ 0
C12677 _0322_ _1009_/a_27_47# 0
C12678 _0343_ _0426_ 0
C12679 net205 comp0.B\[6\] 0
C12680 _0476_ _0959_/a_217_297# 0.00489f
C12681 _0217_ _0462_ 0.02603f
C12682 _0330_ _0726_/a_51_297# 0
C12683 _0251_ _0519_/a_299_297# 0
C12684 hold9/a_49_47# hold9/a_285_47# 0.22264f
C12685 _0416_ _0278_ 0
C12686 _1056_/a_592_47# acc0.A\[9\] 0
C12687 net148 _0523_/a_299_297# 0.05915f
C12688 _1035_/a_1059_315# clknet_1_1__leaf__0463_ 0.00882f
C12689 _1035_/a_634_159# net122 0
C12690 _0753_/a_79_21# net46 0
C12691 _0992_/a_27_47# net37 0
C12692 _0992_/a_891_413# hold70/a_49_47# 0.00267f
C12693 _0992_/a_466_413# hold70/a_391_47# 0
C12694 clknet_0__0465_ net47 0.1549f
C12695 VPWR _0486_ 1.59078f
C12696 hold53/a_285_47# net200 0.01228f
C12697 _0251_ output65/a_27_47# 0
C12698 _0598_/a_382_297# _0598_/a_297_47# 0
C12699 clkbuf_1_0__f__0459_/a_110_47# _0507_/a_27_297# 0.00384f
C12700 _1015_/a_634_159# _0181_ 0.00939f
C12701 _0987_/a_27_47# _0987_/a_193_47# 0.96607f
C12702 _0238_ _0748_/a_299_297# 0
C12703 _1034_/a_381_47# comp0.B\[2\] 0.01618f
C12704 pp[7] acc0.A\[7\] 0
C12705 control0.state\[1\] _0175_ 0.00256f
C12706 pp[7] _0989_/a_1059_315# 0
C12707 _0343_ _0185_ 0.00113f
C12708 net123 VPWR 0.43262f
C12709 _0125_ _1008_/a_634_159# 0
C12710 acc0.A\[27\] _1008_/a_891_413# 0.00551f
C12711 _0992_/a_634_159# net67 0.00112f
C12712 _0341_ clknet_1_1__leaf__0462_ 0.01116f
C12713 _1000_/a_634_159# VPWR 0.18153f
C12714 VPWR input32/a_75_212# 0.26736f
C12715 _0093_ _0797_/a_207_413# 0.0099f
C12716 _0480_ _0488_ 0.3817f
C12717 _0983_/a_891_413# _0181_ 0.00543f
C12718 _0796_/a_297_297# net41 0
C12719 _1072_/a_1059_315# _0466_ 0
C12720 _0211_ comp0.B\[5\] 0.0307f
C12721 _0657_/a_109_297# clknet_1_1__leaf__0465_ 0.00198f
C12722 _0465_ _0847_/a_109_297# 0
C12723 _0149_ clknet_0__0464_ 0
C12724 hold89/a_285_47# clk 0.05035f
C12725 _0298_ net6 0.39168f
C12726 _1000_/a_27_47# clkbuf_0__0461_/a_110_47# 0
C12727 hold23/a_391_47# hold28/a_49_47# 0.00144f
C12728 hold35/a_49_47# acc0.A\[10\] 0.00247f
C12729 _1029_/a_27_47# _1029_/a_193_47# 0.97453f
C12730 _0254_ _0350_ 0
C12731 hold2/a_285_47# net247 0
C12732 _0370_ _0460_ 0.02697f
C12733 hold52/a_391_47# _0216_ 0
C12734 output65/a_27_47# net58 0
C12735 _0352_ _0772_/a_79_21# 0.15752f
C12736 _0296_ net6 0
C12737 _0679_/a_68_297# net52 0
C12738 _0095_ net42 0.2684f
C12739 _0179_ A[12] 0
C12740 pp[30] _1031_/a_1017_47# 0
C12741 _1032_/a_381_47# clknet_1_0__leaf__0461_ 0.00973f
C12742 _0666_/a_113_47# _0298_ 0.00963f
C12743 net144 A[11] 0.03177f
C12744 hold57/a_285_47# net36 0
C12745 net175 _0530_/a_384_47# 0.01033f
C12746 net61 _0639_/a_109_297# 0.00324f
C12747 _0343_ _0998_/a_1059_315# 0.00407f
C12748 _0722_/a_79_21# clknet_1_1__leaf__0462_ 0.0017f
C12749 _1008_/a_891_413# _0364_ 0.00394f
C12750 net64 _0831_/a_35_297# 0.00106f
C12751 comp0.B\[13\] _1045_/a_27_47# 0.0017f
C12752 _0399_ _0580_/a_27_297# 0.03056f
C12753 _0172_ net148 0
C12754 _0645_/a_285_47# _0996_/a_193_47# 0
C12755 clknet_1_0__leaf__0465_ _0536_/a_245_297# 0
C12756 _1017_/a_193_47# _1016_/a_891_413# 0
C12757 _1017_/a_466_413# _1016_/a_466_413# 0.00104f
C12758 hold55/a_391_47# _0178_ 0
C12759 _0520_/a_109_297# _0180_ 0.01052f
C12760 _0231_ _0376_ 0
C12761 acc0.A\[8\] _0988_/a_381_47# 0
C12762 _0254_ _0621_/a_35_297# 0
C12763 _0402_ _0422_ 0.19324f
C12764 _0998_/a_466_413# acc0.A\[17\] 0
C12765 _0324_ _0687_/a_59_75# 0
C12766 acc0.A\[21\] net49 0.58585f
C12767 _0578_/a_109_47# acc0.A\[20\] 0
C12768 _0643_/a_253_297# _0255_ 0
C12769 _1016_/a_27_47# _0158_ 0
C12770 net166 _1060_/a_27_47# 0
C12771 net229 _0345_ 0
C12772 _1037_/a_193_47# clknet_1_1__leaf__0463_ 0
C12773 _0756_/a_47_47# _1023_/a_634_159# 0
C12774 net21 _0176_ 0.06104f
C12775 net86 net45 0.00662f
C12776 _0998_/a_193_47# clkbuf_1_1__f__0461_/a_110_47# 0.01155f
C12777 _0555_/a_51_297# _0555_/a_149_47# 0.02487f
C12778 clknet_1_0__leaf__0459_ _0675_/a_68_297# 0
C12779 _0363_ net96 0
C12780 A[12] _0513_/a_81_21# 0
C12781 _0427_ acc0.A\[9\] 0.04047f
C12782 hold41/a_49_47# _1057_/a_27_47# 0
C12783 net2 _0186_ 0.14413f
C12784 _0415_ _0092_ 0
C12785 _0113_ clkbuf_1_1__f__0457_/a_110_47# 0
C12786 hold38/a_49_47# clknet_0_clk 0
C12787 _1067_/a_193_47# _1065_/a_1059_315# 0
C12788 _1067_/a_27_47# _1065_/a_891_413# 0
C12789 _0399_ _0790_/a_117_297# 0
C12790 _0846_/a_51_297# _0843_/a_68_297# 0
C12791 net58 _0986_/a_193_47# 0.03305f
C12792 _0299_ _0797_/a_297_47# 0.00223f
C12793 hold47/a_391_47# clknet_1_0__leaf__0465_ 0.0056f
C12794 _0308_ _1009_/a_193_47# 0
C12795 _1033_/a_891_413# _1033_/a_1017_47# 0.00617f
C12796 _1033_/a_193_47# _0131_ 0.2529f
C12797 hold87/a_391_47# _0263_ 0
C12798 _0985_/a_27_47# VPWR 0.65025f
C12799 net63 _0987_/a_634_159# 0
C12800 _0352_ net51 0.15641f
C12801 _0965_/a_47_47# _0478_ 0.40179f
C12802 _0841_/a_297_297# _0345_ 0.00557f
C12803 _1012_/a_891_413# _1012_/a_1017_47# 0.00617f
C12804 _0130_ _1033_/a_466_413# 0
C12805 _0856_/a_79_21# hold60/a_49_47# 0
C12806 net118 clknet_1_1__leaf_clk 0
C12807 _0846_/a_512_297# _0219_ 0
C12808 net226 _0485_ 0
C12809 _0244_ _0582_/a_27_297# 0
C12810 _0102_ _0105_ 0
C12811 hold55/a_49_47# hold55/a_285_47# 0.22264f
C12812 net76 _0988_/a_975_413# 0
C12813 _0753_/a_297_297# VPWR 0.29324f
C12814 _1054_/a_27_47# hold83/a_391_47# 0
C12815 _0248_ _0462_ 0.08144f
C12816 clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0457_ 0
C12817 _1009_/a_891_413# _0219_ 0.05913f
C12818 hold86/a_391_47# net233 0.14294f
C12819 _1050_/a_381_47# acc0.A\[4\] 0.01617f
C12820 _0459_ hold72/a_285_47# 0.01808f
C12821 net15 _0987_/a_466_413# 0
C12822 clkbuf_1_0__f__0463_/a_110_47# _0465_ 0
C12823 hold54/a_49_47# _0457_ 0.00235f
C12824 _1055_/a_561_413# acc0.A\[9\] 0
C12825 _0088_ _0181_ 0.02436f
C12826 hold26/a_391_47# _0202_ 0
C12827 _1041_/a_891_413# net152 0.00226f
C12828 _1041_/a_1059_315# net32 0
C12829 hold100/a_391_47# _0458_ 0
C12830 VPWR _0677_/a_47_47# 0.38209f
C12831 _0718_/a_47_47# _0353_ 0
C12832 _0967_/a_109_93# _0946_/a_30_53# 0
C12833 net62 _0347_ 0
C12834 _0946_/a_30_53# _0487_ 0.00866f
C12835 _0163_ _0215_ 0.0013f
C12836 _0346_ clkbuf_0__0460_/a_110_47# 0
C12837 net36 _0159_ 0
C12838 _0450_ _0347_ 0
C12839 _0517_/a_81_21# clknet_1_1__leaf__0465_ 0.00279f
C12840 _0508_/a_81_21# net228 0.05912f
C12841 comp0.B\[4\] B[5] 0
C12842 _0229_ _0606_/a_215_297# 0
C12843 VPWR _0544_/a_149_47# 0
C12844 _0993_/a_193_47# net79 0.00438f
C12845 _0983_/a_466_413# _1018_/a_634_159# 0
C12846 hold87/a_285_47# _0459_ 0
C12847 comp0.B\[14\] _1045_/a_891_413# 0
C12848 net34 _0483_ 0
C12849 VPWR _1034_/a_1059_315# 0.3816f
C12850 clknet_1_0__leaf__0460_ _1067_/a_634_159# 0
C12851 _0179_ _1057_/a_193_47# 0
C12852 net198 _1043_/a_193_47# 0.02976f
C12853 net18 _1043_/a_27_47# 0.0287f
C12854 _0960_/a_27_47# control0.count\[1\] 0.16031f
C12855 _0343_ _0983_/a_27_47# 0.00782f
C12856 _0531_/a_27_297# _0531_/a_109_47# 0.00393f
C12857 _0996_/a_27_47# _0507_/a_109_297# 0
C12858 clknet_0__0458_ _0345_ 0.3103f
C12859 net68 _0112_ 0
C12860 _0553_/a_149_47# _0463_ 0
C12861 hold6/a_391_47# _1043_/a_466_413# 0
C12862 _1053_/a_891_413# input12/a_75_212# 0
C12863 _1053_/a_634_159# A[5] 0.00131f
C12864 _0179_ net140 0.00109f
C12865 net87 hold40/a_391_47# 0
C12866 net46 _0250_ 0
C12867 net21 net130 0.01377f
C12868 _1002_/a_193_47# acc0.A\[20\] 0
C12869 _0998_/a_634_159# _0998_/a_466_413# 0.23992f
C12870 _0998_/a_193_47# _0998_/a_1059_315# 0.03405f
C12871 _0998_/a_27_47# _0998_/a_891_413# 0.03089f
C12872 hold32/a_391_47# VPWR 0.22198f
C12873 pp[17] _0708_/a_68_297# 0.01135f
C12874 output44/a_27_47# net60 0
C12875 net57 hold61/a_49_47# 0
C12876 _0956_/a_304_297# _0208_ 0.00166f
C12877 comp0.B\[15\] _0173_ 0.00398f
C12878 net58 _0845_/a_109_47# 0
C12879 clknet_1_1__leaf__0459_ net60 0.00168f
C12880 _0349_ net208 0
C12881 _1055_/a_634_159# _0369_ 0
C12882 net64 _0988_/a_381_47# 0.01613f
C12883 net45 _1018_/a_1017_47# 0
C12884 _1059_/a_466_413# _0459_ 0.00289f
C12885 hold64/a_391_47# _0345_ 0.01353f
C12886 _1031_/a_1017_47# _0339_ 0
C12887 _1003_/a_193_47# _0369_ 0
C12888 _0796_/a_215_47# _0400_ 0
C12889 clknet_1_1__leaf__0459_ net5 0.02634f
C12890 _0498_/a_51_297# _1061_/a_634_159# 0.00128f
C12891 net110 _1023_/a_27_47# 0
C12892 hold56/a_49_47# _1033_/a_27_47# 0
C12893 _0662_/a_299_297# _0986_/a_193_47# 0
C12894 comp0.B\[13\] net132 0
C12895 _0769_/a_384_47# clknet_1_0__leaf__0461_ 0
C12896 clknet_0__0463_ _0955_/a_32_297# 0
C12897 _0280_ net228 0
C12898 hold87/a_391_47# clknet_1_0__leaf__0461_ 0.00192f
C12899 hold38/a_391_47# _0955_/a_32_297# 0.01532f
C12900 VPWR _0507_/a_109_47# 0
C12901 _1019_/a_27_47# _1019_/a_466_413# 0.26005f
C12902 _1019_/a_193_47# _1019_/a_634_159# 0.12729f
C12903 net44 _1012_/a_1059_315# 0.0106f
C12904 _1046_/a_193_47# net132 0.00374f
C12905 _1046_/a_1059_315# _1046_/a_1017_47# 0
C12906 _1000_/a_634_159# clknet_1_0__leaf__0459_ 0
C12907 _0218_ _0774_/a_68_297# 0.16674f
C12908 _0557_/a_51_297# net171 0
C12909 _0949_/a_59_75# clkbuf_0_clk/a_110_47# 0.01323f
C12910 _1056_/a_1059_315# _0153_ 0
C12911 _0809_/a_81_21# hold70/a_285_47# 0
C12912 clkbuf_0__0464_/a_110_47# net10 0
C12913 clknet_1_0__leaf__0463_ B[6] 0.00998f
C12914 _0837_/a_81_21# _0172_ 0.17319f
C12915 net133 _0533_/a_109_297# 0
C12916 net61 output58/a_27_47# 0.02272f
C12917 VPWR _1012_/a_27_47# 0.71251f
C12918 net34 control0.count\[1\] 0
C12919 VPWR hold82/a_285_47# 0.27904f
C12920 _0221_ _0335_ 0.70506f
C12921 VPWR _0330_ 0.51042f
C12922 _0218_ _0085_ 0
C12923 _0343_ _0225_ 0.047f
C12924 net215 _0122_ 0.21391f
C12925 _0684_/a_59_75# net55 0.16258f
C12926 _0565_/a_245_297# _0175_ 0
C12927 _0548_/a_51_297# _1040_/a_1059_315# 0
C12928 _0473_ _0496_/a_27_47# 0.02655f
C12929 net205 net26 0.10058f
C12930 _0982_/a_891_413# clkbuf_0__0457_/a_110_47# 0
C12931 acc0.A\[9\] net142 0.22116f
C12932 net196 net195 0.00136f
C12933 net9 _1049_/a_634_159# 0.00325f
C12934 net175 _1049_/a_891_413# 0.00109f
C12935 _0343_ _0436_ 0.24272f
C12936 _0183_ acc0.A\[18\] 0.09467f
C12937 output55/a_27_47# net242 0
C12938 pp[27] _0729_/a_68_297# 0
C12939 _0557_/a_51_297# net24 0
C12940 _0210_ comp0.B\[5\] 0.07893f
C12941 net160 comp0.B\[6\] 0.14509f
C12942 _0775_/a_510_47# _0352_ 0.00633f
C12943 acc0.A\[31\] _1031_/a_27_47# 0
C12944 hold15/a_285_47# _1031_/a_1059_315# 0.0129f
C12945 _0457_ _1032_/a_1017_47# 0
C12946 net105 _0208_ 0.00591f
C12947 net44 net85 0
C12948 _0336_ net209 0
C12949 hold76/a_285_47# _0247_ 0
C12950 control0.state\[0\] clknet_0_clk 0.09516f
C12951 _1021_/a_27_47# _0578_/a_27_297# 0
C12952 hold88/a_49_47# hold88/a_391_47# 0.00188f
C12953 _0179_ _0154_ 0.00787f
C12954 VPWR _0242_ 0.75426f
C12955 _1024_/a_27_47# pp[24] 0.00123f
C12956 _1024_/a_634_159# net52 0.00723f
C12957 _1024_/a_891_413# output52/a_27_47# 0.00113f
C12958 clkload3/a_110_47# net84 0
C12959 VPWR _0999_/a_592_47# 0
C12960 _0459_ _0392_ 0
C12961 _1052_/a_975_413# acc0.A\[6\] 0
C12962 _1052_/a_466_413# _0193_ 0
C12963 _0581_/a_109_297# net206 0.02099f
C12964 _0990_/a_27_47# _0990_/a_1059_315# 0.04875f
C12965 _0990_/a_193_47# _0990_/a_466_413# 0.07855f
C12966 _0347_ _0687_/a_59_75# 0
C12967 _0732_/a_209_297# VPWR 0.20952f
C12968 clknet_0__0458_ clkload1/a_268_47# 0
C12969 comp0.B\[2\] net201 0.00571f
C12970 _0267_ _0849_/a_79_21# 0.00711f
C12971 _0313_ hold90/a_49_47# 0
C12972 net168 _0519_/a_299_297# 0.05857f
C12973 net125 _0180_ 0
C12974 hold7/a_285_47# _0525_/a_299_297# 0
C12975 _0984_/a_891_413# net58 0.00498f
C12976 hold27/a_391_47# comp0.B\[8\] 0.01857f
C12977 _0264_ _0263_ 0.0065f
C12978 clkbuf_1_0__f__0463_/a_110_47# net174 0
C12979 _0172_ _0542_/a_240_47# 0.02331f
C12980 _0174_ _0546_/a_51_297# 0.12574f
C12981 clkbuf_0__0465_/a_110_47# net62 0.00946f
C12982 net36 acc0.A\[0\] 0.01998f
C12983 net203 _0173_ 0.47812f
C12984 hold19/a_391_47# net166 0.13432f
C12985 hold56/a_391_47# _0132_ 0
C12986 _0343_ _0990_/a_592_47# 0
C12987 _0985_/a_381_47# acc0.A\[3\] 0.00706f
C12988 _0433_ _0828_/a_113_297# 0
C12989 acc0.A\[25\] _1007_/a_193_47# 0
C12990 _0967_/a_109_93# _0487_ 0
C12991 _0967_/a_215_297# _0485_ 0.38301f
C12992 _0346_ _1014_/a_891_413# 0.01064f
C12993 _0484_ _0162_ 0.32771f
C12994 _0343_ _0793_/a_149_47# 0.00131f
C12995 net75 acc0.A\[6\] 0
C12996 _0343_ clknet_0__0459_ 0.01187f
C12997 clknet_1_1__leaf__0463_ _1062_/a_193_47# 0
C12998 hold88/a_285_47# _0086_ 0
C12999 _1049_/a_381_47# _0147_ 0.12885f
C13000 _1049_/a_466_413# acc0.A\[3\] 0
C13001 _0552_/a_150_297# _0175_ 0
C13002 clknet_1_1__leaf__0459_ acc0.A\[11\] 0.01154f
C13003 clknet_0__0465_ _0294_ 0
C13004 hold9/a_285_47# _0739_/a_79_21# 0.00244f
C13005 _0194_ _0193_ 0
C13006 _0818_/a_193_47# acc0.A\[9\] 0
C13007 hold9/a_391_47# _0347_ 0.00172f
C13008 _0461_ _0195_ 0.00307f
C13009 _0229_ hold3/a_49_47# 0
C13010 _0747_/a_215_47# _0104_ 0
C13011 net248 _0989_/a_634_159# 0
C13012 _0598_/a_79_21# _0352_ 0.00387f
C13013 VPWR _0197_ 0.72598f
C13014 _1070_/a_1059_315# _1070_/a_891_413# 0.31086f
C13015 _1070_/a_193_47# _1070_/a_975_413# 0
C13016 _1070_/a_466_413# _1070_/a_381_47# 0.03733f
C13017 _1052_/a_634_159# _0150_ 0.03783f
C13018 _0137_ acc0.A\[15\] 0
C13019 _1053_/a_891_413# _1053_/a_975_413# 0.00851f
C13020 _1053_/a_27_47# net139 0.22665f
C13021 _1053_/a_381_47# _1053_/a_561_413# 0.00123f
C13022 pp[17] _1030_/a_634_159# 0
C13023 net44 _1030_/a_1059_315# 0.09497f
C13024 _1057_/a_561_413# acc0.A\[10\] 0
C13025 _1015_/a_1059_315# net118 0
C13026 clknet_1_0__leaf__0465_ _1050_/a_561_413# 0
C13027 _0960_/a_109_47# control0.count\[2\] 0
C13028 net45 _0998_/a_381_47# 0.00204f
C13029 acc0.A\[22\] _1023_/a_1059_315# 0.00353f
C13030 _0217_ _1023_/a_891_413# 0
C13031 _0816_/a_150_297# clknet_1_1__leaf__0465_ 0
C13032 _0198_ _1061_/a_1059_315# 0
C13033 _1032_/a_1059_315# _0208_ 0
C13034 hold43/a_391_47# _0216_ 0.04017f
C13035 _1066_/a_466_413# control0.sh 0.00278f
C13036 _1014_/a_27_47# _0465_ 0
C13037 hold37/a_49_47# acc0.A\[4\] 0.07788f
C13038 _1062_/a_27_47# _0468_ 0.00164f
C13039 hold33/a_285_47# net36 0
C13040 _0217_ hold59/a_391_47# 0.06121f
C13041 _0183_ hold59/a_49_47# 0
C13042 VPWR _1030_/a_27_47# 0.60874f
C13043 _0995_/a_27_47# net43 0
C13044 clknet_1_1__leaf__0463_ _0561_/a_245_297# 0
C13045 _0756_/a_47_47# _0377_ 0
C13046 _0559_/a_51_297# _1034_/a_891_413# 0
C13047 _0263_ net170 0
C13048 net7 _1040_/a_27_47# 0
C13049 _0935_/a_27_47# _0492_/a_27_47# 0
C13050 input10/a_75_212# input18/a_75_212# 0.01223f
C13051 _1061_/a_193_47# _0492_/a_27_47# 0
C13052 net1 _0166_ 0
C13053 _1068_/a_381_47# _0166_ 0.11632f
C13054 _0749_/a_81_21# _0345_ 0.01098f
C13055 _1030_/a_891_413# _1030_/a_1017_47# 0.00617f
C13056 _0414_ _0403_ 0.35287f
C13057 VPWR A[6] 0.34719f
C13058 _0328_ acc0.A\[25\] 0.05608f
C13059 _0997_/a_634_159# net83 0
C13060 _1038_/a_891_413# _0552_/a_68_297# 0.00141f
C13061 hold63/a_391_47# hold53/a_285_47# 0
C13062 hold63/a_285_47# hold53/a_391_47# 0
C13063 clknet_1_0__leaf__0458_ _0261_ 0.02449f
C13064 _0274_ _0399_ 0.02434f
C13065 _0376_ _0225_ 0.20414f
C13066 hold27/a_391_47# _1046_/a_466_413# 0
C13067 net123 _1036_/a_27_47# 0
C13068 net138 acc0.A\[6\] 0
C13069 _0592_/a_68_297# hold4/a_49_47# 0
C13070 VPWR net190 0.27847f
C13071 net121 net122 0.00486f
C13072 clknet_1_0__leaf__0465_ _0623_/a_109_297# 0
C13073 _1056_/a_27_47# _1056_/a_1059_315# 0.04875f
C13074 _1056_/a_193_47# _1056_/a_466_413# 0.07482f
C13075 _1032_/a_466_413# net17 0.00567f
C13076 _0092_ _0347_ 0
C13077 _0402_ _0423_ 0
C13078 _0390_ _0242_ 0
C13079 net61 clkbuf_1_0__f__0465_/a_110_47# 0.01765f
C13080 _0310_ _0746_/a_384_47# 0
C13081 _0458_ _0256_ 0
C13082 hold28/a_49_47# hold71/a_391_47# 0
C13083 VPWR _0153_ 0.76449f
C13084 clkbuf_1_0__f__0459_/a_110_47# _0185_ 0.00284f
C13085 _0320_ _0364_ 0.05251f
C13086 _0987_/a_634_159# _0987_/a_1017_47# 0
C13087 _0987_/a_466_413# _0987_/a_592_47# 0.00553f
C13088 _0264_ clknet_1_0__leaf__0461_ 0.00485f
C13089 _0307_ _0777_/a_47_47# 0.00249f
C13090 hold74/a_49_47# _0398_ 0
C13091 _0114_ clknet_1_1__leaf__0465_ 0
C13092 hold47/a_285_47# _0149_ 0
C13093 hold47/a_391_47# net137 0
C13094 _0924_/a_27_47# _0181_ 0
C13095 net211 _0183_ 0.05077f
C13096 net44 net45 0.01594f
C13097 _0741_/a_109_297# clknet_1_0__leaf__0460_ 0
C13098 _0312_ _0367_ 0
C13099 _0235_ _0462_ 0.00783f
C13100 clknet_1_1__leaf__0458_ _0525_/a_81_21# 0
C13101 clknet_1_1__leaf__0459_ hold81/a_391_47# 0.00837f
C13102 clkload2/a_110_47# clknet_1_0__leaf__0464_ 0
C13103 _0661_/a_27_297# VPWR 0.1317f
C13104 _0558_/a_150_297# clknet_1_1__leaf__0463_ 0
C13105 acc0.A\[1\] _1047_/a_381_47# 0
C13106 _0199_ _1047_/a_193_47# 0.0241f
C13107 net62 _0824_/a_59_75# 0
C13108 _1047_/a_1059_315# net218 0
C13109 net86 VPWR 0.46684f
C13110 _1004_/a_466_413# _1004_/a_381_47# 0.03733f
C13111 _1004_/a_193_47# _1004_/a_975_413# 0
C13112 _1004_/a_1059_315# _1004_/a_891_413# 0.31086f
C13113 _0549_/a_68_297# net28 0
C13114 clknet_0__0458_ _0836_/a_68_297# 0
C13115 _0317_ clkbuf_0__0462_/a_110_47# 0
C13116 net47 _0986_/a_27_47# 0
C13117 _1027_/a_1059_315# _1008_/a_27_47# 0
C13118 _1027_/a_193_47# _1008_/a_466_413# 0
C13119 _1027_/a_27_47# _1008_/a_1059_315# 0
C13120 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0464_/a_110_47# 0.00554f
C13121 net157 _1049_/a_466_413# 0
C13122 acc0.A\[30\] hold61/a_391_47# 0.01954f
C13123 acc0.A\[31\] _0712_/a_79_21# 0
C13124 hold23/a_391_47# clkbuf_1_0__f__0464_/a_110_47# 0.01439f
C13125 hold18/a_391_47# _0465_ 0.01458f
C13126 _1067_/a_193_47# hold93/a_49_47# 0
C13127 _1067_/a_27_47# hold93/a_285_47# 0
C13128 _0680_/a_80_21# _0312_ 0.19366f
C13129 _0369_ hold93/a_391_47# 0
C13130 clknet_1_0__leaf__0465_ _1053_/a_634_159# 0.00629f
C13131 _1029_/a_466_413# _1029_/a_592_47# 0.00553f
C13132 _1029_/a_634_159# _1029_/a_1017_47# 0
C13133 net58 hold18/a_285_47# 0
C13134 _0583_/a_109_297# net102 0
C13135 _1019_/a_27_47# _0352_ 0
C13136 _0538_/a_51_297# _0954_/a_32_297# 0.00112f
C13137 clknet_1_0__leaf__0458_ _0509_/a_27_47# 0.00198f
C13138 hold87/a_285_47# _0267_ 0
C13139 _0195_ _0997_/a_1059_315# 0
C13140 _0228_ _0378_ 0
C13141 clkbuf_1_1__f__0460_/a_110_47# _0219_ 0
C13142 pp[15] net6 0
C13143 _0328_ _0737_/a_117_297# 0.00239f
C13144 _0817_/a_368_297# _0345_ 0.00121f
C13145 _0314_ clknet_0__0462_ 0.002f
C13146 clkload0/X _1072_/a_1059_315# 0
C13147 _0346_ _0795_/a_81_21# 0.18759f
C13148 _0351_ _0778_/a_68_297# 0
C13149 _0399_ _0117_ 0.12225f
C13150 hold66/a_285_47# net241 0
C13151 hold66/a_49_47# _0219_ 0.00146f
C13152 acc0.A\[4\] _0987_/a_381_47# 0.00355f
C13153 _0387_ _0294_ 0.00589f
C13154 _0961_/a_199_47# _0479_ 0.00151f
C13155 _0195_ _0465_ 0.05342f
C13156 _1020_/a_193_47# _0217_ 0
C13157 _1020_/a_634_159# net150 0
C13158 clkbuf_1_1__f__0460_/a_110_47# _0728_/a_59_75# 0
C13159 net72 clkbuf_0__0458_/a_110_47# 0.00104f
C13160 _0324_ _0352_ 0.04224f
C13161 _0180_ _0186_ 1.29936f
C13162 _0747_/a_79_21# _0326_ 0.00138f
C13163 net219 _0347_ 0.01547f
C13164 _0399_ net43 0.06509f
C13165 output66/a_27_47# acc0.A\[9\] 0
C13166 net44 _0587_/a_27_47# 0.1822f
C13167 _0237_ net51 0.00792f
C13168 clknet_1_0__leaf__0459_ _0242_ 0.09568f
C13169 _1016_/a_27_47# _1016_/a_634_159# 0.13601f
C13170 _0856_/a_510_47# _0465_ 0
C13171 acc0.A\[2\] _0195_ 0.23715f
C13172 _0483_ _1068_/a_466_413# 0
C13173 control0.count\[3\] _1068_/a_891_413# 0
C13174 hold11/a_49_47# _1061_/a_27_47# 0
C13175 _0379_ _1023_/a_1059_315# 0
C13176 _0756_/a_47_47# net109 0
C13177 clknet_1_1__leaf__0460_ hold69/a_285_47# 0.02844f
C13178 _0101_ _0103_ 0
C13179 _1033_/a_1059_315# comp0.B\[15\] 0
C13180 _1028_/a_634_159# _1028_/a_592_47# 0
C13181 _0236_ _0373_ 0.54723f
C13182 net188 hold42/a_285_47# 0.03458f
C13183 _0407_ clknet_1_1__leaf__0461_ 0
C13184 net58 _0856_/a_215_47# 0
C13185 _0343_ _0996_/a_1059_315# 0.00272f
C13186 _0369_ _0989_/a_561_413# 0
C13187 clknet_1_0__leaf__0458_ net47 0.13496f
C13188 _0765_/a_297_297# _0460_ 0.00187f
C13189 net56 _0701_/a_80_21# 0.00349f
C13190 _0812_/a_79_21# _0812_/a_510_47# 0.00844f
C13191 _0812_/a_297_297# _0812_/a_215_47# 0
C13192 _0765_/a_510_47# clknet_1_0__leaf__0457_ 0
C13193 VPWR _0990_/a_27_47# 0.45001f
C13194 _0999_/a_27_47# _0399_ 0
C13195 _0999_/a_193_47# _0398_ 0
C13196 _0369_ _0992_/a_561_413# 0
C13197 net63 net73 0
C13198 _0432_ _0186_ 0.0162f
C13199 net160 net26 0.04007f
C13200 VPWR _1018_/a_1017_47# 0
C13201 _0130_ _0131_ 0
C13202 hold55/a_391_47# comp0.B\[1\] 0
C13203 _0110_ _0720_/a_68_297# 0
C13204 net207 _0178_ 0
C13205 _0083_ _0636_/a_59_75# 0
C13206 _0798_/a_113_297# net41 0
C13207 VPWR _1049_/a_975_413# 0.00478f
C13208 net15 A[4] 0.00408f
C13209 _0224_ _0225_ 0.24494f
C13210 _0500_/a_27_47# net36 0
C13211 net237 _0366_ 0
C13212 clkbuf_0__0463_/a_110_47# _0177_ 0.00587f
C13213 VPWR _0209_ 0.29394f
C13214 _0516_/a_109_297# _0181_ 0.05826f
C13215 net140 hold83/a_49_47# 0.02182f
C13216 _0796_/a_215_47# clkbuf_0__0459_/a_110_47# 0
C13217 net20 hold51/a_49_47# 0.13617f
C13218 _1041_/a_381_47# net31 0.01626f
C13219 hold4/a_285_47# _0103_ 0
C13220 _0647_/a_377_297# VPWR 0.00575f
C13221 _0460_ _1006_/a_466_413# 0.00925f
C13222 VPWR _1066_/a_975_413# 0.00499f
C13223 hold97/a_285_47# _1008_/a_891_413# 0
C13224 net167 _1072_/a_193_47# 0
C13225 acc0.A\[14\] _0400_ 0.09922f
C13226 output67/a_27_47# net67 0.2015f
C13227 hold37/a_285_47# clknet_1_0__leaf__0465_ 0.01245f
C13228 acc0.A\[30\] clknet_1_1__leaf__0462_ 0.07853f
C13229 VPWR _1068_/a_975_413# 0.00418f
C13230 _0964_/a_109_297# _0482_ 0.01416f
C13231 _1053_/a_1059_315# A[4] 0.00163f
C13232 clknet_1_1__leaf__0459_ _0303_ 0.00165f
C13233 _0218_ hold72/a_391_47# 0.07081f
C13234 _0258_ net248 0.01035f
C13235 net149 _0632_/a_113_47# 0
C13236 _1056_/a_27_47# VPWR 0.65003f
C13237 VPWR _0671_/a_113_297# 0.18499f
C13238 hold14/a_285_47# clknet_1_1__leaf__0463_ 0.01635f
C13239 _0993_/a_1059_315# _0091_ 0
C13240 clkbuf_1_0__f__0459_/a_110_47# _0983_/a_27_47# 0
C13241 _0512_/a_27_297# _0512_/a_109_297# 0.17136f
C13242 _0770_/a_79_21# _0770_/a_382_297# 0.00145f
C13243 clknet_1_1__leaf__0463_ input27/a_75_212# 0.0033f
C13244 _0661_/a_277_297# clknet_1_1__leaf__0465_ 0
C13245 _0855_/a_81_21# VPWR 0.20421f
C13246 output54/a_27_47# VPWR 0.24838f
C13247 _0204_ net196 0
C13248 _0140_ _1043_/a_975_413# 0
C13249 clknet_1_0__leaf__0464_ _0148_ 0.05074f
C13250 clknet_1_0__leaf__0465_ _1046_/a_975_413# 0
C13251 _0697_/a_217_297# _0319_ 0.04598f
C13252 _0293_ _0990_/a_1059_315# 0
C13253 _0170_ _1071_/a_561_413# 0
C13254 _0996_/a_466_413# net5 0.02001f
C13255 _0996_/a_193_47# _0185_ 0
C13256 clknet_0_clk _1068_/a_193_47# 0.03839f
C13257 net139 A[5] 0
C13258 _0343_ pp[4] 0
C13259 _0998_/a_466_413# net84 0.01018f
C13260 _0551_/a_27_47# _0178_ 0.14526f
C13261 _1020_/a_634_159# control0.add 0
C13262 net178 _1055_/a_27_47# 0
C13263 _0305_ _0304_ 0
C13264 clknet_1_1__leaf__0459_ _0281_ 0.10435f
C13265 clknet_1_0__leaf__0460_ _0756_/a_285_47# 0
C13266 net38 _0418_ 0
C13267 _0157_ _0459_ 0
C13268 _0396_ _0306_ 0.00158f
C13269 _0159_ _1061_/a_27_47# 0.13017f
C13270 net247 _1061_/a_1059_315# 0
C13271 _0498_/a_51_297# net147 0.0071f
C13272 net7 _1061_/a_466_413# 0
C13273 _0404_ _0403_ 0.34573f
C13274 _0704_/a_68_297# net239 0
C13275 _0984_/a_1059_315# net47 0
C13276 _0096_ _0181_ 0
C13277 clknet_0__0463_ _0474_ 0.01569f
C13278 net190 _0569_/a_109_47# 0
C13279 _0350_ net223 0.3025f
C13280 hold38/a_391_47# _0474_ 0.00206f
C13281 _0176_ _0173_ 0.23354f
C13282 _0478_ clknet_0_clk 0
C13283 _0174_ _1044_/a_1017_47# 0
C13284 _1019_/a_27_47# net207 0.08446f
C13285 _1019_/a_193_47# net105 0.04232f
C13286 _1019_/a_1059_315# _1019_/a_1017_47# 0
C13287 _0714_/a_51_297# _0714_/a_240_47# 0.03076f
C13288 clknet_1_0__leaf__0462_ hold63/a_285_47# 0.00321f
C13289 hold18/a_49_47# _0261_ 0.00393f
C13290 net86 clknet_1_0__leaf__0459_ 0.13866f
C13291 hold42/a_285_47# _0155_ 0.00315f
C13292 net51 _1005_/a_27_47# 0.00115f
C13293 _0467_ comp0.B\[5\] 0
C13294 _0705_/a_59_75# _0334_ 0.00169f
C13295 _0730_/a_215_47# acc0.A\[27\] 0.00915f
C13296 _0553_/a_149_47# clkbuf_1_0__f__0463_/a_110_47# 0
C13297 _1051_/a_466_413# acc0.A\[4\] 0
C13298 hold83/a_285_47# acc0.A\[6\] 0.00838f
C13299 _0548_/a_245_297# net174 0.00291f
C13300 _0726_/a_149_47# _0726_/a_240_47# 0.06872f
C13301 hold9/a_49_47# acc0.A\[28\] 0
C13302 _1058_/a_561_413# net67 0
C13303 hold24/a_391_47# _0207_ 0.0243f
C13304 _0327_ _0332_ 0.44617f
C13305 _0575_/a_109_297# net176 0
C13306 net242 _1010_/a_634_159# 0
C13307 _0533_/a_27_297# _0178_ 0.00381f
C13308 _0182_ _0499_/a_59_75# 0
C13309 net9 net135 0
C13310 _1013_/a_1059_315# _0220_ 0
C13311 hold5/a_285_47# hold5/a_391_47# 0.41909f
C13312 _1015_/a_27_47# _0584_/a_27_297# 0
C13313 hold58/a_49_47# _1035_/a_891_413# 0.0037f
C13314 hold58/a_285_47# _1035_/a_1059_315# 0.01042f
C13315 _0820_/a_79_21# _0179_ 0
C13316 _0655_/a_109_93# hold81/a_285_47# 0
C13317 _1070_/a_27_47# _0976_/a_76_199# 0
C13318 _0982_/a_891_413# _0350_ 0.01606f
C13319 hold38/a_49_47# _1065_/a_27_47# 0.00166f
C13320 acc0.A\[1\] net149 0.12163f
C13321 comp0.B\[5\] comp0.B\[0\] 0
C13322 _0739_/a_79_21# _0739_/a_297_297# 0.01735f
C13323 VPWR _0998_/a_381_47# 0.07064f
C13324 _1020_/a_27_47# hold40/a_49_47# 0
C13325 acc0.A\[29\] hold50/a_391_47# 0
C13326 hold99/a_285_47# _0091_ 0
C13327 clknet_1_0__leaf__0465_ _0987_/a_561_413# 0
C13328 net115 _1028_/a_1059_315# 0
C13329 _1029_/a_27_47# acc0.A\[28\] 0.0062f
C13330 _0347_ _0739_/a_215_47# 0.1226f
C13331 _0990_/a_466_413# clknet_1_1__leaf__0465_ 0
C13332 _0110_ net116 0
C13333 _0347_ _0352_ 1.30991f
C13334 _0465_ _1048_/a_193_47# 0.00371f
C13335 net110 net52 0
C13336 _0965_/a_47_47# VPWR 0.31112f
C13337 _1054_/a_27_47# net9 0
C13338 _0687_/a_59_75# _0106_ 0
C13339 _0292_ _0785_/a_81_21# 0.19509f
C13340 _0990_/a_891_413# _0990_/a_1017_47# 0.00617f
C13341 _0990_/a_193_47# _0088_ 0.41035f
C13342 net125 _0498_/a_51_297# 0.02711f
C13343 _1039_/a_27_47# _0159_ 0.0017f
C13344 _0386_ _0614_/a_29_53# 0.01037f
C13345 net42 _0219_ 0.25927f
C13346 hold81/a_285_47# _0418_ 0
C13347 _0546_/a_51_297# comp0.B\[9\] 0
C13348 _0546_/a_240_47# net127 0
C13349 _1002_/a_561_413# _0460_ 0
C13350 _1002_/a_592_47# clknet_1_0__leaf__0457_ 0
C13351 acc0.A\[2\] _1048_/a_193_47# 0
C13352 _0793_/a_51_297# _0793_/a_149_47# 0.02487f
C13353 acc0.A\[27\] hold8/a_49_47# 0
C13354 _0190_ acc0.A\[10\] 0
C13355 _0315_ acc0.A\[23\] 0.00251f
C13356 _0273_ _0621_/a_35_297# 0
C13357 _0598_/a_79_21# _0237_ 0.03324f
C13358 net42 _0669_/a_111_297# 0
C13359 pp[30] _0720_/a_150_297# 0
C13360 clkbuf_1_0__f__0459_/a_110_47# clknet_0__0459_ 0.3166f
C13361 _0564_/a_68_297# _0175_ 0.10076f
C13362 _0104_ _0352_ 0
C13363 _1050_/a_634_159# _0180_ 0
C13364 _0743_/a_245_297# _0368_ 0
C13365 net233 _0268_ 0.0041f
C13366 acc0.A\[16\] _1060_/a_1059_315# 0
C13367 _0967_/a_403_297# _0476_ 0.01409f
C13368 comp0.B\[7\] _1039_/a_193_47# 0
C13369 comp0.B\[10\] _0139_ 0.00225f
C13370 _0110_ hold92/a_285_47# 0
C13371 net200 _1025_/a_1059_315# 0
C13372 hold68/a_285_47# _0575_/a_27_297# 0.00104f
C13373 _0147_ acc0.A\[3\] 0.02364f
C13374 _1034_/a_193_47# comp0.B\[6\] 0.02868f
C13375 hold21/a_49_47# net63 0.00166f
C13376 _0465_ _0846_/a_149_47# 0.00119f
C13377 hold25/a_285_47# net174 0
C13378 _0343_ _0462_ 0.04575f
C13379 net97 hold80/a_391_47# 0
C13380 _1051_/a_634_159# _1051_/a_1059_315# 0
C13381 _1051_/a_27_47# _1051_/a_381_47# 0.06222f
C13382 _1051_/a_193_47# _1051_/a_891_413# 0.19489f
C13383 net44 VPWR 2.44619f
C13384 clknet_1_1__leaf_clk _0175_ 0
C13385 _1056_/a_466_413# clknet_1_1__leaf__0465_ 0
C13386 _0802_/a_59_75# VPWR 0.23889f
C13387 _0742_/a_384_47# _0219_ 0
C13388 clkbuf_1_0__f__0465_/a_110_47# _0431_ 0.00195f
C13389 acc0.A\[14\] _0849_/a_510_47# 0.00445f
C13390 _0462_ net95 0.00182f
C13391 _1070_/a_466_413# control0.count\[1\] 0.00165f
C13392 _1070_/a_975_413# VPWR 0.00502f
C13393 _1070_/a_381_47# _0168_ 0.12066f
C13394 net106 _1033_/a_381_47# 0
C13395 _1045_/a_193_47# _1045_/a_592_47# 0.00135f
C13396 _1045_/a_466_413# _1045_/a_561_413# 0.00772f
C13397 _1045_/a_634_159# _1045_/a_975_413# 0
C13398 hold90/a_285_47# _0360_ 0.05965f
C13399 _0680_/a_80_21# _0746_/a_299_297# 0
C13400 _0680_/a_217_297# _0746_/a_81_21# 0
C13401 _0584_/a_109_297# _0566_/a_27_47# 0
C13402 _0183_ net177 0.04294f
C13403 VPWR _1043_/a_466_413# 0.2538f
C13404 _0678_/a_68_297# _0394_ 0.05684f
C13405 hold21/a_285_47# net15 0.00362f
C13406 _0294_ _0986_/a_27_47# 0
C13407 _1028_/a_27_47# _0350_ 0
C13408 _1018_/a_193_47# _0399_ 0.00253f
C13409 _1043_/a_466_413# _1043_/a_561_413# 0.00772f
C13410 _1043_/a_634_159# _1043_/a_975_413# 0
C13411 _0573_/a_27_47# _0465_ 0.00259f
C13412 net87 net1 0.00174f
C13413 _0535_/a_150_297# net10 0.00175f
C13414 hold46/a_391_47# _0176_ 0.00417f
C13415 net133 _0532_/a_81_21# 0
C13416 hold88/a_49_47# acc0.A\[8\] 0.0535f
C13417 _0372_ _0219_ 0
C13418 _0195_ clknet_0__0464_ 0
C13419 _0218_ _0264_ 0.03113f
C13420 _1030_/a_193_47# net208 0
C13421 _0384_ clknet_1_0__leaf__0457_ 0
C13422 _1004_/a_975_413# VPWR 0.00516f
C13423 _1021_/a_891_413# _1002_/a_891_413# 0.00316f
C13424 _0518_/a_109_47# _0180_ 0
C13425 _0216_ net239 0
C13426 _1054_/a_634_159# _1054_/a_466_413# 0.23992f
C13427 _1054_/a_193_47# _1054_/a_1059_315# 0.03294f
C13428 _1054_/a_27_47# _1054_/a_891_413# 0.03224f
C13429 _0775_/a_510_47# _0392_ 0.0017f
C13430 _1071_/a_27_47# control0.count\[0\] 0.0066f
C13431 _1071_/a_1059_315# clknet_1_0__leaf_clk 0
C13432 _1015_/a_27_47# _1015_/a_634_159# 0.14145f
C13433 clkbuf_1_0__f__0458_/a_110_47# _0465_ 0.01071f
C13434 hold100/a_285_47# _0182_ 0
C13435 _0983_/a_634_159# VPWR 0.19357f
C13436 acc0.A\[0\] hold60/a_391_47# 0.00101f
C13437 _0234_ net50 0
C13438 _0174_ _1042_/a_891_413# 0.02366f
C13439 _0454_ _0263_ 0
C13440 net182 _0153_ 0
C13441 _0730_/a_79_21# _1010_/a_466_413# 0
C13442 _0730_/a_215_47# _1010_/a_193_47# 0
C13443 net202 net17 0
C13444 _0982_/a_466_413# acc0.A\[1\] 0
C13445 net247 _0631_/a_109_297# 0
C13446 clknet_1_1__leaf__0462_ _1027_/a_27_47# 0.01599f
C13447 pp[27] _0357_ 0
C13448 clknet_1_1__leaf__0463_ net17 0.03082f
C13449 _0987_/a_592_47# _0085_ 0.00188f
C13450 acc0.A\[30\] hold92/a_49_47# 0.00261f
C13451 _0783_/a_215_47# clkbuf_1_1__f__0461_/a_110_47# 0.00246f
C13452 _0689_/a_68_297# _0686_/a_27_53# 0
C13453 _1038_/a_27_47# _1038_/a_466_413# 0.27314f
C13454 _1038_/a_193_47# _1038_/a_634_159# 0.12497f
C13455 _0556_/a_68_297# _1037_/a_193_47# 0.00237f
C13456 _0283_ _0671_/a_113_297# 0
C13457 _0293_ VPWR 0.18469f
C13458 hold88/a_391_47# net76 0.0021f
C13459 _0411_ _0797_/a_27_413# 0
C13460 control0.state\[2\] _1064_/a_1059_315# 0.08429f
C13461 _0676_/a_113_47# _0219_ 0
C13462 _0856_/a_297_297# net47 0
C13463 input13/a_75_212# input14/a_75_212# 0.00176f
C13464 _0218_ net170 0
C13465 _0343_ _0297_ 0
C13466 control0.state\[0\] _1065_/a_27_47# 0
C13467 acc0.A\[8\] _0987_/a_891_413# 0
C13468 net157 _0147_ 0
C13469 _0341_ _0218_ 0.01957f
C13470 pp[29] hold80/a_285_47# 0.02232f
C13471 clknet_1_0__leaf__0458_ _0848_/a_109_297# 0
C13472 _0515_/a_299_297# acc0.A\[10\] 0
C13473 _1059_/a_381_47# _0158_ 0
C13474 _0983_/a_634_159# _0983_/a_381_47# 0
C13475 _0820_/a_215_47# hold67/a_391_47# 0
C13476 clknet_1_0__leaf__0465_ _1051_/a_1059_315# 0.00556f
C13477 clknet_1_0__leaf__0458_ _0294_ 0
C13478 hold38/a_285_47# comp0.B\[4\] 0
C13479 hold88/a_285_47# _0350_ 0
C13480 clknet_1_0__leaf__0465_ _1045_/a_381_47# 0.00187f
C13481 _0758_/a_215_47# _0350_ 0.01307f
C13482 clknet_1_0__leaf__0465_ net139 0.21716f
C13483 net40 _0995_/a_27_47# 0.00545f
C13484 hold98/a_391_47# _0995_/a_466_413# 0.00171f
C13485 hold98/a_49_47# _0995_/a_891_413# 0
C13486 hold29/a_49_47# VPWR 0.32525f
C13487 clkbuf_1_0__f__0461_/a_110_47# _0246_ 0
C13488 VPWR _0566_/a_27_47# 0.42104f
C13489 hold37/a_391_47# net184 0.13581f
C13490 _0985_/a_193_47# net71 0.00616f
C13491 _0200_ net152 0
C13492 _0538_/a_240_47# comp0.B\[12\] 0
C13493 _1002_/a_27_47# net17 0
C13494 _0244_ net223 0
C13495 output64/a_27_47# pp[6] 0.33644f
C13496 _0349_ _0221_ 0
C13497 _0692_/a_113_47# net52 0
C13498 _0087_ output63/a_27_47# 0
C13499 _1015_/a_466_413# _0566_/a_27_47# 0
C13500 _0606_/a_297_297# _0237_ 0
C13501 comp0.B\[8\] net152 0
C13502 _0742_/a_81_21# acc0.A\[23\] 0
C13503 _1056_/a_193_47# hold35/a_285_47# 0.00369f
C13504 _1056_/a_27_47# hold35/a_391_47# 0
C13505 _1056_/a_634_159# hold35/a_49_47# 0.00169f
C13506 _0488_ _1068_/a_27_47# 0
C13507 net90 _1007_/a_27_47# 0
C13508 clknet_1_0__leaf__0459_ _0998_/a_381_47# 0
C13509 _0637_/a_311_297# _0268_ 0.01696f
C13510 acc0.A\[10\] _0091_ 0
C13511 hold97/a_285_47# _0320_ 0
C13512 _0831_/a_35_297# _0369_ 0.01406f
C13513 _0280_ _0644_/a_47_47# 0
C13514 hold33/a_285_47# _1039_/a_27_47# 0
C13515 _1003_/a_1059_315# _0217_ 0.02693f
C13516 net64 hold88/a_49_47# 0.30195f
C13517 acc0.A\[14\] clkbuf_0__0459_/a_110_47# 0.16318f
C13518 net162 net163 0.00554f
C13519 _0330_ _0697_/a_80_21# 0
C13520 _1013_/a_891_413# _0218_ 0.00745f
C13521 _0785_/a_81_21# _0785_/a_299_297# 0.08213f
C13522 _0454_ clknet_1_0__leaf__0461_ 0
C13523 _1016_/a_891_413# _1016_/a_975_413# 0.00851f
C13524 _1016_/a_381_47# _1016_/a_561_413# 0.00123f
C13525 _1004_/a_891_413# net176 0.01107f
C13526 _0331_ _0317_ 0.00522f
C13527 net56 _0330_ 0.04283f
C13528 _0521_/a_384_47# _0180_ 0
C13529 clknet_0__0459_ _0996_/a_193_47# 0.00272f
C13530 _0483_ _0166_ 0
C13531 _0432_ net62 0.03467f
C13532 _0458_ clknet_0__0465_ 0
C13533 acc0.A\[16\] _0294_ 0.00575f
C13534 net113 _1026_/a_193_47# 0.00384f
C13535 _1028_/a_891_413# acc0.A\[28\] 0.01145f
C13536 net49 _0381_ 0
C13537 _0176_ net153 0.00138f
C13538 _0300_ acc0.A\[13\] 0.54924f
C13539 _0329_ _0701_/a_209_297# 0.04399f
C13540 _0476_ hold56/a_285_47# 0
C13541 _0208_ _0560_/a_68_297# 0
C13542 _0203_ hold51/a_285_47# 0.00226f
C13543 _0999_/a_1017_47# _0096_ 0
C13544 _0327_ _0701_/a_209_47# 0
C13545 _0846_/a_51_297# _0263_ 0
C13546 _0343_ _0725_/a_303_47# 0
C13547 hold97/a_391_47# clknet_1_1__leaf__0462_ 0
C13548 _0733_/a_79_199# _0219_ 0.0063f
C13549 _0749_/a_384_47# _0346_ 0.00117f
C13550 clknet_0__0462_ _0360_ 0.04179f
C13551 _0326_ _0745_/a_193_47# 0
C13552 _0514_/a_109_297# net2 0.00625f
C13553 _0455_ net47 0.02902f
C13554 _0179_ _0511_/a_81_21# 0.00365f
C13555 net39 _0994_/a_891_413# 0.0474f
C13556 _0534_/a_81_21# _0534_/a_384_47# 0.00138f
C13557 _0849_/a_79_21# _0347_ 0.00687f
C13558 hold28/a_285_47# _0532_/a_299_297# 0
C13559 _0134_ _1037_/a_193_47# 0
C13560 _1032_/a_634_159# _0352_ 0
C13561 hold62/a_49_47# hold62/a_391_47# 0.00188f
C13562 _1059_/a_381_47# acc0.A\[14\] 0.00519f
C13563 net44 clknet_1_0__leaf__0459_ 0
C13564 _0538_/a_512_297# net20 0
C13565 _1041_/a_381_47# net7 0.01659f
C13566 clknet_1_1__leaf__0459_ _1057_/a_193_47# 0
C13567 _1057_/a_634_159# acc0.A\[11\] 0
C13568 _0403_ _0419_ 0.23271f
C13569 _1002_/a_27_47# acc0.A\[21\] 0
C13570 hold54/a_49_47# _0130_ 0
C13571 hold39/a_49_47# _0561_/a_51_297# 0.06178f
C13572 _0499_/a_59_75# _0495_/a_68_297# 0.00598f
C13573 _0221_ _0701_/a_209_297# 0
C13574 net193 net152 0
C13575 net96 clknet_1_1__leaf__0462_ 0
C13576 _0753_/a_297_297# _0345_ 0.00129f
C13577 input3/a_75_212# net3 0.11645f
C13578 _0663_/a_27_413# _0812_/a_79_21# 0
C13579 _1056_/a_27_47# net182 0.09975f
C13580 _1056_/a_1059_315# _1056_/a_1017_47# 0
C13581 _0323_ _0691_/a_68_297# 0.10601f
C13582 _0744_/a_27_47# net217 0
C13583 _1004_/a_1059_315# hold68/a_285_47# 0
C13584 _0096_ clknet_1_1__leaf__0461_ 0.22219f
C13585 _0734_/a_47_47# _1009_/a_27_47# 0
C13586 _1054_/a_381_47# VPWR 0.07588f
C13587 _0791_/a_199_47# _0406_ 0
C13588 _0108_ net57 0
C13589 _0517_/a_299_297# net16 0.02477f
C13590 output43/a_27_47# _0797_/a_207_413# 0
C13591 _0618_/a_79_21# net52 0
C13592 acc0.A\[5\] _0987_/a_466_413# 0
C13593 clknet_1_0__leaf__0462_ _1025_/a_592_47# 0
C13594 _0601_/a_68_297# clkbuf_1_0__f__0460_/a_110_47# 0
C13595 net53 _0219_ 0.00582f
C13596 _0369_ _1063_/a_193_47# 0
C13597 _0163_ _1065_/a_193_47# 0.53312f
C13598 _0512_/a_373_47# net3 0.00196f
C13599 _0513_/a_81_21# _0511_/a_81_21# 0
C13600 _1038_/a_891_413# VPWR 0.18138f
C13601 _0949_/a_59_75# _0487_ 0.00333f
C13602 _1041_/a_891_413# A[15] 0
C13603 _0222_ net51 0.99566f
C13604 hold39/a_49_47# _0133_ 0.03693f
C13605 VPWR _0655_/a_369_297# 0
C13606 _0446_ net10 0
C13607 _0719_/a_27_47# _0369_ 0.02613f
C13608 _1067_/a_193_47# clknet_1_0__leaf__0457_ 0.04802f
C13609 _0369_ _0460_ 0.11464f
C13610 _0152_ _0518_/a_27_297# 0
C13611 _0983_/a_634_159# clknet_1_0__leaf__0459_ 0
C13612 clknet_1_0__leaf__0460_ _0618_/a_297_297# 0.001f
C13613 _0695_/a_472_297# _0250_ 0.00566f
C13614 _0627_/a_369_297# _0346_ 0
C13615 _0369_ _1060_/a_193_47# 0
C13616 _0374_ _0377_ 0.05134f
C13617 _0241_ _0616_/a_292_297# 0
C13618 hold86/a_391_47# _0264_ 0
C13619 clknet_0__0463_ _0563_/a_51_297# 0.01545f
C13620 clkbuf_1_1__f__0463_/a_110_47# _0563_/a_149_47# 0.00154f
C13621 _0757_/a_68_297# _0757_/a_150_297# 0.00477f
C13622 hold31/a_49_47# _0988_/a_27_47# 0
C13623 _1019_/a_1059_315# clkbuf_1_0__f__0461_/a_110_47# 0
C13624 net56 _1030_/a_27_47# 0
C13625 _1001_/a_891_413# _0216_ 0
C13626 _1031_/a_27_47# _1030_/a_634_159# 0
C13627 _1031_/a_193_47# _1030_/a_193_47# 0
C13628 _1031_/a_634_159# _1030_/a_27_47# 0
C13629 _0714_/a_512_297# _0111_ 0
C13630 _0714_/a_240_47# net225 0.02304f
C13631 _0817_/a_585_47# _0346_ 0
C13632 net35 _1071_/a_561_413# 0
C13633 _1008_/a_634_159# net244 0.00233f
C13634 input6/a_75_212# _0277_ 0
C13635 A[14] _0297_ 0.00154f
C13636 net45 net102 0
C13637 _0179_ _0087_ 0.0026f
C13638 comp0.B\[13\] _1042_/a_891_413# 0
C13639 net245 _0300_ 0
C13640 clknet_0__0457_ _0457_ 0.0117f
C13641 _1012_/a_193_47# _0395_ 0
C13642 _0404_ acc0.A\[13\] 0.02109f
C13643 _1032_/a_27_47# comp0.B\[15\] 0
C13644 _0172_ _0140_ 0.00966f
C13645 _0180_ _0987_/a_634_159# 0
C13646 _0498_/a_51_297# _0497_/a_68_297# 0.00117f
C13647 _0149_ acc0.A\[4\] 0
C13648 _1038_/a_193_47# _0550_/a_149_47# 0
C13649 _0382_ hold3/a_49_47# 0
C13650 _0237_ hold3/a_391_47# 0.03828f
C13651 clknet_1_0__leaf__0460_ _0181_ 0.29198f
C13652 clknet_0_clk clkbuf_1_1__f_clk/a_110_47# 0.36881f
C13653 net43 _0306_ 0.08036f
C13654 _0343_ _0995_/a_561_413# 0
C13655 _0554_/a_68_297# _1037_/a_193_47# 0
C13656 _0712_/a_79_21# _0708_/a_68_297# 0.00133f
C13657 _0551_/a_27_47# comp0.B\[1\] 0
C13658 _1014_/a_975_413# clknet_1_0__leaf__0461_ 0
C13659 net33 _0163_ 0.00157f
C13660 _1025_/a_27_47# _1025_/a_466_413# 0.27314f
C13661 _1025_/a_193_47# _1025_/a_634_159# 0.11949f
C13662 _0858_/a_27_47# _0182_ 0.04567f
C13663 _0354_ net227 0
C13664 clknet_1_1__leaf__0463_ B[2] 0.00183f
C13665 hold64/a_49_47# _0869_/a_27_47# 0.00862f
C13666 _1012_/a_27_47# _0345_ 0
C13667 hold82/a_285_47# _0345_ 0.00167f
C13668 _0330_ _0345_ 0
C13669 comp0.B\[1\] _1032_/a_891_413# 0
C13670 net242 net96 0
C13671 _0287_ _0286_ 0.00462f
C13672 _0199_ _0178_ 0.47443f
C13673 net34 _1064_/a_975_413# 0.00187f
C13674 clknet_0__0465_ clkbuf_1_1__f__0458_/a_110_47# 0.00438f
C13675 hold55/a_285_47# net202 0.00735f
C13676 net233 net222 0
C13677 _0183_ _0461_ 0.06004f
C13678 hold58/a_391_47# _0133_ 0
C13679 VPWR _0522_/a_27_297# 0.21396f
C13680 net187 _0391_ 0
C13681 _1070_/a_27_47# _0488_ 0.00402f
C13682 hold31/a_285_47# clknet_1_1__leaf__0458_ 0
C13683 _1020_/a_381_47# _0181_ 0
C13684 comp0.B\[0\] hold84/a_49_47# 0
C13685 _0347_ hold72/a_285_47# 0.00149f
C13686 _1059_/a_1059_315# net228 0
C13687 _0388_ _0393_ 0
C13688 net214 _0181_ 0
C13689 _0179_ net181 0.11579f
C13690 _0999_/a_27_47# _0306_ 0
C13691 _0739_/a_215_47# _0106_ 0
C13692 _1046_/a_634_159# net10 0.0168f
C13693 clknet_0__0457_ _1001_/a_381_47# 0
C13694 _0467_ _1065_/a_381_47# 0.01676f
C13695 _0515_/a_384_47# _0181_ 0
C13696 _0352_ _0106_ 0
C13697 hold95/a_285_47# hold95/a_391_47# 0.41909f
C13698 _0088_ clknet_1_1__leaf__0465_ 0
C13699 _0396_ _0778_/a_68_297# 0.11141f
C13700 hold86/a_285_47# clknet_1_0__leaf__0458_ 0
C13701 input31/a_75_212# net127 0
C13702 net206 _0632_/a_113_47# 0
C13703 _1003_/a_27_47# control0.state\[2\] 0
C13704 _0996_/a_634_159# _0996_/a_466_413# 0.23992f
C13705 _0996_/a_193_47# _0996_/a_1059_315# 0.03405f
C13706 _0996_/a_27_47# _0996_/a_891_413# 0.03224f
C13707 _0813_/a_109_297# _0181_ 0
C13708 _0195_ _0115_ 0.0033f
C13709 _0174_ _0498_/a_512_297# 0
C13710 A[11] net66 0
C13711 VPWR _0829_/a_109_297# 0.00394f
C13712 _0242_ _0345_ 0
C13713 comp0.B\[1\] _0533_/a_27_297# 0
C13714 _0748_/a_299_297# _0679_/a_68_297# 0
C13715 _0999_/a_891_413# _0219_ 0
C13716 _0999_/a_592_47# _0345_ 0
C13717 clknet_1_0__leaf__0464_ _1048_/a_27_47# 0.00481f
C13718 hold10/a_285_47# clknet_1_1__leaf__0457_ 0.01328f
C13719 output46/a_27_47# net50 0
C13720 net46 output50/a_27_47# 0.00941f
C13721 _0646_/a_285_47# acc0.A\[13\] 0.08625f
C13722 _0646_/a_47_47# net5 0.12101f
C13723 _0159_ _0953_/a_32_297# 0.00303f
C13724 clknet_1_0__leaf__0465_ acc0.A\[8\] 0
C13725 _0376_ _0754_/a_245_297# 0.00163f
C13726 net64 pp[2] 0.00274f
C13727 clknet_1_1__leaf__0463_ _0165_ 0
C13728 hold56/a_49_47# net203 0.00157f
C13729 _0559_/a_512_297# _0175_ 0.00302f
C13730 hold76/a_285_47# _0248_ 0
C13731 _0346_ acc0.A\[10\] 0.00196f
C13732 net136 _0180_ 0
C13733 _0267_ _0449_ 0
C13734 VPWR _0996_/a_381_47# 0.07725f
C13735 hold24/a_49_47# _0553_/a_149_47# 0
C13736 _0317_ _1008_/a_27_47# 0
C13737 _1065_/a_381_47# comp0.B\[0\] 0
C13738 _0274_ _0346_ 0.01694f
C13739 _0726_/a_245_297# acc0.A\[29\] 0
C13740 _0643_/a_253_47# _0640_/a_109_53# 0
C13741 control0.count\[3\] clkbuf_1_0__f_clk/a_110_47# 0.01249f
C13742 _0123_ acc0.A\[25\] 0.13941f
C13743 _1037_/a_975_413# net28 0.00127f
C13744 _0395_ clknet_1_1__leaf__0461_ 0.04021f
C13745 _1051_/a_27_47# acc0.A\[5\] 0
C13746 net66 _0744_/a_27_47# 0.01667f
C13747 _1051_/a_1059_315# net137 0
C13748 _1051_/a_466_413# _0149_ 0.00196f
C13749 hold22/a_391_47# _1054_/a_27_47# 0.0042f
C13750 hold22/a_285_47# _1054_/a_193_47# 0.0148f
C13751 _1045_/a_891_413# _1044_/a_1059_315# 0.00349f
C13752 _1045_/a_1059_315# _1044_/a_891_413# 0.01061f
C13753 _0111_ net41 0
C13754 _0743_/a_240_47# _0250_ 0.0015f
C13755 _0107_ clknet_0__0460_ 0
C13756 _0803_/a_68_297# clknet_1_1__leaf__0459_ 0.00155f
C13757 net58 _0445_ 0.1021f
C13758 _0274_ net65 0.00249f
C13759 _0762_/a_297_297# net51 0.00156f
C13760 _1030_/a_466_413# _0353_ 0
C13761 _0837_/a_266_47# _0346_ 0.01124f
C13762 _0992_/a_466_413# acc0.A\[10\] 0.0066f
C13763 _1051_/a_381_47# net131 0
C13764 _0294_ _0288_ 0
C13765 net62 _0986_/a_381_47# 0.01704f
C13766 net22 _1040_/a_634_159# 0
C13767 net106 comp0.B\[1\] 0.01417f
C13768 _0168_ control0.count\[1\] 0.0648f
C13769 clkbuf_1_0__f__0464_/a_110_47# _0148_ 0.00334f
C13770 net203 _1032_/a_27_47# 0
C13771 net23 _1067_/a_975_413# 0
C13772 net164 clknet_1_0__leaf_clk 0.00514f
C13773 _0101_ hold66/a_49_47# 0.04536f
C13774 _0399_ _0990_/a_634_159# 0.01585f
C13775 _1072_/a_381_47# clknet_1_0__leaf_clk 0
C13776 _0689_/a_68_297# _0320_ 0.10376f
C13777 _0787_/a_80_21# _0993_/a_27_47# 0.0011f
C13778 VPWR net196 0.61353f
C13779 _0298_ input6/a_75_212# 0
C13780 _0714_/a_51_297# net117 0
C13781 net40 _0299_ 0.25158f
C13782 net245 _0404_ 0
C13783 _0984_/a_891_413# _0158_ 0
C13784 _1002_/a_466_413# net240 0
C13785 _1002_/a_27_47# _0165_ 0
C13786 clknet_1_1__leaf__0459_ _0673_/a_337_297# 0
C13787 _0369_ _0796_/a_79_21# 0.1123f
C13788 VPWR _1015_/a_1017_47# 0
C13789 hold49/a_391_47# clknet_1_1__leaf__0464_ 0.00483f
C13790 clknet_1_1__leaf__0459_ _0672_/a_215_47# 0
C13791 clknet_1_1__leaf__0460_ _0776_/a_109_297# 0
C13792 _1003_/a_193_47# _0467_ 0
C13793 _0458_ _0529_/a_109_47# 0
C13794 _0361_ _0323_ 0.00248f
C13795 hold20/a_49_47# net91 0
C13796 clknet_0__0464_ _0540_/a_240_47# 0
C13797 _1030_/a_27_47# _0345_ 0.04085f
C13798 _0362_ acc0.A\[27\] 0.02994f
C13799 clknet_1_0__leaf__0463_ _1040_/a_634_159# 0.00163f
C13800 hold3/a_285_47# _1005_/a_193_47# 0
C13801 _0275_ _0428_ 0.24767f
C13802 VPWR clknet_0_clk 2.40796f
C13803 acc0.A\[1\] net206 0.23234f
C13804 _0294_ _0247_ 0.00265f
C13805 _0119_ _1002_/a_561_413# 0
C13806 _0402_ _0369_ 0
C13807 pp[25] pp[24] 0.09033f
C13808 _1032_/a_193_47# _1032_/a_381_47# 0.10164f
C13809 _1032_/a_634_159# _1032_/a_891_413# 0.03684f
C13810 _1032_/a_27_47# _1032_/a_561_413# 0.0027f
C13811 _1054_/a_634_159# net169 0.03496f
C13812 _1054_/a_466_413# net140 0
C13813 _0568_/a_27_297# _0568_/a_373_47# 0.01338f
C13814 _1015_/a_891_413# _1015_/a_975_413# 0.00851f
C13815 _1015_/a_381_47# _1015_/a_561_413# 0.00123f
C13816 _0717_/a_209_297# hold80/a_285_47# 0
C13817 _0717_/a_80_21# hold80/a_391_47# 0
C13818 _1038_/a_634_159# net29 0
C13819 _0713_/a_27_47# _1015_/a_193_47# 0
C13820 net69 VPWR 0.56663f
C13821 _0557_/a_149_47# _0208_ 0.02934f
C13822 _0357_ _1010_/a_561_413# 0
C13823 _0108_ _1010_/a_1059_315# 0
C13824 _0598_/a_79_21# _0222_ 0
C13825 net68 _0182_ 0.00157f
C13826 _0080_ acc0.A\[1\] 0.06513f
C13827 _0753_/a_381_47# clknet_1_0__leaf__0460_ 0.00118f
C13828 _0198_ net149 0
C13829 _0347_ _0392_ 0.15014f
C13830 _0735_/a_109_297# VPWR 0.00643f
C13831 net65 pp[5] 0
C13832 _0375_ _0228_ 0
C13833 _0405_ _0408_ 0.02723f
C13834 _0343_ _1031_/a_561_413# 0
C13835 net190 _0345_ 0
C13836 _0183_ _0465_ 0.03566f
C13837 _1014_/a_634_159# net149 0.03551f
C13838 _0744_/a_27_47# _0350_ 0.219f
C13839 _1038_/a_27_47# net172 0.08144f
C13840 _1038_/a_193_47# net124 0.00655f
C13841 _1038_/a_1059_315# _1038_/a_1017_47# 0
C13842 net19 _0541_/a_150_297# 0.00147f
C13843 _1039_/a_891_413# _0210_ 0
C13844 _0211_ _1037_/a_891_413# 0
C13845 _0611_/a_68_297# acc0.A\[19\] 0.02791f
C13846 input33/a_75_212# _1066_/a_1059_315# 0
C13847 net33 _1066_/a_27_47# 0.04651f
C13848 hold35/a_285_47# clknet_1_1__leaf__0465_ 0
C13849 hold46/a_285_47# _0548_/a_51_297# 0
C13850 _0312_ net95 0
C13851 net70 _0267_ 0
C13852 _0731_/a_81_21# net216 0
C13853 _0172_ _1043_/a_634_159# 0
C13854 _0319_ _1008_/a_1017_47# 0
C13855 _1067_/a_1059_315# net107 0.00483f
C13856 _1067_/a_381_47# clknet_1_0__leaf__0461_ 0
C13857 input1/a_27_47# init 0.00129f
C13858 _0183_ acc0.A\[2\] 0
C13859 _0655_/a_369_297# _0283_ 0
C13860 pp[30] _0336_ 0.04369f
C13861 _0661_/a_27_297# _0345_ 0.0416f
C13862 _0661_/a_27_297# _0814_/a_27_47# 0
C13863 _0268_ _0849_/a_297_297# 0
C13864 _0637_/a_311_297# net222 0
C13865 _0399_ _0433_ 0
C13866 _0346_ hold73/a_285_47# 0
C13867 clknet_1_0__leaf__0465_ _1044_/a_891_413# 0
C13868 net61 net10 0
C13869 net49 _0468_ 0.00172f
C13870 _0983_/a_381_47# net69 0
C13871 _0490_ _0486_ 0
C13872 net167 control0.state\[2\] 0
C13873 hold16/a_49_47# _1030_/a_27_47# 0.00533f
C13874 hold36/a_49_47# hold36/a_391_47# 0.00188f
C13875 _0289_ _0673_/a_253_297# 0.0066f
C13876 _0287_ _0673_/a_103_199# 0.1394f
C13877 _0661_/a_205_297# _0295_ 0
C13878 net9 _0523_/a_299_297# 0.01079f
C13879 _0854_/a_79_21# _0451_ 0
C13880 _0261_ _0448_ 0.00157f
C13881 net245 _0995_/a_592_47# 0.00147f
C13882 control0.count\[3\] control0.count\[2\] 0
C13883 _0715_/a_27_47# _0275_ 0.09641f
C13884 VPWR _0840_/a_150_297# 0.00211f
C13885 _0137_ _0171_ 0.00176f
C13886 _0461_ hold40/a_285_47# 0.00139f
C13887 _0454_ _0218_ 0.11875f
C13888 _0984_/a_891_413# acc0.A\[14\] 0
C13889 clknet_1_1__leaf__0460_ _1008_/a_193_47# 0
C13890 net31 _0206_ 0.04668f
C13891 hold45/a_285_47# net4 0.00744f
C13892 hold64/a_391_47# clknet_1_0__leaf__0457_ 0.00169f
C13893 _0997_/a_891_413# net42 0.0485f
C13894 hold37/a_285_47# _0148_ 0
C13895 _0550_/a_245_297# _0550_/a_240_47# 0
C13896 _0371_ _1006_/a_27_47# 0
C13897 net216 _1006_/a_193_47# 0
C13898 _0113_ _0566_/a_27_47# 0
C13899 net106 _1032_/a_634_159# 0.00154f
C13900 acc0.A\[12\] _1058_/a_466_413# 0.02907f
C13901 _0226_ _0765_/a_79_21# 0
C13902 _0466_ _1068_/a_1017_47# 0.0016f
C13903 hold32/a_285_47# _1055_/a_193_47# 0.01463f
C13904 hold32/a_391_47# _1055_/a_27_47# 0
C13905 _1048_/a_1059_315# _1047_/a_891_413# 0
C13906 _0467_ _0471_ 0
C13907 _0767_/a_59_75# _0387_ 0.12275f
C13908 net89 _0183_ 0
C13909 hold14/a_285_47# _0556_/a_68_297# 0.00241f
C13910 _1004_/a_1017_47# net50 0.00191f
C13911 _1054_/a_1059_315# acc0.A\[6\] 0
C13912 clkbuf_1_1__f__0462_/a_110_47# _0219_ 0
C13913 _0294_ _0505_/a_109_297# 0.00278f
C13914 _0465_ acc0.A\[15\] 0.19055f
C13915 VPWR _0955_/a_220_297# 0.006f
C13916 _0520_/a_27_297# net12 0
C13917 _0954_/a_32_297# comp0.B\[10\] 0
C13918 _0388_ net206 0
C13919 _0578_/a_27_297# _0352_ 0.01466f
C13920 hold33/a_285_47# _0953_/a_32_297# 0.00299f
C13921 _1061_/a_381_47# acc0.A\[15\] 0
C13922 _0616_/a_78_199# _0246_ 0.07594f
C13923 _0240_ _0614_/a_29_53# 0.08059f
C13924 _1036_/a_193_47# _0175_ 0.00764f
C13925 _0361_ net237 0
C13926 net76 acc0.A\[8\] 0
C13927 acc0.A\[2\] acc0.A\[15\] 0.00252f
C13928 _0998_/a_561_413# _0096_ 0
C13929 _0567_/a_27_297# _0567_/a_109_47# 0.00393f
C13930 _0314_ _0352_ 0
C13931 net21 _0542_/a_51_297# 0
C13932 clknet_0__0458_ _0635_/a_27_47# 0
C13933 net78 _0291_ 0
C13934 net204 _0176_ 0.08475f
C13935 clknet_1_0__leaf__0462_ _0223_ 0
C13936 _0414_ VPWR 0.53167f
C13937 _0354_ net208 0
C13938 clknet_0__0465_ _0291_ 0.0789f
C13939 hold23/a_49_47# _0182_ 0
C13940 clkload0/a_27_47# _1068_/a_1059_315# 0
C13941 hold54/a_285_47# comp0.B\[15\] 0.00398f
C13942 _0471_ comp0.B\[0\] 0
C13943 net97 _1029_/a_27_47# 0
C13944 _0217_ hold4/a_391_47# 0.02878f
C13945 _0183_ hold4/a_49_47# 0.04668f
C13946 acc0.A\[22\] hold4/a_285_47# 0.06432f
C13947 hold86/a_49_47# hold18/a_285_47# 0
C13948 _0172_ net9 0.02762f
C13949 _0328_ clkbuf_1_1__f__0460_/a_110_47# 0.00159f
C13950 _1052_/a_1059_315# net11 0.02328f
C13951 _0216_ net149 0.12925f
C13952 net66 _0350_ 0.55123f
C13953 _0539_/a_68_297# input19/a_75_212# 0
C13954 _0982_/a_27_47# _1014_/a_891_413# 0.00295f
C13955 _0982_/a_193_47# _1014_/a_1059_315# 0.00743f
C13956 _0143_ net20 0
C13957 net21 _0142_ 0
C13958 hold27/a_49_47# _0176_ 0
C13959 _0785_/a_81_21# clkbuf_1_1__f__0465_/a_110_47# 0
C13960 _0195_ _1017_/a_891_413# 0.03457f
C13961 hold64/a_285_47# _1001_/a_891_413# 0
C13962 clk _0978_/a_373_47# 0
C13963 _0179_ net154 0.84025f
C13964 hold42/a_391_47# VPWR 0.16892f
C13965 _0677_/a_47_47# _0394_ 0
C13966 _0677_/a_285_47# _0308_ 0
C13967 _0677_/a_129_47# _0306_ 0
C13968 _1057_/a_891_413# VPWR 0.18236f
C13969 _1048_/a_891_413# _0186_ 0
C13970 VPWR net102 0.39801f
C13971 hold29/a_391_47# net50 0.06786f
C13972 clkbuf_1_1__f__0462_/a_110_47# _1008_/a_634_159# 0
C13973 _0231_ _0377_ 0
C13974 _0233_ net241 0
C13975 _0991_/a_27_47# _0350_ 0.00673f
C13976 _0717_/a_80_21# _0336_ 0.00187f
C13977 _0362_ _1009_/a_634_159# 0.00378f
C13978 _0275_ _0258_ 0.17379f
C13979 acc0.A\[5\] _0085_ 0.17783f
C13980 _0343_ hold78/a_49_47# 0.00189f
C13981 comp0.B\[10\] _0540_/a_245_297# 0
C13982 _0367_ _1007_/a_634_159# 0
C13983 _0366_ _1007_/a_1059_315# 0.07879f
C13984 acc0.A\[17\] _0219_ 0.03163f
C13985 _0188_ net192 0
C13986 net1 _1064_/a_891_413# 0
C13987 _0322_ clknet_0__0460_ 0.33418f
C13988 hold5/a_391_47# net32 0
C13989 _0339_ _0336_ 0.0246f
C13990 comp0.B\[10\] net173 0
C13991 _0179_ _0465_ 0.05427f
C13992 _0805_/a_181_47# _0402_ 0.00295f
C13993 hold69/a_285_47# hold69/a_391_47# 0.41909f
C13994 _1050_/a_1059_315# clknet_1_1__leaf__0464_ 0.00481f
C13995 _0671_/a_113_297# _0345_ 0.00133f
C13996 _0976_/a_76_199# _0976_/a_218_374# 0.00557f
C13997 net35 _0169_ 0
C13998 _0800_/a_51_297# _0800_/a_512_297# 0.0116f
C13999 net28 _0173_ 0
C14000 _0327_ clknet_0__0460_ 0.0125f
C14001 net44 net56 0
C14002 net35 _1072_/a_592_47# 0
C14003 hold57/a_285_47# _0174_ 0.04046f
C14004 _0172_ _0175_ 0.00214f
C14005 hold87/a_391_47# _0268_ 0
C14006 _0313_ _0574_/a_27_297# 0
C14007 _0855_/a_81_21# _0345_ 0.01891f
C14008 _1017_/a_1059_315# _0369_ 0
C14009 _0225_ _1023_/a_634_159# 0
C14010 _1052_/a_1059_315# hold7/a_391_47# 0
C14011 _0152_ _0191_ 0.12891f
C14012 pp[17] _1031_/a_27_47# 0
C14013 _0304_ _0671_/a_199_47# 0
C14014 _0179_ acc0.A\[2\] 0.09198f
C14015 _0473_ comp0.B\[12\] 0.00844f
C14016 VPWR _0699_/a_150_297# 0.00144f
C14017 _0672_/a_510_47# _0303_ 0.00175f
C14018 _0607_/a_109_297# _0352_ 0.05286f
C14019 acc0.A\[14\] hold91/a_391_47# 0.00346f
C14020 _0965_/a_285_47# _0488_ 0
C14021 _0965_/a_129_47# _0466_ 0.00325f
C14022 hold14/a_285_47# _0134_ 0.00315f
C14023 net178 _0988_/a_1059_315# 0.05932f
C14024 _0458_ _0845_/a_193_297# 0.00351f
C14025 _0217_ _0582_/a_109_47# 0.00482f
C14026 _0183_ _0582_/a_27_297# 0.18543f
C14027 _0982_/a_891_413# hold18/a_391_47# 0
C14028 clknet_1_0__leaf__0458_ _0458_ 0.05085f
C14029 _0815_/a_113_297# _0991_/a_466_413# 0
C14030 net64 net76 0
C14031 _0343_ _0129_ 0.12679f
C14032 _1012_/a_27_47# _0394_ 0
C14033 _0983_/a_1059_315# _0399_ 0.04459f
C14034 _0457_ _1067_/a_1017_47# 0
C14035 _0749_/a_81_21# clknet_1_0__leaf__0457_ 0
C14036 net51 _1022_/a_466_413# 0
C14037 net60 _0219_ 0
C14038 hold58/a_391_47# _0208_ 0
C14039 VPWR _0300_ 0.46381f
C14040 clkbuf_1_1__f__0464_/a_110_47# comp0.B\[12\] 0.00868f
C14041 clknet_1_0__leaf__0463_ _1061_/a_891_413# 0
C14042 hold68/a_285_47# net176 0.03672f
C14043 net215 hold29/a_285_47# 0
C14044 hold54/a_285_47# net203 0
C14045 _0428_ _0517_/a_81_21# 0
C14046 _0260_ _0267_ 0
C14047 net5 _0219_ 0.02376f
C14048 hold15/a_285_47# _0705_/a_59_75# 0
C14049 _0498_/a_240_47# _0177_ 0
C14050 _0180_ net73 0
C14051 _0781_/a_68_297# _0094_ 0
C14052 _0523_/a_81_21# _0522_/a_27_297# 0
C14053 _0210_ _1037_/a_891_413# 0.00153f
C14054 net47 _0444_ 0
C14055 _1025_/a_1059_315# _1025_/a_1017_47# 0
C14056 _0201_ net22 0
C14057 _0764_/a_384_47# _0460_ 0
C14058 _1030_/a_193_47# _0221_ 0
C14059 net78 _0290_ 0
C14060 hold69/a_49_47# _0462_ 0.009f
C14061 _0973_/a_27_297# _1067_/a_466_413# 0
C14062 clknet_0__0465_ _0290_ 0
C14063 net55 output55/a_27_47# 0.17858f
C14064 hold25/a_391_47# _0136_ 0
C14065 net69 _0453_ 0
C14066 net149 net247 0.02719f
C14067 _0982_/a_891_413# _0195_ 0.00271f
C14068 VPWR _0193_ 0.30421f
C14069 control0.count\[1\] _0976_/a_439_47# 0
C14070 clk _0972_/a_93_21# 0
C14071 _0516_/a_109_297# clknet_1_1__leaf__0465_ 0
C14072 _0617_/a_68_297# _0617_/a_150_297# 0.00477f
C14073 hold49/a_49_47# comp0.B\[12\] 0.12718f
C14074 hold49/a_285_47# comp0.B\[11\] 0.00198f
C14075 net132 net10 0.0943f
C14076 _0236_ _1006_/a_193_47# 0
C14077 net38 _0417_ 0
C14078 _0467_ control0.reset 0.00165f
C14079 _0119_ _0369_ 0
C14080 _0313_ _0326_ 0
C14081 acc0.A\[14\] _0670_/a_510_47# 0.0046f
C14082 net205 net185 0
C14083 _1055_/a_27_47# _0153_ 0
C14084 _0366_ clkbuf_1_0__f__0462_/a_110_47# 0
C14085 hold57/a_285_47# _0208_ 0.01443f
C14086 _0218_ _0779_/a_79_21# 0.05052f
C14087 VPWR _0827_/a_27_47# 0.00489f
C14088 hold5/a_391_47# net10 0.02961f
C14089 _0174_ _0159_ 0.07558f
C14090 _0402_ _0993_/a_27_47# 0.00296f
C14091 net36 net104 0.00426f
C14092 _0581_/a_109_297# _0247_ 0.00609f
C14093 comp0.B\[5\] control0.sh 0.79304f
C14094 _0123_ net210 0
C14095 net1 hold84/a_49_47# 0
C14096 hold63/a_49_47# acc0.A\[25\] 0.29952f
C14097 hold68/a_49_47# hold68/a_285_47# 0.22264f
C14098 _0820_/a_79_21# _0292_ 0.00111f
C14099 net146 _0505_/a_373_47# 0
C14100 _1052_/a_1059_315# clknet_1_1__leaf__0458_ 0
C14101 acc0.A\[16\] _1016_/a_466_413# 0
C14102 hold79/a_285_47# _0978_/a_27_297# 0.00259f
C14103 _0714_/a_245_297# _0342_ 0.00131f
C14104 hold31/a_49_47# _0642_/a_215_297# 0
C14105 acc0.A\[27\] _0324_ 0
C14106 _0812_/a_297_297# net67 0.00572f
C14107 net37 net228 0.18748f
C14108 clknet_1_0__leaf__0463_ _1039_/a_891_413# 0.00336f
C14109 _1057_/a_975_413# clknet_1_1__leaf__0465_ 0.00126f
C14110 VPWR _1036_/a_561_413# 0.003f
C14111 hold54/a_391_47# _0533_/a_109_297# 0
C14112 _0304_ clkbuf_1_1__f__0459_/a_110_47# 0.00316f
C14113 hold24/a_285_47# _0136_ 0.0111f
C14114 clknet_0__0457_ _0982_/a_1059_315# 0
C14115 control0.reset comp0.B\[0\] 1.05371f
C14116 net98 _0308_ 0
C14117 _0536_/a_149_47# net173 0
C14118 _1044_/a_634_159# _1044_/a_381_47# 0
C14119 _0355_ _0127_ 0
C14120 clkbuf_0__0462_/a_110_47# _0462_ 0.32841f
C14121 hold11/a_285_47# _0536_/a_240_47# 0
C14122 _1038_/a_634_159# comp0.B\[6\] 0.00389f
C14123 _0157_ _0347_ 0
C14124 hold41/a_285_47# _1058_/a_27_47# 0.01543f
C14125 _0815_/a_113_297# _0401_ 0.04832f
C14126 _0815_/a_199_47# _0290_ 0.01065f
C14127 clkload2/Y net132 0.00205f
C14128 _0502_/a_27_47# VPWR 0.37344f
C14129 net131 _1044_/a_561_413# 0
C14130 _0217_ net47 0.3604f
C14131 _0548_/a_240_47# _0206_ 0
C14132 _0512_/a_27_297# net67 0.02102f
C14133 output36/a_27_47# _1038_/a_27_47# 0.03759f
C14134 pp[16] net42 0
C14135 _0999_/a_27_47# _0778_/a_68_297# 0
C14136 net44 _0345_ 0.02661f
C14137 _0108_ clkbuf_1_1__f__0460_/a_110_47# 0.00288f
C14138 _0819_/a_81_21# _0990_/a_27_47# 0
C14139 _0802_/a_59_75# _0345_ 0
C14140 pp[19] _1023_/a_1059_315# 0
C14141 net46 _1023_/a_381_47# 0
C14142 _0195_ _1028_/a_27_47# 0.42253f
C14143 _1067_/a_466_413# net17 0.00576f
C14144 _1051_/a_1059_315# _0148_ 0.00186f
C14145 hold49/a_285_47# _0202_ 0.02177f
C14146 net49 _0762_/a_79_21# 0
C14147 _1057_/a_27_47# _1057_/a_466_413# 0.27314f
C14148 _1057_/a_193_47# _1057_/a_634_159# 0.11072f
C14149 _0404_ VPWR 2.1101f
C14150 _0259_ _0627_/a_369_297# 0
C14151 VPWR _0754_/a_149_47# 0
C14152 clknet_1_0__leaf__0459_ net102 0.01049f
C14153 _0816_/a_68_297# _0346_ 0
C14154 clknet_1_1__leaf__0459_ _0669_/a_29_53# 0.00117f
C14155 _0324_ _0364_ 0
C14156 pp[17] _0712_/a_79_21# 0
C14157 _0100_ net240 0
C14158 _0800_/a_51_297# _0995_/a_193_47# 0
C14159 _0575_/a_109_47# pp[24] 0
C14160 _1059_/a_193_47# _1059_/a_634_159# 0.11072f
C14161 _1059_/a_27_47# _1059_/a_466_413# 0.27314f
C14162 pp[8] pp[1] 0.17991f
C14163 output42/a_27_47# clknet_1_1__leaf__0459_ 0
C14164 _0441_ _0465_ 0
C14165 _0662_/a_384_47# _0424_ 0
C14166 _0458_ _0532_/a_299_297# 0
C14167 _0849_/a_297_297# net222 0
C14168 hold100/a_391_47# net247 0.14418f
C14169 pp[15] input6/a_75_212# 0
C14170 _0517_/a_299_297# net142 0.01363f
C14171 net248 _0987_/a_27_47# 0
C14172 _0310_ _0775_/a_215_47# 0
C14173 net140 net169 0.00163f
C14174 _1032_/a_1059_315# net202 0
C14175 _0568_/a_373_47# _0128_ 0
C14176 _1015_/a_1017_47# _0113_ 0.00147f
C14177 _0344_ _1030_/a_193_47# 0
C14178 net124 net29 0
C14179 _1057_/a_891_413# _0283_ 0
C14180 _0982_/a_466_413# net247 0
C14181 pp[12] pp[13] 0.18478f
C14182 _1032_/a_1059_315# clknet_1_1__leaf__0463_ 0
C14183 _0951_/a_109_93# clknet_1_0__leaf__0457_ 0
C14184 _0569_/a_27_297# _0127_ 0.12525f
C14185 _0569_/a_373_47# acc0.A\[29\] 0.0013f
C14186 acc0.A\[20\] _0604_/a_113_47# 0
C14187 _1065_/a_27_47# clkbuf_1_1__f_clk/a_110_47# 0.00876f
C14188 _0179_ _1058_/a_634_159# 0
C14189 acc0.A\[14\] _0505_/a_109_47# 0.00492f
C14190 hold46/a_49_47# _0540_/a_240_47# 0
C14191 hold46/a_285_47# _0540_/a_149_47# 0
C14192 _0388_ _0773_/a_35_297# 0.26981f
C14193 net100 net149 0.22691f
C14194 _0244_ _0773_/a_285_297# 0
C14195 _0679_/a_68_297# _0246_ 0.16708f
C14196 net44 hold16/a_49_47# 0
C14197 _0718_/a_47_47# _0336_ 0.02255f
C14198 _0172_ net129 0
C14199 control0.add clknet_1_0__leaf__0461_ 0
C14200 hold86/a_391_47# _0846_/a_51_297# 0
C14201 _0551_/a_27_47# _0180_ 0.02707f
C14202 _0343_ _1055_/a_891_413# 0
C14203 _0125_ _1028_/a_193_47# 0.00114f
C14204 acc0.A\[27\] _1028_/a_1059_315# 0.00116f
C14205 comp0.B\[14\] _0954_/a_304_297# 0.00206f
C14206 _0646_/a_285_47# VPWR 0.00547f
C14207 net101 VPWR 0.38541f
C14208 hold11/a_285_47# _1046_/a_27_47# 0.00754f
C14209 _0293_ _0345_ 0.07487f
C14210 _0293_ _0814_/a_27_47# 0.0248f
C14211 _0268_ net170 0.00145f
C14212 hold17/a_49_47# _0488_ 0
C14213 acc0.A\[20\] _0603_/a_68_297# 0.19814f
C14214 acc0.A\[20\] hold73/a_391_47# 0.02797f
C14215 _1052_/a_27_47# _0186_ 0.01154f
C14216 _1020_/a_592_47# net1 0
C14217 _0216_ _0758_/a_79_21# 0
C14218 _1003_/a_193_47# net1 0
C14219 _0997_/a_1017_47# net43 0.00134f
C14220 _0570_/a_109_47# clknet_1_1__leaf__0462_ 0
C14221 _0570_/a_27_297# net113 0.03261f
C14222 acc0.A\[9\] _0347_ 0.30129f
C14223 _0230_ _0103_ 0.04181f
C14224 pp[1] _0988_/a_891_413# 0
C14225 VPWR _0995_/a_592_47# 0
C14226 _0399_ _0266_ 0
C14227 net186 _1033_/a_27_47# 0.00103f
C14228 _0284_ _0993_/a_381_47# 0.0017f
C14229 _0244_ _0350_ 0
C14230 hold78/a_391_47# net45 0.01012f
C14231 clknet_1_1__leaf__0460_ _0318_ 0.06823f
C14232 hold101/a_285_47# acc0.A\[4\] 0
C14233 _0225_ _0377_ 0.0034f
C14234 _0731_/a_81_21# _0370_ 0.03832f
C14235 hold64/a_285_47# net149 0
C14236 clkbuf_1_0__f__0464_/a_110_47# _1048_/a_27_47# 0.00117f
C14237 net7 _0206_ 0.02246f
C14238 VPWR _0228_ 1.32346f
C14239 _0663_/a_297_47# _0290_ 0.00144f
C14240 _0663_/a_207_413# _0401_ 0
C14241 _0663_/a_27_413# _0425_ 0
C14242 _1014_/a_27_47# clkbuf_0__0457_/a_110_47# 0.00287f
C14243 _0458_ hold18/a_49_47# 0
C14244 _1051_/a_381_47# _0525_/a_81_21# 0
C14245 _0259_ _0274_ 0
C14246 _0550_/a_149_47# _0137_ 0
C14247 _0533_/a_27_297# _0180_ 0.14118f
C14248 _0533_/a_109_47# acc0.A\[1\] 0
C14249 _0533_/a_109_297# _0182_ 0.02107f
C14250 _0951_/a_209_311# _1062_/a_634_159# 0
C14251 _0951_/a_109_93# _1062_/a_466_413# 0.0015f
C14252 hold43/a_285_47# net190 0.01022f
C14253 _0179_ clknet_0__0464_ 0.01567f
C14254 net227 _0353_ 0
C14255 control0.state\[0\] clknet_1_0__leaf_clk 0.088f
C14256 acc0.A\[1\] hold71/a_285_47# 0.05843f
C14257 _0182_ hold71/a_49_47# 0.01032f
C14258 _0183_ _1060_/a_634_159# 0.00233f
C14259 hold33/a_285_47# _0174_ 0
C14260 clknet_1_1__leaf__0459_ _0511_/a_81_21# 0
C14261 output65/a_27_47# acc0.A\[8\] 0
C14262 _1000_/a_1017_47# _0461_ 0
C14263 _0511_/a_299_297# acc0.A\[11\] 0.00428f
C14264 _0211_ net27 0.03535f
C14265 _0316_ acc0.A\[27\] 0.03088f
C14266 pp[8] hold34/a_49_47# 0.04883f
C14267 hold65/a_49_47# _0258_ 0.00118f
C14268 hold65/a_391_47# _0257_ 0.00262f
C14269 _0263_ clknet_1_1__leaf__0457_ 0
C14270 _0369_ _0373_ 0.02438f
C14271 _0275_ net72 0.41067f
C14272 _0133_ clkbuf_1_1__f__0463_/a_110_47# 0.06332f
C14273 _1031_/a_27_47# _0567_/a_109_297# 0
C14274 _1031_/a_193_47# _0567_/a_27_297# 0
C14275 _0234_ hold94/a_49_47# 0.00395f
C14276 hold88/a_49_47# _0369_ 0
C14277 _0239_ _0218_ 0
C14278 _0546_/a_245_297# net152 0.0022f
C14279 _0546_/a_149_47# _0205_ 0.00154f
C14280 _0546_/a_51_297# net32 0.10994f
C14281 _1047_/a_891_413# clkbuf_1_1__f__0457_/a_110_47# 0.00988f
C14282 _1047_/a_27_47# clknet_1_1__leaf__0457_ 0.00358f
C14283 _0346_ clknet_0__0460_ 0
C14284 VPWR _1023_/a_561_413# 0.00292f
C14285 clknet_1_1__leaf__0462_ hold50/a_391_47# 0.00586f
C14286 _0991_/a_634_159# _0991_/a_592_47# 0
C14287 _0992_/a_1059_315# _0187_ 0
C14288 comp0.B\[14\] _0540_/a_240_47# 0.00398f
C14289 _0554_/a_150_297# _0208_ 0
C14290 VPWR net16 0.45264f
C14291 _0726_/a_149_47# _0219_ 0.01553f
C14292 acc0.A\[27\] _0347_ 1.09014f
C14293 _0627_/a_297_297# _0186_ 0
C14294 _0370_ _1006_/a_193_47# 0
C14295 _0195_ _0727_/a_193_47# 0
C14296 _0794_/a_110_297# _0300_ 0
C14297 _0997_/a_27_47# clknet_1_1__leaf__0461_ 0
C14298 _0216_ _1029_/a_1059_315# 0.00383f
C14299 hold11/a_391_47# _0177_ 0
C14300 _0210_ _0475_ 0
C14301 clknet_0_clk comp0.B\[3\] 0
C14302 hold78/a_391_47# _0587_/a_27_47# 0
C14303 net48 _0228_ 0.02352f
C14304 _1059_/a_1059_315# _0644_/a_47_47# 0
C14305 _0799_/a_209_297# net5 0
C14306 _0982_/a_466_413# net100 0
C14307 net68 _1014_/a_466_413# 0.00271f
C14308 VPWR _1065_/a_27_47# 0.44512f
C14309 _1004_/a_634_159# acc0.A\[23\] 0
C14310 net82 _0183_ 0.00315f
C14311 _0316_ _0364_ 0
C14312 _0159_ _1046_/a_193_47# 0
C14313 _1001_/a_561_413# _0183_ 0
C14314 _1001_/a_592_47# _0217_ 0
C14315 _0195_ _1016_/a_193_47# 0
C14316 clknet_1_0__leaf__0462_ _0216_ 1.02101f
C14317 net123 _1037_/a_466_413# 0.00158f
C14318 hold47/a_49_47# net134 0
C14319 _0399_ _0996_/a_975_413# 0
C14320 _0984_/a_27_47# _0269_ 0
C14321 net203 _0562_/a_68_297# 0
C14322 _0530_/a_384_47# _0465_ 0
C14323 clkbuf_1_1__f__0462_/a_110_47# net94 0
C14324 B[3] control0.sh 0
C14325 _1021_/a_1059_315# _0183_ 0.00915f
C14326 net1 _0471_ 0.03468f
C14327 _0352_ _0360_ 0
C14328 _0347_ _0364_ 0.12557f
C14329 A[13] net6 0.03022f
C14330 _1060_/a_634_159# acc0.A\[15\] 0
C14331 _0366_ net51 0
C14332 _0174_ net20 0.27897f
C14333 _1058_/a_975_413# acc0.A\[10\] 0
C14334 _0647_/a_47_47# _0301_ 0
C14335 _0367_ net93 0.00713f
C14336 _0315_ _0105_ 0.03015f
C14337 _0099_ _0771_/a_382_47# 0
C14338 _0195_ acc0.A\[4\] 0
C14339 _0546_/a_51_297# _1042_/a_1059_315# 0
C14340 hold57/a_391_47# _0555_/a_51_297# 0
C14341 _0579_/a_109_297# _0713_/a_27_47# 0
C14342 net53 _1007_/a_193_47# 0.0019f
C14343 acc0.A\[6\] net13 0
C14344 _0661_/a_205_297# _0346_ 0
C14345 _0110_ _0347_ 0.222f
C14346 _0976_/a_505_21# _0466_ 0.10334f
C14347 _0388_ _0387_ 0.00128f
C14348 _0800_/a_240_47# _0413_ 0.04691f
C14349 _0800_/a_51_297# _0093_ 0.10258f
C14350 clknet_1_1__leaf__0457_ clknet_1_0__leaf__0461_ 0
C14351 _0279_ net6 0
C14352 _0195_ clkbuf_0__0457_/a_110_47# 0
C14353 _0733_/a_79_199# _0328_ 0.02489f
C14354 _0424_ net47 0
C14355 _0225_ net109 0.03101f
C14356 _0404_ _0283_ 0
C14357 _0508_/a_81_21# net229 0.00396f
C14358 _0180_ _0529_/a_27_297# 0.13493f
C14359 _0655_/a_369_297# _0345_ 0
C14360 net201 _0563_/a_240_47# 0
C14361 _1011_/a_27_47# _1011_/a_466_413# 0.25987f
C14362 _1011_/a_193_47# _1011_/a_634_159# 0.11897f
C14363 _1016_/a_27_47# _0369_ 0.0047f
C14364 VPWR _0830_/a_510_47# 0
C14365 _0713_/a_27_47# _0399_ 0
C14366 net64 output65/a_27_47# 0
C14367 VPWR _0323_ 0.84928f
C14368 _0310_ _0359_ 0
C14369 VPWR init 0.32347f
C14370 _1034_/a_27_47# net23 0
C14371 net232 _0972_/a_250_297# 0
C14372 clknet_0__0465_ _0986_/a_1059_315# 0.00705f
C14373 _0350_ _1006_/a_634_159# 0.03545f
C14374 _0714_/a_51_297# _0216_ 0.00148f
C14375 _0714_/a_512_297# _0195_ 0
C14376 _0216_ _1019_/a_891_413# 0
C14377 _0666_/a_113_47# _0279_ 0
C14378 _0183_ _0115_ 0.01128f
C14379 _0815_/a_113_297# _0089_ 0.05588f
C14380 _0217_ net93 0
C14381 net82 acc0.A\[15\] 0.00842f
C14382 _1021_/a_27_47# hold73/a_49_47# 0
C14383 _1043_/a_891_413# hold51/a_285_47# 0.00163f
C14384 _1043_/a_1059_315# hold51/a_391_47# 0.00124f
C14385 clknet_1_0__leaf__0462_ hold96/a_391_47# 0.0366f
C14386 _0243_ net36 0.00248f
C14387 net51 net151 0
C14388 _0200_ comp0.B\[12\] 0
C14389 _1020_/a_466_413# VPWR 0.25495f
C14390 _0350_ _0986_/a_634_159# 0.00499f
C14391 hold74/a_285_47# _0459_ 0.00473f
C14392 hold12/a_285_47# VPWR 0.31999f
C14393 _0971_/a_299_297# _1063_/a_466_413# 0.00162f
C14394 hold41/a_49_47# pp[9] 0
C14395 net101 clknet_1_0__leaf__0459_ 0.01092f
C14396 _0399_ _0612_/a_59_75# 0
C14397 clk _0975_/a_59_75# 0.02407f
C14398 _0835_/a_215_47# _0255_ 0.04393f
C14399 _0486_ control0.count\[0\] 0
C14400 _0955_/a_32_297# comp0.B\[5\] 0.07655f
C14401 net162 _0220_ 0.07976f
C14402 _0955_/a_220_297# comp0.B\[3\] 0
C14403 net53 _0328_ 0.14507f
C14404 clkbuf_1_0__f__0461_/a_110_47# _0264_ 0
C14405 _0404_ _0794_/a_110_297# 0.00898f
C14406 _0789_/a_544_297# _0297_ 0.00143f
C14407 _0789_/a_75_199# _0300_ 0.17692f
C14408 _0305_ _0748_/a_81_21# 0
C14409 _0680_/a_80_21# _0294_ 0.16261f
C14410 _0523_/a_81_21# _0193_ 0.19233f
C14411 _0609_/a_109_297# _0248_ 0
C14412 _0429_ hold65/a_391_47# 0
C14413 _0216_ net206 0
C14414 _1025_/a_975_413# acc0.A\[25\] 0
C14415 clknet_1_1__leaf__0459_ _0799_/a_80_21# 0.00452f
C14416 net65 _0828_/a_113_297# 0.00255f
C14417 control0.count\[3\] clkload0/a_27_47# 0
C14418 net55 _1010_/a_634_159# 0
C14419 _1020_/a_381_47# _1015_/a_27_47# 0
C14420 _1020_/a_27_47# _1015_/a_381_47# 0
C14421 net70 _0347_ 0
C14422 _0163_ _0880_/a_27_47# 0
C14423 hold101/a_391_47# clknet_1_0__leaf__0465_ 0.03126f
C14424 _0165_ _1067_/a_466_413# 0.02519f
C14425 _0179_ _1060_/a_634_159# 0
C14426 control0.state\[2\] _0974_/a_448_47# 0
C14427 _0486_ _0974_/a_544_297# 0.0027f
C14428 clkbuf_0__0463_/a_110_47# _0495_/a_68_297# 0.00648f
C14429 net54 _1008_/a_381_47# 0
C14430 _0217_ _0294_ 0.0381f
C14431 net39 pp[12] 0.01592f
C14432 _0255_ _0523_/a_299_297# 0
C14433 clknet_0__0457_ _1019_/a_381_47# 0.00127f
C14434 _1010_/a_193_47# _0347_ 0.03585f
C14435 net43 net221 0
C14436 net125 _0181_ 0
C14437 _0159_ comp0.B\[9\] 0
C14438 _1051_/a_193_47# clknet_1_1__leaf__0464_ 0.00338f
C14439 hold63/a_49_47# net210 0
C14440 _0800_/a_149_47# _0404_ 0
C14441 net55 _1009_/a_466_413# 0
C14442 _0368_ hold90/a_49_47# 0
C14443 _0959_/a_80_21# _0164_ 0
C14444 VPWR _0419_ 0.23093f
C14445 _1045_/a_466_413# clknet_1_1__leaf__0464_ 0
C14446 _1036_/a_193_47# _1036_/a_381_47# 0.0982f
C14447 _1036_/a_634_159# _1036_/a_891_413# 0.03684f
C14448 _1036_/a_27_47# _1036_/a_561_413# 0.0027f
C14449 _0090_ net37 0
C14450 _0290_ _0986_/a_27_47# 0
C14451 net84 _0219_ 0
C14452 _0346_ _0990_/a_634_159# 0
C14453 _1030_/a_891_413# hold61/a_391_47# 0.00323f
C14454 control0.sh hold84/a_49_47# 0.29171f
C14455 _0517_/a_299_297# _0988_/a_27_47# 0
C14456 _0517_/a_81_21# _0988_/a_193_47# 0
C14457 _1012_/a_634_159# _0778_/a_68_297# 0
C14458 _0578_/a_27_297# _0578_/a_373_47# 0.01338f
C14459 _1049_/a_634_159# net11 0
C14460 _0591_/a_109_297# _0223_ 0.0122f
C14461 _0725_/a_209_297# _0725_/a_209_47# 0
C14462 _0725_/a_80_21# _0725_/a_303_47# 0.01146f
C14463 _0274_ _0253_ 0.16073f
C14464 net248 clkbuf_1_0__f__0465_/a_110_47# 0.02606f
C14465 acc0.A\[16\] net166 0.02821f
C14466 _0463_ clkbuf_1_0__f__0463_/a_110_47# 0.02426f
C14467 pp[28] _0723_/a_207_413# 0.00848f
C14468 _0176_ _0205_ 0.03979f
C14469 _0966_/a_109_297# _0966_/a_27_47# 0
C14470 net133 clknet_1_1__leaf__0457_ 0.02558f
C14471 net3 net37 0.16257f
C14472 _0595_/a_109_297# _0217_ 0.00145f
C14473 _0796_/a_297_297# acc0.A\[15\] 0
C14474 net44 _0394_ 0
C14475 _0654_/a_27_413# _0419_ 0
C14476 _0654_/a_297_47# _0417_ 0
C14477 _1044_/a_381_47# net130 0.0013f
C14478 _0195_ net41 0
C14479 _0210_ net27 0.00113f
C14480 net193 comp0.B\[12\] 0
C14481 output36/a_27_47# B[6] 0.01105f
C14482 hold33/a_285_47# comp0.B\[13\] 0
C14483 _1041_/a_1059_315# hold6/a_49_47# 0.001f
C14484 _1041_/a_634_159# hold6/a_391_47# 0.00123f
C14485 _1041_/a_466_413# hold6/a_285_47# 0
C14486 _0137_ _0494_/a_27_47# 0
C14487 net124 comp0.B\[6\] 0
C14488 hold69/a_49_47# _0312_ 0.02329f
C14489 _0965_/a_47_47# _0490_ 0
C14490 control0.count\[3\] _0981_/a_27_297# 0
C14491 _0985_/a_975_413# _0465_ 0
C14492 _0163_ _1062_/a_27_47# 0
C14493 clknet_1_0__leaf__0462_ _1024_/a_193_47# 0.0043f
C14494 _0467_ _1063_/a_193_47# 0.03936f
C14495 VPWR net237 0.16122f
C14496 _1058_/a_27_47# net4 0.07437f
C14497 _0869_/a_27_47# acc0.A\[19\] 0.12103f
C14498 _1021_/a_27_47# _0181_ 0.03408f
C14499 _0399_ _0516_/a_27_297# 0
C14500 _0483_ _0962_/a_109_297# 0
C14501 _0326_ clkbuf_0__0460_/a_110_47# 0.02753f
C14502 VPWR _0843_/a_150_297# 0.00123f
C14503 net36 _1038_/a_975_413# 0
C14504 pp[0] _1038_/a_381_47# 0
C14505 clknet_1_1__leaf_clk _1065_/a_1017_47# 0
C14506 _1049_/a_891_413# _0465_ 0
C14507 _0803_/a_68_297# _0803_/a_150_297# 0.00477f
C14508 _0329_ _0354_ 0
C14509 _0353_ net208 0
C14510 _1012_/a_1059_315# _0720_/a_68_297# 0.00168f
C14511 net224 hold77/a_49_47# 0.00134f
C14512 _0428_ _0990_/a_466_413# 0
C14513 _0427_ _0990_/a_1059_315# 0
C14514 hold86/a_285_47# _0448_ 0.03424f
C14515 _0585_/a_27_297# clknet_1_1__leaf__0457_ 0.00117f
C14516 pp[27] _0356_ 0
C14517 net46 acc0.A\[23\] 0.16983f
C14518 hold34/a_391_47# _0186_ 0
C14519 _1054_/a_27_47# _0989_/a_27_47# 0.00206f
C14520 _0467_ _0460_ 0.00803f
C14521 _0255_ _0172_ 0
C14522 hold20/a_49_47# _0217_ 0
C14523 _0736_/a_139_47# _0363_ 0
C14524 _0570_/a_27_297# hold8/a_285_47# 0
C14525 _0327_ _0355_ 0
C14526 _1057_/a_27_47# net189 0.09365f
C14527 _1057_/a_1059_315# _1057_/a_1017_47# 0
C14528 _0378_ net51 0.06894f
C14529 acc0.A\[2\] _1049_/a_891_413# 0
C14530 _0174_ clkbuf_1_1__f__0463_/a_110_47# 0
C14531 _0269_ _0986_/a_561_413# 0
C14532 net63 _0524_/a_27_297# 0
C14533 net59 _0352_ 0.00684f
C14534 _0195_ _0534_/a_299_297# 0.05586f
C14535 VPWR _1064_/a_1017_47# 0
C14536 _0209_ net171 0.03446f
C14537 _0607_/a_109_47# clknet_0__0461_ 0
C14538 _0579_/a_27_297# _0579_/a_109_47# 0.00393f
C14539 net57 hold62/a_391_47# 0
C14540 _0433_ _0346_ 0
C14541 _0195_ hold62/a_285_47# 0.01274f
C14542 _1059_/a_1059_315# _1059_/a_1017_47# 0
C14543 _1059_/a_193_47# net145 0.004f
C14544 _1059_/a_27_47# _0157_ 0.11969f
C14545 _0789_/a_75_199# _0404_ 0.19852f
C14546 comp0.B\[0\] _1063_/a_193_47# 0
C14547 hold78/a_391_47# VPWR 0.1654f
C14548 _0528_/a_299_297# net170 0.05874f
C14549 _0568_/a_109_297# _0219_ 0.00713f
C14550 _0510_/a_27_297# _0186_ 0.11662f
C14551 _0218_ control0.add 0.06605f
C14552 _0981_/a_373_47# VPWR 0
C14553 net65 _0433_ 0.01259f
C14554 _0221_ _0354_ 0.20448f
C14555 _0181_ _1047_/a_1059_315# 0
C14556 _0710_/a_109_297# _0341_ 0.00179f
C14557 _0176_ _1042_/a_193_47# 0
C14558 _0080_ net247 0
C14559 _0312_ clkbuf_0__0462_/a_110_47# 0.00136f
C14560 net214 clknet_1_1__leaf__0465_ 0.03804f
C14561 clknet_1_0__leaf_clk _1068_/a_193_47# 0.00265f
C14562 _0673_/a_337_297# _0673_/a_253_47# 0.00219f
C14563 _0209_ net24 0
C14564 _0179_ net144 0.25779f
C14565 clknet_1_1__leaf__0460_ _1007_/a_27_47# 0
C14566 comp0.B\[13\] net20 0.26363f
C14567 net69 _0345_ 0
C14568 _0369_ _0761_/a_113_47# 0
C14569 _0672_/a_215_47# _0672_/a_510_47# 0.00529f
C14570 comp0.B\[6\] _0494_/a_27_47# 0.00943f
C14571 _0210_ _0136_ 0
C14572 _0693_/a_68_297# clknet_1_0__leaf__0460_ 0
C14573 _0398_ _0096_ 0.00756f
C14574 _1030_/a_891_413# clknet_1_1__leaf__0462_ 0
C14575 hold32/a_285_47# pp[8] 0.03908f
C14576 hold65/a_391_47# clknet_1_1__leaf__0458_ 0.0045f
C14577 _0284_ _0403_ 0.01954f
C14578 net83 _0405_ 0.0016f
C14579 VPWR _0686_/a_27_53# 0.0765f
C14580 _0530_/a_81_21# _0509_/a_27_47# 0
C14581 _0715_/a_27_47# _0990_/a_466_413# 0
C14582 _1054_/a_466_413# _0087_ 0
C14583 VPWR _1008_/a_891_413# 0.18718f
C14584 _0478_ clknet_1_0__leaf_clk 0.67233f
C14585 net163 VPWR 0.4019f
C14586 _0180_ _0196_ 0.02497f
C14587 _0182_ net170 0
C14588 clknet_1_0__leaf__0465_ _0369_ 0
C14589 net158 _1046_/a_891_413# 0
C14590 _0335_ _0723_/a_27_413# 0.20762f
C14591 _0309_ _0218_ 0
C14592 _0457_ comp0.B\[0\] 0.00718f
C14593 _0958_/a_27_47# _0951_/a_209_311# 0
C14594 _0467_ _1062_/a_891_413# 0
C14595 net21 net198 0
C14596 _0576_/a_27_297# hold29/a_391_47# 0.00398f
C14597 net46 _0602_/a_113_47# 0
C14598 _0124_ _0352_ 0
C14599 acc0.A\[13\] _0668_/a_297_47# 0
C14600 clknet_1_0__leaf__0458_ acc0.A\[1\] 0.12285f
C14601 _0126_ net113 0.00113f
C14602 _0438_ _0434_ 0.01858f
C14603 _0305_ _1017_/a_193_47# 0
C14604 _0341_ _1013_/a_27_47# 0
C14605 _0179_ hold47/a_285_47# 0.00408f
C14606 net101 _0113_ 0.00341f
C14607 net144 _0513_/a_81_21# 0
C14608 _1058_/a_975_413# _0188_ 0
C14609 clknet_0__0463_ _0173_ 0.81672f
C14610 clkbuf_1_1__f__0463_/a_110_47# _0208_ 0.18672f
C14611 _0408_ hold91/a_285_47# 0
C14612 _0181_ _0186_ 1.51617f
C14613 _0299_ _0995_/a_27_47# 0.01233f
C14614 _0454_ _0268_ 0
C14615 hold38/a_391_47# _0173_ 0.00117f
C14616 _0460_ _0374_ 0.00178f
C14617 hold33/a_285_47# comp0.B\[9\] 0.04445f
C14618 _1010_/a_27_47# hold95/a_285_47# 0
C14619 _1010_/a_193_47# hold95/a_49_47# 0
C14620 acc0.A\[24\] net51 0
C14621 _1039_/a_193_47# comp0.B\[2\] 0
C14622 clknet_1_0__leaf__0462_ _0577_/a_27_297# 0.02436f
C14623 _0180_ _0199_ 0.18487f
C14624 control0.state\[1\] clk 0.41578f
C14625 comp0.B\[0\] _1062_/a_891_413# 0
C14626 _0274_ output61/a_27_47# 0
C14627 hold69/a_285_47# _0219_ 0
C14628 _0183_ net146 0.2391f
C14629 _0199_ net218 0
C14630 hold19/a_49_47# _0181_ 0
C14631 _0163_ net107 0
C14632 clknet_0__0458_ net233 0.00179f
C14633 _1014_/a_27_47# _0350_ 0
C14634 net204 net28 0.08644f
C14635 hold28/a_391_47# clknet_1_1__leaf__0457_ 0
C14636 VPWR _0563_/a_512_297# 0.00609f
C14637 B[8] _0546_/a_149_47# 0
C14638 _0190_ A[9] 0
C14639 control0.state\[1\] _1063_/a_891_413# 0.03642f
C14640 net207 _1014_/a_1059_315# 0
C14641 net105 _1014_/a_891_413# 0
C14642 hold44/a_49_47# hold44/a_285_47# 0.22264f
C14643 clknet_1_0__leaf__0462_ _1022_/a_592_47# 0
C14644 _1005_/a_634_159# _1005_/a_381_47# 0
C14645 pp[15] pp[18] 0
C14646 _0731_/a_81_21# _0731_/a_384_47# 0.00138f
C14647 net182 net16 0
C14648 _0984_/a_27_47# _0082_ 0.12476f
C14649 _0984_/a_466_413# net222 0
C14650 _1066_/a_27_47# _1062_/a_27_47# 0.07618f
C14651 _1060_/a_27_47# _0507_/a_109_297# 0
C14652 _1060_/a_193_47# _0507_/a_27_297# 0
C14653 _1013_/a_634_159# _1013_/a_466_413# 0.23992f
C14654 _1013_/a_193_47# _1013_/a_1059_315# 0.03405f
C14655 _1013_/a_27_47# _1013_/a_891_413# 0.03224f
C14656 acc0.A\[27\] _0106_ 0.08683f
C14657 _0991_/a_891_413# net67 0.00338f
C14658 _1002_/a_27_47# _1002_/a_193_47# 0.96639f
C14659 _0351_ net209 0
C14660 _0216_ _0356_ 0.00118f
C14661 _0309_ _0775_/a_215_47# 0
C14662 _0181_ clknet_0__0462_ 0
C14663 net243 _0347_ 0.00255f
C14664 _0424_ _0294_ 0.20356f
C14665 _0617_/a_68_297# _0219_ 0
C14666 _0315_ _0359_ 0.26151f
C14667 _0366_ _0324_ 0.11952f
C14668 _0830_/a_297_297# acc0.A\[6\] 0.00559f
C14669 _0985_/a_381_47# _0261_ 0
C14670 _0985_/a_891_413# _0263_ 0
C14671 clknet_1_1__leaf__0459_ _0997_/a_1059_315# 0.00978f
C14672 _1017_/a_27_47# net43 0
C14673 _0283_ _0419_ 0
C14674 net165 _1060_/a_193_47# 0
C14675 _0770_/a_382_297# _0461_ 0
C14676 _0574_/a_373_47# _0216_ 0.0023f
C14677 clknet_1_1__leaf__0459_ _0992_/a_975_413# 0
C14678 _0414_ _0345_ 0
C14679 VPWR _0989_/a_193_47# 0.31294f
C14680 hold32/a_49_47# pp[9] 0.00655f
C14681 net150 net240 0
C14682 _0358_ _0317_ 0
C14683 VPWR hold1/a_285_47# 0.28365f
C14684 _0475_ comp0.B\[0\] 0
C14685 _0274_ _0642_/a_382_47# 0.00367f
C14686 net178 net235 0
C14687 _0080_ net100 0
C14688 hold64/a_285_47# _1019_/a_891_413# 0.00152f
C14689 hold64/a_391_47# _1019_/a_1059_315# 0
C14690 _1038_/a_891_413# _1040_/a_27_47# 0
C14691 _1038_/a_1059_315# _1040_/a_193_47# 0
C14692 _1012_/a_1059_315# hold92/a_285_47# 0.00451f
C14693 VPWR _0992_/a_193_47# 0.31835f
C14694 _0600_/a_253_47# _0223_ 0.03636f
C14695 _0600_/a_103_199# _0232_ 0.08045f
C14696 hold56/a_285_47# hold39/a_391_47# 0
C14697 hold56/a_391_47# hold39/a_285_47# 0
C14698 _0216_ comp0.B\[15\] 0
C14699 _0183_ net223 0
C14700 _0764_/a_384_47# _0373_ 0.01051f
C14701 comp0.B\[10\] net19 0
C14702 net123 _0135_ 0.01033f
C14703 _0768_/a_109_297# _0347_ 0
C14704 _0719_/a_27_47# acc0.A\[19\] 0.04823f
C14705 comp0.B\[9\] net20 0
C14706 _0995_/a_634_159# _0995_/a_592_47# 0
C14707 _0328_ clkbuf_1_1__f__0462_/a_110_47# 0
C14708 hold10/a_391_47# VPWR 0.17682f
C14709 clknet_1_0__leaf__0457_ _0242_ 0
C14710 hold76/a_391_47# net46 0.07459f
C14711 _0106_ _0364_ 0
C14712 _0357_ _0333_ 0.06944f
C14713 _0820_/a_79_21# clkbuf_1_1__f__0465_/a_110_47# 0.0075f
C14714 clknet_1_1__leaf__0463_ _0560_/a_68_297# 0
C14715 _0991_/a_1059_315# acc0.A\[9\] 0
C14716 _0343_ _0582_/a_109_47# 0.00248f
C14717 hold59/a_285_47# acc0.A\[18\] 0.00795f
C14718 net146 acc0.A\[15\] 0.05628f
C14719 _0983_/a_1059_315# _0346_ 0.00146f
C14720 hold18/a_391_47# _0350_ 0.04103f
C14721 _1070_/a_466_413# _0489_ 0
C14722 _1034_/a_27_47# _0213_ 0.02453f
C14723 _1034_/a_1059_315# _0561_/a_149_47# 0
C14724 _1017_/a_634_159# _0675_/a_68_297# 0
C14725 hold64/a_285_47# net206 0.00274f
C14726 _0217_ _0581_/a_109_297# 0.02081f
C14727 net36 net180 0
C14728 VPWR _0427_ 0.39137f
C14729 net32 _1042_/a_891_413# 0.03028f
C14730 _0139_ _1042_/a_634_159# 0
C14731 _1018_/a_466_413# _0459_ 0.00305f
C14732 _0168_ _1069_/a_27_47# 0
C14733 VPWR _1069_/a_634_159# 0.18215f
C14734 _1070_/a_193_47# clknet_1_0__leaf_clk 0.02259f
C14735 control0.state\[1\] _1062_/a_592_47# 0
C14736 VPWR hold60/a_285_47# 0.28362f
C14737 output64/a_27_47# hold31/a_285_47# 0
C14738 _0268_ _0846_/a_51_297# 0.00111f
C14739 _0982_/a_891_413# _0183_ 0.00364f
C14740 hold27/a_285_47# net173 0
C14741 _1034_/a_466_413# _0472_ 0
C14742 _0299_ _0399_ 0
C14743 comp0.B\[12\] _1045_/a_193_47# 0
C14744 net8 _0560_/a_68_297# 0
C14745 _0695_/a_80_21# _0743_/a_51_297# 0
C14746 _0622_/a_193_47# _0252_ 0.00506f
C14747 _1011_/a_193_47# net97 0.00544f
C14748 _1011_/a_1059_315# _1011_/a_1017_47# 0
C14749 input2/a_75_212# acc0.A\[10\] 0.0016f
C14750 VPWR input24/a_75_212# 0.1893f
C14751 _0272_ net62 0.00617f
C14752 _0985_/a_193_47# _0186_ 0.06528f
C14753 _1000_/a_27_47# _0614_/a_29_53# 0
C14754 _0465_ _0171_ 0.00523f
C14755 _0133_ _1034_/a_561_413# 0
C14756 _0274_ _0446_ 0
C14757 _0182_ _0532_/a_81_21# 0.0369f
C14758 acc0.A\[1\] _0532_/a_299_297# 0
C14759 _0195_ _0350_ 0.11461f
C14760 _0719_/a_27_47# _0249_ 0
C14761 _1006_/a_193_47# _1006_/a_466_413# 0.07482f
C14762 _1006_/a_27_47# _1006_/a_1059_315# 0.04755f
C14763 _0179_ comp0.B\[14\] 0
C14764 net232 _0164_ 0.0011f
C14765 _0538_/a_245_297# VPWR 0.00471f
C14766 _0350_ net92 0.13421f
C14767 _0226_ _0764_/a_299_297# 0
C14768 _0111_ _0195_ 0.03693f
C14769 _0249_ _0460_ 0.03456f
C14770 _0972_/a_346_47# _0487_ 0
C14771 _0316_ hold97/a_285_47# 0
C14772 _0984_/a_27_47# _0984_/a_193_47# 0.96557f
C14773 _0201_ _1043_/a_193_47# 0
C14774 clknet_1_0__leaf__0462_ _0756_/a_377_297# 0
C14775 _0212_ _1034_/a_27_47# 0
C14776 _0124_ _1025_/a_466_413# 0
C14777 _0808_/a_81_21# _0808_/a_368_297# 0.01485f
C14778 _1055_/a_561_413# VPWR 0.00332f
C14779 _0118_ VPWR 0.37938f
C14780 net76 _0369_ 0.03262f
C14781 _1001_/a_1059_315# _0242_ 0
C14782 _1003_/a_381_47# VPWR 0.07615f
C14783 _0982_/a_27_47# _0117_ 0
C14784 hold77/a_49_47# hold77/a_391_47# 0.00188f
C14785 hold97/a_49_47# _0739_/a_79_21# 0
C14786 _0955_/a_32_297# hold84/a_49_47# 0
C14787 net98 hold92/a_391_47# 0
C14788 pp[26] clknet_1_1__leaf__0462_ 0
C14789 net54 net113 0
C14790 net35 _1068_/a_1059_315# 0.09743f
C14791 comp0.B\[5\] _0474_ 0.01264f
C14792 hold97/a_285_47# _0347_ 0
C14793 _0712_/a_79_21# _1031_/a_27_47# 0.00238f
C14794 hold74/a_391_47# _0218_ 0
C14795 _0986_/a_193_47# _0986_/a_466_413# 0.07482f
C14796 _0986_/a_27_47# _0986_/a_1059_315# 0.04875f
C14797 net148 _0987_/a_1059_315# 0
C14798 _0300_ _0345_ 0.00449f
C14799 _0361_ clkbuf_1_0__f__0462_/a_110_47# 0.00164f
C14800 net236 _0466_ 0.1182f
C14801 clknet_0__0458_ _0637_/a_311_297# 0
C14802 net55 net96 0.18028f
C14803 _1020_/a_466_413# _0113_ 0
C14804 _0118_ _1015_/a_466_413# 0
C14805 _1017_/a_193_47# _0181_ 0.09837f
C14806 _1023_/a_27_47# _1023_/a_561_413# 0.0027f
C14807 _1023_/a_634_159# _1023_/a_891_413# 0.03684f
C14808 _1023_/a_193_47# _1023_/a_381_47# 0.09799f
C14809 _0179_ net146 0
C14810 _0344_ _0567_/a_27_297# 0.01004f
C14811 _0304_ _0277_ 0
C14812 _1042_/a_1059_315# _1042_/a_891_413# 0.31086f
C14813 _1042_/a_193_47# _1042_/a_975_413# 0
C14814 _1042_/a_466_413# _1042_/a_381_47# 0.03733f
C14815 hold59/a_49_47# hold59/a_285_47# 0.22264f
C14816 acc0.A\[14\] net42 0.06507f
C14817 clknet_1_0__leaf__0458_ net77 0.10833f
C14818 _0181_ _1060_/a_592_47# 0.00191f
C14819 control0.add _0099_ 0.02003f
C14820 _0175_ _0214_ 0.00125f
C14821 _0516_/a_27_297# _0190_ 0.11367f
C14822 _0516_/a_109_47# net16 0.00149f
C14823 _0290_ _0288_ 0.00471f
C14824 _0425_ acc0.A\[9\] 0.03511f
C14825 clknet_1_1__leaf__0464_ _1044_/a_634_159# 0.03972f
C14826 comp0.B\[15\] net247 0
C14827 _0459_ acc0.A\[13\] 0.0017f
C14828 _0343_ net47 3.27134f
C14829 pp[16] net60 0.01489f
C14830 _1017_/a_466_413# _0307_ 0.00212f
C14831 net9 _1061_/a_1059_315# 0
C14832 _0179_ _1050_/a_381_47# 0
C14833 _0093_ _0298_ 0.00169f
C14834 net184 clknet_1_1__leaf__0464_ 0
C14835 _0458_ _0448_ 0
C14836 _1039_/a_381_47# _0171_ 0
C14837 comp0.B\[3\] _1065_/a_27_47# 0.00284f
C14838 _1036_/a_193_47# comp0.B\[4\] 0.0015f
C14839 _1036_/a_1059_315# net161 0
C14840 _0466_ _1064_/a_193_47# 0
C14841 _0852_/a_35_297# _0350_ 0
C14842 net120 _1033_/a_27_47# 0.00484f
C14843 hold18/a_49_47# acc0.A\[1\] 0
C14844 net70 _1059_/a_27_47# 0
C14845 _0984_/a_27_47# net145 0
C14846 _0230_ hold66/a_49_47# 0
C14847 _0153_ _0988_/a_1059_315# 0
C14848 _0107_ hold77/a_285_47# 0
C14849 _0399_ _0619_/a_68_297# 0
C14850 net55 _0315_ 0
C14851 _0716_/a_27_47# _0402_ 0
C14852 pp[29] _1011_/a_27_47# 0
C14853 _1057_/a_193_47# _0511_/a_299_297# 0
C14854 _0992_/a_1059_315# clknet_1_1__leaf__0465_ 0
C14855 VPWR _1040_/a_561_413# 0.00256f
C14856 _0144_ _0142_ 0
C14857 _0324_ _0689_/a_68_297# 0.00337f
C14858 _0294_ _0583_/a_373_47# 0
C14859 clknet_1_0__leaf__0463_ _0136_ 0.00421f
C14860 _0574_/a_27_297# _1024_/a_1059_315# 0
C14861 _1050_/a_1017_47# _0194_ 0
C14862 _0174_ B[9] 0
C14863 _0366_ _0347_ 0
C14864 VPWR net142 0.33497f
C14865 _1036_/a_1059_315# net26 0.01788f
C14866 hold31/a_391_47# clkbuf_1_1__f__0458_/a_110_47# 0.00116f
C14867 _0743_/a_51_297# _0743_/a_512_297# 0.0116f
C14868 control0.count\[3\] _0170_ 0.02809f
C14869 _0177_ clknet_1_1__leaf__0457_ 0.20005f
C14870 _1002_/a_1059_315# _0765_/a_215_47# 0
C14871 _1054_/a_27_47# net11 0.03072f
C14872 _0596_/a_59_75# _0382_ 0
C14873 hold34/a_49_47# A[10] 0.01355f
C14874 hold28/a_285_47# _0530_/a_81_21# 0
C14875 net223 hold40/a_285_47# 0
C14876 _0391_ hold40/a_49_47# 0
C14877 _0571_/a_27_297# _0571_/a_109_47# 0.00393f
C14878 _0662_/a_81_21# _0292_ 0.0031f
C14879 _0399_ _0190_ 0
C14880 _1052_/a_1059_315# net15 0
C14881 _0467_ _0470_ 0.04975f
C14882 control0.sh control0.reset 0.22441f
C14883 _0428_ _0088_ 0.17558f
C14884 _0999_/a_466_413# _0218_ 0.03049f
C14885 _1012_/a_1017_47# net239 0
C14886 _1054_/a_891_413# _0252_ 0
C14887 _0856_/a_297_297# acc0.A\[1\] 0
C14888 VPWR _0320_ 0.64375f
C14889 clknet_1_0__leaf__0464_ _1049_/a_1059_315# 0.0018f
C14890 hold41/a_285_47# A[10] 0
C14891 clknet_0__0465_ _0825_/a_68_297# 0.00143f
C14892 clkbuf_0__0463_/a_110_47# net7 0
C14893 _0734_/a_47_47# clknet_0__0460_ 0
C14894 _1058_/a_466_413# acc0.A\[11\] 0
C14895 hold100/a_49_47# _0181_ 0
C14896 net150 hold3/a_285_47# 0.0087f
C14897 input2/a_75_212# _0510_/a_109_297# 0
C14898 VPWR _1035_/a_634_159# 0.18467f
C14899 _1053_/a_1059_315# _1052_/a_1059_315# 0
C14900 _1001_/a_27_47# net45 0
C14901 _0504_/a_27_47# _0465_ 0.01721f
C14902 hold22/a_391_47# _0437_ 0
C14903 _0404_ _0345_ 0.03035f
C14904 _0224_ hold4/a_391_47# 0
C14905 _0754_/a_51_297# net241 0.09221f
C14906 _0754_/a_149_47# _0345_ 0.00167f
C14907 _0754_/a_245_297# _0377_ 0.00192f
C14908 _0982_/a_193_47# _0181_ 0.49714f
C14909 _0179_ _1053_/a_193_47# 0
C14910 _0236_ _0764_/a_81_21# 0
C14911 _0992_/a_27_47# _0286_ 0
C14912 _0992_/a_193_47# _0283_ 0
C14913 _0470_ comp0.B\[0\] 0.01911f
C14914 _1056_/a_1059_315# output66/a_27_47# 0
C14915 hold37/a_391_47# _0142_ 0.00171f
C14916 acc0.A\[21\] hold73/a_285_47# 0
C14917 _0266_ _0346_ 0.01918f
C14918 _0187_ _0186_ 0.02417f
C14919 _0504_/a_27_47# acc0.A\[2\] 0
C14920 _0183_ _0487_ 0
C14921 clknet_1_0__leaf__0465_ _0138_ 0
C14922 _1064_/a_27_47# _1064_/a_634_159# 0.13601f
C14923 _0456_ _0465_ 0.00344f
C14924 _0837_/a_81_21# _0256_ 0
C14925 _0350_ net90 0
C14926 _0097_ _0347_ 0.02408f
C14927 clknet_1_1__leaf__0459_ _0786_/a_80_21# 0.00376f
C14928 clk _1068_/a_634_159# 0
C14929 clkbuf_0_clk/a_110_47# _1068_/a_891_413# 0
C14930 _1018_/a_193_47# _1017_/a_27_47# 0
C14931 _1018_/a_27_47# _1017_/a_193_47# 0
C14932 clknet_0__0457_ hold71/a_391_47# 0
C14933 _0837_/a_81_21# _0987_/a_1059_315# 0.00697f
C14934 _1038_/a_1059_315# _0207_ 0.02449f
C14935 _1038_/a_891_413# net171 0.00215f
C14936 _0304_ _0296_ 0
C14937 _0769_/a_81_21# _0771_/a_27_413# 0
C14938 VPWR _0818_/a_193_47# 0
C14939 _0587_/a_27_47# hold92/a_285_47# 0
C14940 _0829_/a_27_47# _0434_ 0
C14941 _0990_/a_27_47# _0988_/a_1059_315# 0
C14942 _1051_/a_193_47# net148 0
C14943 net1 _1063_/a_193_47# 0
C14944 _0454_ net222 0
C14945 _0231_ _0460_ 0
C14946 _1033_/a_193_47# comp0.B\[0\] 0.02493f
C14947 _1053_/a_561_413# net12 0
C14948 _0535_/a_150_297# hold6/a_49_47# 0
C14949 VPWR _0994_/a_561_413# 0.00292f
C14950 _0343_ _1060_/a_1059_315# 0.00368f
C14951 _0324_ net112 0
C14952 net159 _1068_/a_466_413# 0
C14953 control0.state\[0\] _0970_/a_27_297# 0.00827f
C14954 _0490_ clknet_0_clk 0.00874f
C14955 net1 _0460_ 0.03766f
C14956 hold19/a_49_47# clknet_1_1__leaf__0461_ 0
C14957 _0226_ _0183_ 0
C14958 clknet_0__0465_ _0841_/a_79_21# 0.00248f
C14959 clknet_1_0__leaf__0458_ _0854_/a_297_297# 0
C14960 _1028_/a_27_47# net156 0
C14961 hold5/a_285_47# net20 0
C14962 _0461_ _1015_/a_561_413# 0
C14963 _0324_ acc0.A\[24\] 0.36194f
C14964 net62 _0181_ 0.00402f
C14965 _0553_/a_51_297# _0209_ 0.10887f
C14966 net157 control0.reset 0
C14967 _0118_ clknet_1_0__leaf__0459_ 0.03265f
C14968 _1010_/a_891_413# _0350_ 0.06108f
C14969 _0576_/a_27_297# net50 0.00199f
C14970 _0477_ _0951_/a_209_311# 0.00914f
C14971 _0181_ _0450_ 0
C14972 hold13/a_391_47# _1034_/a_1059_315# 0
C14973 hold13/a_285_47# _1034_/a_891_413# 0
C14974 _0259_ _0990_/a_634_159# 0
C14975 net101 _0345_ 0.0014f
C14976 _0338_ net209 0
C14977 _0222_ _1005_/a_975_413# 0
C14978 _0180_ _0449_ 0
C14979 _0195_ _0244_ 0
C14980 _0565_/a_512_297# _0173_ 0
C14981 _0287_ _0809_/a_384_47# 0
C14982 net61 _0274_ 0.03551f
C14983 net157 _1061_/a_891_413# 0.02016f
C14984 _0846_/a_149_47# _0350_ 0.00143f
C14985 hold70/a_49_47# net37 0.28377f
C14986 _0544_/a_51_297# _0543_/a_68_297# 0
C14987 _0800_/a_51_297# _0997_/a_27_47# 0
C14988 VPWR _0720_/a_68_297# 0.16924f
C14989 _1056_/a_27_47# _0988_/a_1059_315# 0
C14990 _0995_/a_891_413# _0219_ 0
C14991 _0227_ _0618_/a_297_297# 0
C14992 _0457_ net1 0.2366f
C14993 net230 _0179_ 0.17086f
C14994 _0695_/a_300_47# _0312_ 0
C14995 _0695_/a_217_297# _0323_ 0.01218f
C14996 _0180_ _0498_/a_149_47# 0
C14997 net247 hold71/a_285_47# 0.04002f
C14998 net138 _1053_/a_27_47# 0
C14999 _0183_ _1016_/a_193_47# 0
C15000 net108 _0183_ 0
C15001 clknet_1_0__leaf__0462_ _0120_ 0.04331f
C15002 _1031_/a_634_159# _1031_/a_592_47# 0
C15003 _0531_/a_109_297# _1047_/a_466_413# 0
C15004 net45 _0459_ 1.1782f
C15005 comp0.B\[14\] _0141_ 0
C15006 net68 clkbuf_1_1__f__0457_/a_110_47# 0.00594f
C15007 net67 hold70/a_391_47# 0.04588f
C15008 hold30/a_49_47# _0756_/a_285_47# 0
C15009 input2/a_75_212# _0188_ 0
C15010 _1041_/a_634_159# VPWR 0.18276f
C15011 acc0.A\[7\] _0829_/a_27_47# 0
C15012 net31 _0139_ 0
C15013 _0415_ _0403_ 0.32848f
C15014 _1022_/a_27_47# _1005_/a_27_47# 0
C15015 _0316_ _0689_/a_68_297# 0
C15016 _0369_ clkbuf_0__0459_/a_110_47# 0.01599f
C15017 pp[15] _0995_/a_193_47# 0.00605f
C15018 _1005_/a_381_47# net91 0
C15019 _1005_/a_891_413# _0103_ 0.0554f
C15020 _0388_ _0247_ 0
C15021 net213 net49 0
C15022 _0325_ _0315_ 0
C15023 _1060_/a_466_413# net5 0
C15024 _1060_/a_193_47# _0185_ 0.0011f
C15025 _0191_ A[8] 0
C15026 _0976_/a_505_21# _1069_/a_1059_315# 0
C15027 _1054_/a_27_47# clknet_1_1__leaf__0458_ 0
C15028 net1 _1062_/a_891_413# 0
C15029 _1002_/a_634_159# _1002_/a_1017_47# 0
C15030 _1002_/a_466_413# _1002_/a_592_47# 0.00553f
C15031 clkbuf_1_0__f__0458_/a_110_47# _0350_ 0.19044f
C15032 _1027_/a_193_47# _0365_ 0
C15033 _0183_ clkbuf_0__0457_/a_110_47# 0.02693f
C15034 _0640_/a_465_297# VPWR 0
C15035 net29 _1040_/a_1059_315# 0
C15036 _0984_/a_975_413# clknet_1_0__leaf__0458_ 0.00107f
C15037 _0623_/a_109_297# _0440_ 0
C15038 _0820_/a_79_21# _0820_/a_297_297# 0.01735f
C15039 _0174_ _1041_/a_1017_47# 0
C15040 _0965_/a_47_47# control0.count\[0\] 0
C15041 _0340_ _0704_/a_68_297# 0
C15042 _0710_/a_109_297# acc0.A\[30\] 0
C15043 _1028_/a_27_47# acc0.A\[26\] 0
C15044 _0154_ _1055_/a_1059_315# 0
C15045 VPWR _0997_/a_975_413# 0.00418f
C15046 _0409_ _0400_ 0
C15047 acc0.A\[12\] _0422_ 0.00231f
C15048 _0662_/a_299_297# _0785_/a_81_21# 0
C15049 _0713_/a_27_47# _0346_ 0.00305f
C15050 _0217_ _1019_/a_592_47# 0
C15051 net203 net186 0
C15052 _0362_ _0361_ 0.00869f
C15053 net54 hold8/a_285_47# 0.01222f
C15054 _1041_/a_193_47# _0550_/a_51_297# 0
C15055 hold77/a_285_47# _0327_ 0
C15056 _0664_/a_297_47# clknet_1_1__leaf__0459_ 0
C15057 _1035_/a_561_413# _0175_ 0
C15058 _0765_/a_510_47# _0385_ 0.00331f
C15059 _0305_ net219 0
C15060 _0372_ net216 0
C15061 pp[28] _1011_/a_1059_315# 0
C15062 VPWR _1061_/a_1017_47# 0
C15063 output66/a_27_47# VPWR 0.33769f
C15064 clknet_1_0__leaf__0463_ _1046_/a_381_47# 0
C15065 _0343_ net93 0.04676f
C15066 control0.count\[1\] _0977_/a_75_212# 0
C15067 _0168_ _0489_ 0.00705f
C15068 _0399_ _0306_ 0.00135f
C15069 VPWR _0668_/a_297_47# 0.00543f
C15070 _1034_/a_891_413# _0132_ 0
C15071 net103 _0675_/a_68_297# 0
C15072 _0971_/a_384_47# _0487_ 0
C15073 _1036_/a_27_47# input24/a_75_212# 0
C15074 control0.state\[1\] net240 0.00143f
C15075 _1035_/a_975_413# control0.sh 0
C15076 _0176_ clknet_1_1__leaf__0464_ 0.24919f
C15077 _0176_ _0548_/a_149_47# 0.00414f
C15078 _1000_/a_193_47# _0393_ 0.01724f
C15079 clknet_1_0__leaf__0465_ net134 0.00517f
C15080 clknet_1_0__leaf__0458_ _0198_ 0
C15081 _0343_ _0796_/a_510_47# 0.00105f
C15082 comp0.B\[12\] _1044_/a_27_47# 0
C15083 _0811_/a_384_47# _0296_ 0
C15084 control0.state\[2\] _0484_ 0.00168f
C15085 control0.count\[1\] _1069_/a_975_413# 0.00112f
C15086 VPWR clknet_1_0__leaf_clk 3.95529f
C15087 _0985_/a_891_413# _0218_ 0
C15088 hold39/a_49_47# clknet_1_1__leaf__0463_ 0.00407f
C15089 net53 _0123_ 0.07093f
C15090 _1018_/a_1059_315# _0218_ 0
C15091 _1030_/a_1059_315# _0220_ 0.02401f
C15092 _1030_/a_466_413# _0336_ 0
C15093 _0414_ _0994_/a_27_47# 0.00395f
C15094 _0695_/a_217_297# net237 0
C15095 _0323_ _0743_/a_149_47# 0
C15096 hold30/a_285_47# net110 0
C15097 _0172_ hold1/a_49_47# 0
C15098 _0369_ _1005_/a_466_413# 0
C15099 _1011_/a_975_413# net57 0
C15100 _1017_/a_193_47# clknet_1_1__leaf__0461_ 0
C15101 _0572_/a_27_297# _0572_/a_373_47# 0.01338f
C15102 _0107_ _0322_ 0.00116f
C15103 _0216_ _1006_/a_27_47# 0.03051f
C15104 _0343_ _0294_ 0.11772f
C15105 _1006_/a_891_413# _1006_/a_1017_47# 0.00617f
C15106 _0179_ _0987_/a_381_47# 0.00114f
C15107 _1006_/a_634_159# net92 0
C15108 _0698_/a_113_297# _0324_ 0
C15109 _0656_/a_59_75# _0288_ 0.11218f
C15110 VPWR net116 0.45558f
C15111 _0107_ _0327_ 0
C15112 _0993_/a_891_413# net246 0.00229f
C15113 output65/a_27_47# _0369_ 0.00199f
C15114 _0221_ _0353_ 0.16882f
C15115 _0323_ _0345_ 0
C15116 clknet_1_0__leaf__0460_ _0754_/a_240_47# 0
C15117 _0984_/a_634_159# _0984_/a_1017_47# 0
C15118 _0984_/a_466_413# _0984_/a_592_47# 0.00553f
C15119 hold10/a_285_47# _0172_ 0
C15120 net180 _1061_/a_27_47# 0
C15121 _0294_ net95 0
C15122 _0347_ net112 0
C15123 net155 acc0.A\[25\] 0
C15124 _0808_/a_266_47# _0419_ 0.06468f
C15125 _0808_/a_266_297# _0091_ 0
C15126 _0439_ _0988_/a_27_47# 0.00755f
C15127 _0438_ _0988_/a_466_413# 0
C15128 clkload0/X _0466_ 0
C15129 _0347_ acc0.A\[24\] 0.33349f
C15130 VPWR _0988_/a_27_47# 0.63415f
C15131 _0514_/a_27_297# acc0.A\[10\] 0.06205f
C15132 hold97/a_285_47# _0106_ 0.00304f
C15133 _0982_/a_1059_315# net165 0
C15134 comp0.B\[6\] hold84/a_391_47# 0
C15135 _1039_/a_1017_47# VPWR 0
C15136 _0285_ hold81/a_49_47# 0
C15137 hold78/a_49_47# _1031_/a_1059_315# 0
C15138 _0730_/a_215_47# VPWR 0.00228f
C15139 _0404_ _0791_/a_113_297# 0
C15140 _0986_/a_891_413# _0986_/a_1017_47# 0.00617f
C15141 net168 _1054_/a_634_159# 0.00219f
C15142 _1056_/a_193_47# _0186_ 0.03246f
C15143 clknet_1_1__leaf_clk clknet_1_0__leaf__0461_ 0.00302f
C15144 VPWR hold92/a_285_47# 0.31974f
C15145 _0118_ _0113_ 0
C15146 hold43/a_391_47# acc0.A\[29\] 0
C15147 _1023_/a_891_413# net109 0
C15148 _1023_/a_1059_315# net177 0
C15149 _1023_/a_193_47# acc0.A\[23\] 0
C15150 _0990_/a_381_47# net47 0.00611f
C15151 _1037_/a_1059_315# _0175_ 0.00112f
C15152 net45 _0220_ 0.00113f
C15153 _0369_ _1006_/a_193_47# 0
C15154 _0512_/a_109_297# acc0.A\[10\] 0
C15155 hold32/a_285_47# A[10] 0
C15156 _0094_ _0507_/a_109_297# 0
C15157 _0753_/a_381_47# _0227_ 0
C15158 clkbuf_1_0__f__0459_/a_110_47# net47 0
C15159 _0697_/a_80_21# _0686_/a_27_53# 0
C15160 _0572_/a_27_297# acc0.A\[27\] 0
C15161 net155 _0571_/a_27_297# 0.07104f
C15162 _0195_ _0571_/a_109_297# 0.01782f
C15163 _0135_ _0209_ 0
C15164 hold58/a_391_47# clknet_1_1__leaf__0463_ 0.01846f
C15165 hold58/a_49_47# net122 0
C15166 net34 _0946_/a_184_297# 0.00401f
C15167 clknet_1_1__leaf__0464_ net130 0.2157f
C15168 _0691_/a_150_297# _0359_ 0
C15169 _0691_/a_68_297# _0324_ 0
C15170 _1011_/a_193_47# _0339_ 0
C15171 _0538_/a_51_297# _0172_ 0.14335f
C15172 _0982_/a_1059_315# acc0.A\[19\] 0
C15173 net36 pp[0] 0.00831f
C15174 _1045_/a_1017_47# net20 0
C15175 _1037_/a_891_413# control0.sh 0.00641f
C15176 net150 _0721_/a_27_47# 0
C15177 net234 clknet_1_0__leaf__0461_ 0
C15178 hold55/a_391_47# _0181_ 0.02775f
C15179 _0179_ acc0.A\[4\] 0.02163f
C15180 net141 pp[4] 0
C15181 net158 net184 0
C15182 _1001_/a_27_47# VPWR 0.56295f
C15183 clknet_1_0__leaf__0464_ net175 0
C15184 hold36/a_285_47# clkbuf_0__0464_/a_110_47# 0.02007f
C15185 _0183_ _0534_/a_299_297# 0
C15186 _0129_ _1031_/a_1059_315# 0
C15187 net163 _1031_/a_634_159# 0
C15188 _0988_/a_27_47# output62/a_27_47# 0
C15189 acc0.A\[16\] _0781_/a_68_297# 0.01567f
C15190 _0340_ _0216_ 0.23869f
C15191 _0128_ hold61/a_285_47# 0.01038f
C15192 _0616_/a_493_297# _0616_/a_215_47# 0
C15193 _1059_/a_1059_315# net229 0
C15194 _0419_ _0345_ 0.08081f
C15195 hold22/a_391_47# _0252_ 0
C15196 net46 clknet_1_0__leaf__0461_ 0.00166f
C15197 _0578_/a_109_297# _1067_/a_1059_315# 0
C15198 net165 _0451_ 0.03285f
C15199 hold42/a_391_47# _0156_ 0
C15200 _0375_ net51 0.04043f
C15201 _1057_/a_891_413# _0156_ 0.00145f
C15202 _1038_/a_1059_315# _1037_/a_1059_315# 0
C15203 net187 _0369_ 0
C15204 _0257_ _0835_/a_215_47# 0.07068f
C15205 _0626_/a_68_297# _0255_ 0
C15206 pp[15] _0093_ 0.0036f
C15207 clknet_0__0457_ net187 0.452f
C15208 VPWR hold8/a_49_47# 0.30827f
C15209 clkbuf_0__0457_/a_110_47# hold40/a_285_47# 0
C15210 net44 _0588_/a_113_47# 0
C15211 net182 net142 0.00928f
C15212 _0225_ _0460_ 0.0022f
C15213 _0997_/a_1059_315# _0095_ 0
C15214 _0556_/a_150_297# clknet_1_1__leaf__0463_ 0
C15215 comp0.B\[5\] _0549_/a_68_297# 0.0027f
C15216 hold99/a_391_47# net246 0.1316f
C15217 _0852_/a_285_47# _0264_ 0.00212f
C15218 hold24/a_391_47# _0176_ 0
C15219 _0776_/a_109_297# _0776_/a_27_47# 0
C15220 _0216_ _0737_/a_35_297# 0
C15221 _0238_ control0.add 0
C15222 _0607_/a_27_297# _0310_ 0
C15223 _0743_/a_149_47# net237 0.00107f
C15224 _0729_/a_68_297# acc0.A\[29\] 0.00199f
C15225 _1053_/a_193_47# hold83/a_49_47# 0.00957f
C15226 _1053_/a_27_47# hold83/a_285_47# 0
C15227 _0770_/a_297_47# _0719_/a_27_47# 0
C15228 _0579_/a_109_297# _0346_ 0.00292f
C15229 net57 _0334_ 0.82978f
C15230 acc0.A\[15\] net41 0.09544f
C15231 _1065_/a_27_47# _1065_/a_1059_315# 0.04875f
C15232 _1065_/a_193_47# _1065_/a_466_413# 0.07482f
C15233 _0395_ _0308_ 0.00196f
C15234 _0217_ _0760_/a_129_47# 0.00139f
C15235 net150 _0760_/a_285_47# 0
C15236 _0183_ _0760_/a_47_47# 0.00629f
C15237 net232 _1066_/a_466_413# 0
C15238 hold30/a_391_47# _0120_ 0.00906f
C15239 _0121_ acc0.A\[22\] 0.00107f
C15240 _0787_/a_209_47# _0281_ 0.00139f
C15241 _0787_/a_80_21# _0418_ 0
C15242 _0587_/a_27_47# _0220_ 0.01075f
C15243 _0998_/a_27_47# _0218_ 0.03548f
C15244 _1036_/a_193_47# _1035_/a_193_47# 0
C15245 _1036_/a_634_159# _1035_/a_27_47# 0.00294f
C15246 _0532_/a_299_297# _0198_ 0.01146f
C15247 A[4] input15/a_75_212# 0.00986f
C15248 input11/a_75_212# A[8] 0.00126f
C15249 net202 _1067_/a_1059_315# 0
C15250 _0601_/a_68_297# acc0.A\[23\] 0.17826f
C15251 _0216_ _0722_/a_297_297# 0
C15252 _0985_/a_27_47# _0270_ 0
C15253 _0707_/a_75_199# _0707_/a_201_297# 0.15956f
C15254 hold79/a_49_47# _1070_/a_27_47# 0
C15255 _1057_/a_381_47# _0992_/a_1059_315# 0
C15256 _0399_ _0346_ 0.2867f
C15257 net237 _0345_ 0.10516f
C15258 _0954_/a_114_297# _1042_/a_193_47# 0
C15259 _0954_/a_220_297# _1042_/a_27_47# 0
C15260 _0305_ _0352_ 0.02938f
C15261 clknet_1_1__leaf__0463_ _1067_/a_1059_315# 0.01136f
C15262 net152 _0540_/a_51_297# 0
C15263 _0508_/a_81_21# hold82/a_285_47# 0
C15264 VPWR _1047_/a_193_47# 0.30872f
C15265 _0811_/a_81_21# _0811_/a_384_47# 0.00138f
C15266 hold17/a_285_47# clknet_1_0__leaf_clk 0.00196f
C15267 _0627_/a_215_53# clknet_0__0465_ 0.01071f
C15268 _0349_ _0352_ 0.43976f
C15269 VPWR _0957_/a_304_297# 0.00455f
C15270 _0236_ _0372_ 0.02064f
C15271 _0181_ net219 0
C15272 _0373_ _0374_ 0.04725f
C15273 _0332_ hold95/a_391_47# 0
C15274 hold101/a_49_47# hold101/a_391_47# 0.00188f
C15275 _0985_/a_27_47# _0858_/a_27_47# 0
C15276 _0399_ net65 0.17804f
C15277 hold57/a_285_47# net8 0
C15278 control0.count\[3\] net35 0.20818f
C15279 VPWR _1007_/a_1059_315# 0.37608f
C15280 _0399_ _0989_/a_466_413# 0.00461f
C15281 VPWR net121 0.57989f
C15282 _0260_ _0180_ 0
C15283 _0172_ _1040_/a_381_47# 0.00787f
C15284 _0710_/a_381_47# _0339_ 0
C15285 _0966_/a_109_297# _0170_ 0
C15286 _1058_/a_381_47# VPWR 0.07542f
C15287 _0179_ _1051_/a_466_413# 0.00401f
C15288 _0403_ _0347_ 0.20418f
C15289 net241 _0219_ 0.12028f
C15290 _0534_/a_299_297# acc0.A\[15\] 0
C15291 VPWR _0420_ 0.22206f
C15292 _0178_ _1049_/a_193_47# 0
C15293 output56/a_27_47# _0704_/a_68_297# 0
C15294 _1055_/a_27_47# net16 0.00625f
C15295 _1064_/a_891_413# _1064_/a_975_413# 0.00851f
C15296 _1064_/a_381_47# _1064_/a_561_413# 0.00123f
C15297 _0316_ _0698_/a_113_297# 0.01401f
C15298 clk clknet_1_1__leaf_clk 0
C15299 acc0.A\[27\] _0360_ 0
C15300 _0274_ _0431_ 0.06572f
C15301 hold78/a_391_47# _0345_ 0
C15302 clknet_1_0__leaf__0458_ _0852_/a_285_297# 0.00283f
C15303 pp[27] output56/a_27_47# 0.01289f
C15304 _0442_ _0271_ 0
C15305 hold27/a_285_47# clknet_1_1__leaf__0457_ 0.0012f
C15306 VPWR _0459_ 0.93991f
C15307 _0669_/a_29_53# _0669_/a_111_297# 0.005f
C15308 control0.add _0721_/a_27_47# 0
C15309 clknet_1_1__leaf_clk _1063_/a_891_413# 0
C15310 net112 _1025_/a_27_47# 0.01102f
C15311 _1002_/a_27_47# _1067_/a_1059_315# 0
C15312 VPWR hold80/a_285_47# 0.28636f
C15313 _0260_ _0432_ 0
C15314 clkbuf_1_0__f__0459_/a_110_47# _1060_/a_1059_315# 0.01627f
C15315 _0959_/a_217_297# clknet_1_1__leaf_clk 0
C15316 _0343_ _1017_/a_561_413# 0
C15317 _1002_/a_891_413# _0369_ 0.0024f
C15318 _0234_ acc0.A\[21\] 0
C15319 _0192_ hold83/a_285_47# 0
C15320 net230 hold83/a_49_47# 0
C15321 _1025_/a_27_47# acc0.A\[24\] 0
C15322 _0438_ _0186_ 0.12916f
C15323 clknet_1_0__leaf__0462_ _0753_/a_79_21# 0
C15324 _0385_ _0384_ 0
C15325 _0130_ comp0.B\[0\] 0
C15326 net14 VPWR 0.67527f
C15327 net159 _0166_ 0
C15328 net34 _0967_/a_297_297# 0
C15329 control0.state\[1\] _0967_/a_403_297# 0
C15330 control0.state\[0\] _0967_/a_487_297# 0.00112f
C15331 net34 _0162_ 0.14879f
C15332 _0257_ _0172_ 0
C15333 hold65/a_285_47# net63 0
C15334 _0985_/a_634_159# net61 0
C15335 _0985_/a_27_47# net233 0
C15336 _1013_/a_634_159# _0339_ 0
C15337 _0323_ net52 0
C15338 _0636_/a_59_75# _0186_ 0.00472f
C15339 hold24/a_49_47# clkbuf_1_0__f__0463_/a_110_47# 0.02055f
C15340 _1017_/a_381_47# acc0.A\[17\] 0
C15341 _0404_ _0994_/a_27_47# 0
C15342 _0352_ hold73/a_49_47# 0.00605f
C15343 _1008_/a_891_413# _0345_ 0
C15344 _0360_ _0364_ 0.02477f
C15345 clknet_1_0__leaf__0458_ net247 0.07278f
C15346 hold13/a_49_47# comp0.B\[2\] 0
C15347 _0222_ _1022_/a_27_47# 0.01486f
C15348 _0118_ _0579_/a_373_47# 0
C15349 net163 _0345_ 0
C15350 _0854_/a_215_47# _0454_ 0.05456f
C15351 _0963_/a_285_297# _1070_/a_891_413# 0
C15352 _1017_/a_1059_315# clkbuf_1_1__f__0461_/a_110_47# 0
C15353 _0313_ _1026_/a_193_47# 0
C15354 hold74/a_391_47# _1016_/a_1059_315# 0.01554f
C15355 _0316_ _0691_/a_68_297# 0
C15356 _0479_ clk 0
C15357 _0346_ _0808_/a_266_297# 0.00103f
C15358 _0322_ _0327_ 0.02979f
C15359 _0413_ _0997_/a_634_159# 0
C15360 hold28/a_49_47# net175 0.03328f
C15361 hold36/a_391_47# _0143_ 0.04931f
C15362 _0498_/a_51_297# _0498_/a_149_47# 0.02487f
C15363 _0830_/a_215_47# _0437_ 0.01383f
C15364 _0830_/a_79_21# _0087_ 0.05048f
C15365 _0830_/a_510_47# net212 0.00259f
C15366 _0246_ _0242_ 0
C15367 _0841_/a_79_21# _0986_/a_27_47# 0.00136f
C15368 clknet_1_1__leaf__0460_ _1028_/a_27_47# 0
C15369 _0179_ net217 0.03047f
C15370 _0313_ hold97/a_49_47# 0.00178f
C15371 _1015_/a_1059_315# clknet_1_0__leaf__0461_ 0.00908f
C15372 net1 _0958_/a_303_47# 0.00187f
C15373 clknet_1_0__leaf__0465_ _1052_/a_975_413# 0
C15374 net8 _0159_ 0.00105f
C15375 _1034_/a_27_47# _0131_ 0
C15376 _1034_/a_193_47# net119 0
C15377 _0409_ clkbuf_0__0459_/a_110_47# 0
C15378 _0179_ A[11] 0
C15379 _1037_/a_1017_47# VPWR 0
C15380 _0557_/a_245_297# _0557_/a_240_47# 0
C15381 _0441_ acc0.A\[4\] 0
C15382 _0217_ net166 0
C15383 _0332_ acc0.A\[28\] 0.008f
C15384 _0596_/a_59_75# net91 0.02418f
C15385 _0514_/a_109_297# _0181_ 0.05782f
C15386 _0289_ _0402_ 0.14426f
C15387 _0195_ _1014_/a_27_47# 0
C15388 _0255_ _0252_ 0.00176f
C15389 A[13] input6/a_75_212# 0.01105f
C15390 _0180_ _0524_/a_27_297# 0.10225f
C15391 VPWR _0265_ 0.45708f
C15392 VPWR clkbuf_1_0__f__0462_/a_110_47# 1.26502f
C15393 _0121_ _0379_ 0
C15394 _0361_ _0324_ 0.23808f
C15395 _0516_/a_109_47# net142 0.00147f
C15396 _0845_/a_109_47# _0844_/a_79_21# 0
C15397 clknet_1_0__leaf__0465_ net22 0.00224f
C15398 clknet_1_0__leaf__0458_ _0844_/a_382_297# 0
C15399 hold51/a_49_47# hold51/a_391_47# 0.00188f
C15400 _0837_/a_81_21# clknet_0__0465_ 0
C15401 net17 net201 0.09203f
C15402 net11 _0523_/a_299_297# 0.01065f
C15403 net26 hold84/a_391_47# 0
C15404 hold7/a_285_47# acc0.A\[6\] 0
C15405 _1001_/a_27_47# clknet_1_0__leaf__0459_ 0
C15406 _0512_/a_109_47# _0181_ 0.00405f
C15407 clknet_1_1__leaf_clk _1062_/a_592_47# 0.00172f
C15408 clknet_1_0__leaf__0465_ net75 0
C15409 _1018_/a_27_47# net219 0.00209f
C15410 _1018_/a_381_47# _0581_/a_27_297# 0
C15411 _0158_ net5 0.0014f
C15412 input31/a_75_212# input7/a_75_212# 0.01252f
C15413 _0482_ _0486_ 0
C15414 _1008_/a_27_47# _1008_/a_466_413# 0.27314f
C15415 _1008_/a_193_47# _1008_/a_634_159# 0.11072f
C15416 _0488_ _1069_/a_891_413# 0
C15417 _0466_ _1069_/a_1059_315# 0
C15418 _0249_ _0373_ 0
C15419 _1021_/a_561_413# clknet_1_1__leaf_clk 0
C15420 _0179_ _0744_/a_27_47# 0.00359f
C15421 hold16/a_49_47# net163 0
C15422 hold16/a_391_47# _0129_ 0
C15423 pp[27] _0707_/a_315_47# 0
C15424 _0718_/a_47_47# _1011_/a_193_47# 0
C15425 _1041_/a_1017_47# comp0.B\[9\] 0
C15426 _1002_/a_592_47# _0100_ 0.00164f
C15427 _1020_/a_634_159# _1020_/a_975_413# 0
C15428 _1020_/a_466_413# _1020_/a_561_413# 0.00772f
C15429 net40 _0278_ 0.04704f
C15430 hold76/a_49_47# net211 0
C15431 output53/a_27_47# _1025_/a_27_47# 0
C15432 _0405_ _0406_ 0.11112f
C15433 _0390_ _0459_ 0
C15434 _1035_/a_634_159# comp0.B\[3\] 0
C15435 _1035_/a_27_47# comp0.B\[5\] 0
C15436 _0559_/a_51_297# _0561_/a_51_297# 0
C15437 _1003_/a_27_47# hold12/a_49_47# 0.00154f
C15438 _0564_/a_150_297# _0173_ 0
C15439 _0119_ net1 0
C15440 A[11] _0513_/a_81_21# 0
C15441 clkbuf_1_0__f__0464_/a_110_47# _1049_/a_1059_315# 0.01266f
C15442 _0239_ _0607_/a_27_297# 0.10985f
C15443 _0107_ _0346_ 0
C15444 _0226_ _0752_/a_27_413# 0
C15445 _0598_/a_79_21# _0375_ 0
C15446 _0598_/a_297_47# _0234_ 0
C15447 output59/a_27_47# net57 0
C15448 B[10] net10 0.03456f
C15449 clknet_1_0__leaf__0463_ clknet_1_0__leaf__0465_ 0.03323f
C15450 hold28/a_285_47# _0147_ 0.03534f
C15451 hold28/a_391_47# net135 0
C15452 _0983_/a_975_413# net47 0.0025f
C15453 acc0.A\[22\] _0380_ 0
C15454 _0515_/a_81_21# _0515_/a_384_47# 0.00138f
C15455 _0183_ _0350_ 0.07633f
C15456 pp[8] input16/a_75_212# 0.02104f
C15457 _0559_/a_240_47# _0957_/a_32_297# 0.00157f
C15458 _0472_ _0175_ 0.05757f
C15459 _0343_ _0606_/a_215_297# 0
C15460 _1031_/a_1059_315# hold61/a_285_47# 0
C15461 _0188_ _0512_/a_109_297# 0.00169f
C15462 _0346_ _0295_ 0.05694f
C15463 _0180_ _1048_/a_975_413# 0
C15464 _0199_ _1048_/a_891_413# 0
C15465 _0411_ _0300_ 0.00165f
C15466 hold69/a_285_47# _0328_ 0
C15467 clknet_0__0458_ _0264_ 0
C15468 _1013_/a_466_413# net99 0
C15469 _1001_/a_1017_47# net46 0.00187f
C15470 _0457_ net157 0
C15471 _0314_ _0366_ 0.13222f
C15472 _1041_/a_193_47# _0172_ 0.04531f
C15473 _1041_/a_634_159# net30 0
C15474 _0559_/a_51_297# _0133_ 0.10182f
C15475 _0181_ _0352_ 0.02458f
C15476 _1039_/a_381_47# _0494_/a_27_47# 0
C15477 pp[12] A[14] 0
C15478 net227 hold80/a_391_47# 0.1316f
C15479 _0992_/a_193_47# _0345_ 0
C15480 hold7/a_391_47# _0523_/a_299_297# 0
C15481 output56/a_27_47# _0216_ 0.00508f
C15482 _0570_/a_27_297# _0739_/a_79_21# 0
C15483 _0645_/a_129_47# net41 0.00236f
C15484 net111 _0347_ 0
C15485 _0284_ VPWR 0.86567f
C15486 clkbuf_1_1__f__0457_/a_110_47# hold71/a_49_47# 0
C15487 _0475_ control0.sh 0
C15488 net57 _0724_/a_113_297# 0.06909f
C15489 hold21/a_285_47# input15/a_75_212# 0.00429f
C15490 hold94/a_391_47# _0754_/a_149_47# 0
C15491 hold94/a_285_47# _0754_/a_240_47# 0
C15492 _0991_/a_27_47# acc0.A\[15\] 0.00123f
C15493 _0826_/a_27_53# _0826_/a_301_297# 0
C15494 _0440_ _1051_/a_1059_315# 0
C15495 clknet_0__0459_ _0796_/a_79_21# 0.00555f
C15496 clknet_1_0__leaf__0462_ _0752_/a_384_47# 0
C15497 _0197_ _0270_ 0
C15498 hold63/a_49_47# net53 0
C15499 _0990_/a_193_47# net62 0.01434f
C15500 _1072_/a_1059_315# _0468_ 0
C15501 clknet_1_0__leaf__0465_ net138 0.182f
C15502 hold42/a_285_47# _1058_/a_27_47# 0
C15503 _0172_ net11 0.026f
C15504 _1058_/a_466_413# _1057_/a_193_47# 0
C15505 _1058_/a_1059_315# _1057_/a_27_47# 0
C15506 _1058_/a_27_47# _1057_/a_1059_315# 0
C15507 _1058_/a_193_47# _1057_/a_466_413# 0
C15508 _1058_/a_634_159# _1057_/a_634_159# 0
C15509 VPWR _0220_ 0.80404f
C15510 _0273_ _0641_/a_113_47# 0.00937f
C15511 _0458_ _0530_/a_81_21# 0
C15512 _0464_ _0465_ 0.0263f
C15513 clknet_1_1__leaf__0465_ _0186_ 0.42433f
C15514 clknet_1_0__leaf__0458_ net100 0
C15515 B[9] hold5/a_285_47# 0.00389f
C15516 _1056_/a_975_413# VPWR 0.00464f
C15517 _0427_ _0345_ 0
C15518 _0662_/a_81_21# clkbuf_1_1__f__0465_/a_110_47# 0
C15519 _0159_ net10 0
C15520 _1000_/a_381_47# _0347_ 0.01536f
C15521 _1000_/a_466_413# _0352_ 0.02829f
C15522 VPWR _1063_/a_381_47# 0.07064f
C15523 _0996_/a_193_47# _1060_/a_1059_315# 0
C15524 _0284_ _0654_/a_27_413# 0.24989f
C15525 _0285_ _0654_/a_207_413# 0.19076f
C15526 _0369_ _0103_ 0
C15527 net86 _0246_ 0
C15528 net210 net155 0.00321f
C15529 _0572_/a_373_47# _0124_ 0
C15530 acc0.A\[14\] net5 0.02437f
C15531 VPWR _0959_/a_472_297# 0.00413f
C15532 hold36/a_49_47# _0473_ 0
C15533 clknet_1_0__leaf__0459_ _0459_ 0.24218f
C15534 VPWR _0585_/a_109_297# 0.17878f
C15535 _0697_/a_80_21# _0320_ 0.0015f
C15536 comp0.B\[2\] net17 0
C15537 pp[19] output51/a_27_47# 0.00175f
C15538 _0283_ _0420_ 0.18402f
C15539 _0350_ acc0.A\[15\] 0.06708f
C15540 _0856_/a_510_47# _0195_ 0
C15541 _0126_ hold9/a_49_47# 0.04274f
C15542 clknet_1_0__leaf__0462_ _0250_ 0
C15543 _0804_/a_79_21# _0802_/a_59_75# 0.00178f
C15544 _0274_ _0269_ 0.0349f
C15545 _0347_ hold50/a_285_47# 0.02427f
C15546 _1056_/a_193_47# net62 0
C15547 _0984_/a_466_413# net229 0
C15548 clknet_0_clk control0.count\[0\] 0
C15549 VPWR _1060_/a_381_47# 0.07867f
C15550 _0548_/a_51_297# _0548_/a_512_297# 0.0116f
C15551 _1019_/a_1059_315# _0242_ 0
C15552 pp[28] _0707_/a_208_47# 0.0019f
C15553 _0584_/a_27_297# _0208_ 0
C15554 _0385_ _0383_ 0
C15555 hold65/a_49_47# clkbuf_1_0__f__0465_/a_110_47# 0
C15556 _0835_/a_215_47# clknet_1_1__leaf__0458_ 0
C15557 hold84/a_285_47# hold84/a_391_47# 0.41909f
C15558 _0179_ net66 0.44457f
C15559 _0189_ acc0.A\[10\] 0.01851f
C15560 _0985_/a_27_47# hold23/a_49_47# 0.00617f
C15561 _1043_/a_27_47# _0543_/a_68_297# 0
C15562 net10 _0447_ 0
C15563 _0172_ hold7/a_391_47# 0
C15564 _0118_ _0345_ 0.00139f
C15565 net168 net140 0.06327f
C15566 net234 _0218_ 0
C15567 _0402_ _0655_/a_109_93# 0
C15568 _0174_ _1043_/a_381_47# 0.01071f
C15569 clknet_0_clk _0974_/a_544_297# 0.00118f
C15570 _0511_/a_81_21# _0511_/a_299_297# 0.08213f
C15571 _0216_ _0247_ 0.23028f
C15572 hold89/a_285_47# _0486_ 0
C15573 hold89/a_391_47# control0.state\[2\] 0.04689f
C15574 clknet_0_clk clknet_1_0__leaf__0457_ 0
C15575 net65 _0619_/a_68_297# 0.13288f
C15576 _0643_/a_103_199# _0432_ 0
C15577 _0619_/a_68_297# _0989_/a_466_413# 0.00748f
C15578 _0179_ _0991_/a_27_47# 0
C15579 clkbuf_1_0__f__0457_/a_110_47# _0216_ 0
C15580 _0316_ _0361_ 0
C15581 _0704_/a_150_297# acc0.A\[30\] 0.00126f
C15582 _1044_/a_592_47# net20 0
C15583 _0682_/a_68_297# _1025_/a_193_47# 0
C15584 net46 _0218_ 0.06235f
C15585 pp[27] _1010_/a_466_413# 0
C15586 clknet_1_1__leaf__0458_ _0523_/a_299_297# 0
C15587 _0217_ acc0.A\[1\] 0.14327f
C15588 net59 _0110_ 0
C15589 pp[30] _0351_ 0
C15590 comp0.B\[11\] _0139_ 0
C15591 _0326_ _0368_ 0
C15592 hold36/a_49_47# _0186_ 0
C15593 _0404_ _0411_ 0.19856f
C15594 _0124_ acc0.A\[27\] 0
C15595 net155 _0125_ 0
C15596 _0799_/a_80_21# _0219_ 0.0073f
C15597 clknet_1_0__leaf__0465_ _0442_ 0.08649f
C15598 _0457_ _1015_/a_975_413# 0
C15599 _0532_/a_81_21# _1048_/a_1059_315# 0.00186f
C15600 _0402_ _0418_ 0.2836f
C15601 VPWR _0267_ 0.47679f
C15602 _0380_ _0379_ 0.6803f
C15603 _0195_ _0852_/a_35_297# 0
C15604 hold18/a_49_47# net247 0.06774f
C15605 VPWR _0772_/a_79_21# 0.44522f
C15606 _0376_ _0606_/a_215_297# 0
C15607 _0234_ _0606_/a_465_297# 0
C15608 net45 _1017_/a_592_47# 0
C15609 _1020_/a_27_47# _0461_ 0.00121f
C15610 VPWR _1062_/a_1017_47# 0
C15611 _1018_/a_466_413# _0347_ 0
C15612 _1039_/a_592_47# _0172_ 0
C15613 _1021_/a_975_413# VPWR 0.00515f
C15614 hold58/a_49_47# _0557_/a_240_47# 0
C15615 net219 clknet_1_1__leaf__0461_ 0
C15616 _0762_/a_215_47# _0383_ 0.01004f
C15617 net180 _0953_/a_32_297# 0.00511f
C15618 _0179_ _0350_ 0.22943f
C15619 net149 _0526_/a_27_47# 0
C15620 _0424_ _0291_ 0.00448f
C15621 _1000_/a_193_47# _0773_/a_35_297# 0.00909f
C15622 net56 _0720_/a_68_297# 0
C15623 _0346_ _0811_/a_299_297# 0.00872f
C15624 _1009_/a_27_47# _1009_/a_193_47# 0.97445f
C15625 net207 _0181_ 0
C15626 clknet_1_1__leaf__0460_ _0694_/a_113_47# 0
C15627 _0421_ _0296_ 0.02019f
C15628 _0410_ clkbuf_1_1__f__0459_/a_110_47# 0
C15629 _0642_/a_215_297# VPWR 0.18337f
C15630 _1065_/a_891_413# _1065_/a_1017_47# 0.00617f
C15631 B[4] _0175_ 0.00354f
C15632 _0717_/a_80_21# _0707_/a_75_199# 0
C15633 _0508_/a_384_47# _0185_ 0
C15634 hold66/a_391_47# _1005_/a_466_413# 0
C15635 _1036_/a_27_47# net121 0.03908f
C15636 _0186_ _0522_/a_109_297# 0.0116f
C15637 net111 _1025_/a_27_47# 0.23013f
C15638 _1068_/a_891_413# _0487_ 0
C15639 net1 _0485_ 0.11536f
C15640 _0992_/a_1059_315# _0811_/a_81_21# 0
C15641 hold11/a_285_47# _0498_/a_51_297# 0
C15642 net31 net173 0.16743f
C15643 _0707_/a_75_199# _0339_ 0.10576f
C15644 _0707_/a_201_297# _0338_ 0.00327f
C15645 _0707_/a_544_297# _0335_ 0
C15646 comp0.B\[1\] _0565_/a_51_297# 0.01595f
C15647 _0172_ clknet_1_1__leaf__0458_ 0
C15648 _0453_ _0265_ 0.2231f
C15649 _1014_/a_634_159# _1014_/a_592_47# 0
C15650 _1071_/a_634_159# _1071_/a_466_413# 0.23992f
C15651 _1071_/a_193_47# _1071_/a_1059_315# 0.03405f
C15652 _1071_/a_27_47# _1071_/a_891_413# 0.03224f
C15653 _1015_/a_634_159# _0208_ 0.03569f
C15654 _1015_/a_891_413# _0173_ 0
C15655 net27 control0.sh 0.62738f
C15656 VPWR net51 2.03186f
C15657 _0573_/a_27_47# _1014_/a_27_47# 0
C15658 _0985_/a_381_47# _0458_ 0.00728f
C15659 net61 _0828_/a_113_297# 0.01729f
C15660 _0798_/a_199_47# net5 0
C15661 net36 B[1] 0
C15662 _0476_ _1034_/a_1059_315# 0.00234f
C15663 _0179_ _0149_ 0
C15664 _0320_ _0345_ 0.06834f
C15665 _0183_ _0244_ 0.10828f
C15666 _0217_ _0388_ 0
C15667 _0499_/a_145_75# _0175_ 0
C15668 hold54/a_285_47# clknet_0__0463_ 0
C15669 pp[29] _0335_ 0.00494f
C15670 _0362_ VPWR 0.42538f
C15671 _0836_/a_68_297# _0989_/a_193_47# 0
C15672 VPWR _0536_/a_240_47# 0.00139f
C15673 pp[28] acc0.A\[30\] 0
C15674 _0438_ net62 0
C15675 net120 net203 0.02778f
C15676 _0435_ pp[3] 0
C15677 _0437_ _0989_/a_27_47# 0.03866f
C15678 net212 _0989_/a_193_47# 0.00124f
C15679 _0347_ acc0.A\[13\] 0
C15680 hold25/a_49_47# hold25/a_391_47# 0.00188f
C15681 _0305_ _1059_/a_466_413# 0.01177f
C15682 VPWR _0638_/a_109_297# 0.00726f
C15683 _0551_/a_27_47# _0181_ 0
C15684 hold98/a_49_47# net41 0.00832f
C15685 _0098_ net219 0
C15686 net45 _0581_/a_373_47# 0.00156f
C15687 _0719_/a_27_47# _0462_ 0.00589f
C15688 _0285_ _0286_ 0.58309f
C15689 _0284_ _0283_ 0
C15690 _1015_/a_193_47# net17 0.00211f
C15691 net47 acc0.A\[6\] 0
C15692 net2 _0510_/a_373_47# 0
C15693 _1026_/a_561_413# acc0.A\[25\] 0
C15694 _0454_ _0852_/a_285_47# 0.00206f
C15695 net130 net148 0
C15696 _0081_ _0852_/a_35_297# 0
C15697 net36 _1039_/a_634_159# 0.01728f
C15698 _0462_ _0460_ 0.48141f
C15699 net88 _1067_/a_634_159# 0
C15700 _0195_ _1048_/a_193_47# 0
C15701 hold18/a_391_47# _0846_/a_149_47# 0
C15702 hold18/a_285_47# _0846_/a_240_47# 0
C15703 _0390_ _0772_/a_79_21# 0.00581f
C15704 _0770_/a_79_21# _0391_ 0
C15705 _1042_/a_193_47# _0542_/a_51_297# 0
C15706 _1012_/a_193_47# _0352_ 0.04426f
C15707 net54 hold9/a_49_47# 0.01104f
C15708 _0819_/a_81_21# _0427_ 0.00237f
C15709 _0470_ control0.sh 0
C15710 _0343_ _1016_/a_466_413# 0.00557f
C15711 _0172_ _1047_/a_27_47# 0
C15712 _1033_/a_27_47# _0175_ 0
C15713 net188 net3 0
C15714 clknet_1_0__leaf__0462_ _0575_/a_373_47# 0
C15715 _0582_/a_109_297# acc0.A\[18\] 0
C15716 _0831_/a_285_47# acc0.A\[6\] 0
C15717 acc0.A\[22\] _0590_/a_113_47# 0
C15718 clknet_1_0__leaf__0465_ hold83/a_285_47# 0.00199f
C15719 _0294_ clkbuf_0__0461_/a_110_47# 0.022f
C15720 comp0.B\[13\] _0537_/a_68_297# 0.16826f
C15721 net69 _0850_/a_68_297# 0
C15722 _0216_ _1010_/a_466_413# 0
C15723 _0981_/a_109_47# net167 0.00361f
C15724 _0981_/a_373_47# _0490_ 0.00165f
C15725 net48 net51 0.11283f
C15726 acc0.A\[12\] _0276_ 0.00629f
C15727 _1052_/a_466_413# _0180_ 0.00971f
C15728 _0318_ _0219_ 0.04796f
C15729 hold49/a_285_47# net196 0.00968f
C15730 _1016_/a_634_159# acc0.A\[17\] 0
C15731 _1033_/a_891_413# clknet_1_1__leaf_clk 0
C15732 _0963_/a_117_297# control0.count\[1\] 0.002f
C15733 net234 _0112_ 0
C15734 _1037_/a_891_413# _1036_/a_891_413# 0
C15735 _0702_/a_113_47# _0332_ 0
C15736 _0273_ _0435_ 0.14437f
C15737 _0553_/a_240_47# net29 0.06031f
C15738 _0533_/a_27_297# _0181_ 0.05211f
C15739 output37/a_27_47# _1057_/a_891_413# 0
C15740 _0223_ _0367_ 0.00123f
C15741 _0424_ _0290_ 0.03089f
C15742 net175 clkbuf_1_0__f__0464_/a_110_47# 0.00214f
C15743 hold24/a_285_47# hold25/a_49_47# 0
C15744 hold23/a_49_47# _0197_ 0.11837f
C15745 _0130_ net1 0
C15746 _0346_ _0091_ 0.00319f
C15747 net85 _0347_ 0.00398f
C15748 _0607_/a_27_297# _0309_ 0
C15749 _0498_/a_240_47# net7 0.06611f
C15750 net22 _0546_/a_240_47# 0
C15751 _0084_ _0986_/a_193_47# 0.17523f
C15752 _0445_ _0986_/a_466_413# 0
C15753 _0713_/a_27_47# _0782_/a_27_47# 0.00103f
C15754 net214 _0428_ 0.13467f
C15755 net10 net20 0.02681f
C15756 _0357_ acc0.A\[29\] 0.0211f
C15757 _0399_ _0988_/a_634_159# 0.00482f
C15758 net56 net116 0
C15759 comp0.B\[2\] _1033_/a_975_413# 0
C15760 _0464_ clknet_0__0464_ 0.03181f
C15761 _0305_ _0392_ 0
C15762 net150 _1005_/a_561_413# 0
C15763 _0183_ _1005_/a_1059_315# 0
C15764 _0971_/a_81_21# _0950_/a_75_212# 0
C15765 net168 input14/a_75_212# 0
C15766 net190 _1028_/a_975_413# 0
C15767 _0126_ _1028_/a_891_413# 0
C15768 clknet_1_1__leaf__0459_ _0798_/a_113_297# 0.0091f
C15769 _0387_ _0307_ 0
C15770 _0180_ _0194_ 0.22117f
C15771 _1032_/a_634_159# _0565_/a_51_297# 0
C15772 pp[9] _1057_/a_466_413# 0
C15773 _0573_/a_27_47# _0195_ 0
C15774 VPWR _1046_/a_27_47# 0.43681f
C15775 _1022_/a_193_47# _1022_/a_634_159# 0.12729f
C15776 _1022_/a_27_47# _1022_/a_466_413# 0.27314f
C15777 acc0.A\[31\] _1013_/a_466_413# 0
C15778 net162 _1013_/a_193_47# 0
C15779 _0576_/a_373_47# acc0.A\[23\] 0.00226f
C15780 _0178_ _0584_/a_109_297# 0
C15781 _1003_/a_561_413# clknet_1_0__leaf__0460_ 0
C15782 _1021_/a_466_413# _0462_ 0
C15783 _1059_/a_561_413# acc0.A\[15\] 0
C15784 net106 _0181_ 0.12069f
C15785 _0717_/a_303_47# pp[27] 0
C15786 VPWR _0775_/a_510_47# 0.00113f
C15787 clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ 1.66563f
C15788 _0730_/a_79_21# _0331_ 0
C15789 _0811_/a_81_21# _0421_ 0.00378f
C15790 net61 _0433_ 0.26546f
C15791 _0259_ _0399_ 0.0292f
C15792 clknet_1_1__leaf__0461_ _0352_ 0.02876f
C15793 hold20/a_391_47# VPWR 0.19465f
C15794 _0957_/a_32_297# comp0.B\[6\] 0.02513f
C15795 _1018_/a_381_47# _0116_ 0.1266f
C15796 _1018_/a_592_47# net206 0
C15797 _0356_ _0333_ 0.1972f
C15798 _1008_/a_193_47# net94 0.00455f
C15799 _1008_/a_1059_315# _1008_/a_1017_47# 0
C15800 _1055_/a_193_47# _1055_/a_381_47# 0.09799f
C15801 _1055_/a_634_159# _1055_/a_891_413# 0.03684f
C15802 _1055_/a_27_47# _1055_/a_561_413# 0.0027f
C15803 _0774_/a_68_297# _0242_ 0
C15804 B[13] net19 0
C15805 _0337_ _1011_/a_891_413# 0
C15806 pp[16] _0995_/a_891_413# 0
C15807 net53 _1025_/a_975_413# 0.00101f
C15808 _0559_/a_51_297# _0208_ 0.19682f
C15809 _0559_/a_149_47# _0173_ 0.02033f
C15810 net121 comp0.B\[3\] 0
C15811 _0771_/a_27_413# _0771_/a_215_297# 0.14121f
C15812 _1003_/a_27_47# _1003_/a_891_413# 0.03224f
C15813 _1003_/a_193_47# _1003_/a_1059_315# 0.03405f
C15814 _1003_/a_634_159# _1003_/a_466_413# 0.23992f
C15815 hold97/a_49_47# _0321_ 0.00796f
C15816 _1055_/a_1059_315# net181 0
C15817 net23 comp0.B\[6\] 0
C15818 _0855_/a_81_21# _1019_/a_1059_315# 0
C15819 _0679_/a_68_297# _0310_ 0.11485f
C15820 clknet_0__0458_ _0986_/a_1017_47# 0
C15821 hold69/a_49_47# _0294_ 0.0023f
C15822 _0466_ _0974_/a_79_199# 0.07833f
C15823 VPWR _0970_/a_27_297# 0.45948f
C15824 hold58/a_285_47# hold58/a_391_47# 0.41909f
C15825 hold81/a_49_47# net228 0
C15826 _0176_ _0542_/a_240_47# 0.00384f
C15827 _0343_ clkbuf_1_1__f__0458_/a_110_47# 0
C15828 _0155_ net3 0
C15829 _1054_/a_27_47# net15 0.02478f
C15830 _0525_/a_299_297# net148 0
C15831 net46 _0099_ 0.00245f
C15832 _0997_/a_1059_315# _0219_ 0
C15833 _0453_ _0267_ 0
C15834 _0833_/a_510_47# _0439_ 0.00181f
C15835 _1004_/a_891_413# _0758_/a_215_47# 0
C15836 _1004_/a_193_47# _0347_ 0
C15837 _0182_ clknet_1_1__leaf__0457_ 0.29708f
C15838 VPWR _0833_/a_510_47# 0
C15839 net62 clknet_1_1__leaf__0465_ 0
C15840 _0126_ _0739_/a_79_21# 0
C15841 hold87/a_285_47# _0181_ 0.08314f
C15842 _0847_/a_109_297# acc0.A\[15\] 0
C15843 _1054_/a_27_47# _1053_/a_1059_315# 0
C15844 _0799_/a_80_21# _0799_/a_209_297# 0.06257f
C15845 _0465_ _0219_ 0.01366f
C15846 _0559_/a_240_47# _0212_ 0
C15847 _0982_/a_891_413# _0456_ 0.01534f
C15848 _0982_/a_975_413# net234 0
C15849 _0144_ _0147_ 0.00104f
C15850 _0222_ _0756_/a_285_47# 0
C15851 _0598_/a_79_21# VPWR 0.23604f
C15852 _1058_/a_193_47# net189 0.02663f
C15853 _1056_/a_975_413# net182 0
C15854 _0811_/a_81_21# _0809_/a_81_21# 0.00351f
C15855 _0222_ _0749_/a_299_297# 0
C15856 _0557_/a_149_47# _0554_/a_68_297# 0
C15857 acc0.A\[2\] _0219_ 0.00218f
C15858 _0718_/a_47_47# _0707_/a_75_199# 0.00775f
C15859 net43 clknet_0__0461_ 0.22585f
C15860 _0409_ hold91/a_391_47# 0
C15861 VPWR _0178_ 0.73115f
C15862 _0343_ pp[14] 0.04983f
C15863 net236 _0974_/a_79_199# 0
C15864 _0985_/a_891_413# _0268_ 0
C15865 _0985_/a_27_47# hold71/a_49_47# 0
C15866 net45 _0347_ 0.62076f
C15867 hold100/a_49_47# _0452_ 0
C15868 _0098_ _0352_ 0.27059f
C15869 _0399_ net221 0
C15870 _1059_/a_466_413# _0181_ 0
C15871 pp[30] _0338_ 0.00557f
C15872 _1000_/a_1059_315# _0769_/a_81_21# 0
C15873 _0387_ _0780_/a_285_297# 0.00769f
C15874 _0366_ _0360_ 0
C15875 net208 _0336_ 0.04763f
C15876 _0982_/a_193_47# _0452_ 0
C15877 _0982_/a_27_47# _0266_ 0
C15878 _1016_/a_975_413# clknet_1_1__leaf__0461_ 0
C15879 _1048_/a_27_47# _1048_/a_634_159# 0.14145f
C15880 clknet_1_0__leaf_clk _1064_/a_466_413# 0
C15881 _0225_ _0373_ 0
C15882 _1015_/a_466_413# _0178_ 0
C15883 _0717_/a_209_47# pp[28] 0
C15884 _0106_ hold50/a_285_47# 0.00234f
C15885 _0223_ _0742_/a_299_297# 0
C15886 _0179_ clkload2/a_268_47# 0.00113f
C15887 net116 _0345_ 0.00811f
C15888 _0548_/a_51_297# _0138_ 0.10689f
C15889 _0548_/a_240_47# net173 0.04504f
C15890 _0555_/a_51_297# VPWR 0.49304f
C15891 _0556_/a_68_297# _0556_/a_150_297# 0.00477f
C15892 _0506_/a_81_21# net229 0.06169f
C15893 _0251_ _0826_/a_27_53# 0
C15894 _0415_ VPWR 0.38752f
C15895 VPWR _1033_/a_381_47# 0.07064f
C15896 init input23/a_75_212# 0
C15897 _1044_/a_1059_315# _0141_ 0.02588f
C15898 clknet_1_0__leaf__0465_ _1049_/a_381_47# 0
C15899 net1 _0761_/a_113_47# 0
C15900 _0501_/a_27_47# clkbuf_1_1__f__0457_/a_110_47# 0
C15901 net190 net191 0
C15902 VPWR _1050_/a_1017_47# 0
C15903 _0598_/a_79_21# net48 0
C15904 net36 _1041_/a_891_413# 0
C15905 _0286_ _0218_ 0
C15906 _0179_ _0519_/a_384_47# 0
C15907 _0151_ _1054_/a_193_47# 0
C15908 net61 _0636_/a_145_75# 0.00225f
C15909 net45 _0792_/a_209_297# 0
C15910 hold57/a_49_47# hold57/a_285_47# 0.22264f
C15911 input19/a_75_212# _1042_/a_27_47# 0
C15912 _1010_/a_466_413# _1010_/a_561_413# 0.00772f
C15913 _1010_/a_634_159# _1010_/a_975_413# 0
C15914 clknet_1_0__leaf__0462_ _1004_/a_561_413# 0
C15915 _0276_ net42 0.01256f
C15916 _1056_/a_193_47# _0514_/a_109_297# 0
C15917 _0924_/a_27_47# _0174_ 0
C15918 hold55/a_285_47# _1015_/a_193_47# 0.0148f
C15919 hold55/a_391_47# _1015_/a_27_47# 0.0042f
C15920 hold92/a_285_47# _0345_ 0.00219f
C15921 _0465_ _0826_/a_301_297# 0
C15922 _0991_/a_561_413# _0181_ 0
C15923 hold6/a_49_47# _0546_/a_51_297# 0.00372f
C15924 _0978_/a_27_297# _0978_/a_109_297# 0.17136f
C15925 _1040_/a_27_47# _1040_/a_561_413# 0.00163f
C15926 _1040_/a_634_159# _1040_/a_891_413# 0.03684f
C15927 _1040_/a_193_47# _1040_/a_381_47# 0.09503f
C15928 hold36/a_285_47# net194 0
C15929 _0795_/a_81_21# _0795_/a_299_297# 0.08213f
C15930 _0266_ _0446_ 0.01376f
C15931 hold79/a_391_47# _0976_/a_76_199# 0
C15932 _0979_/a_27_297# _0979_/a_109_47# 0.00393f
C15933 _0399_ _0782_/a_27_47# 0.32981f
C15934 _0181_ _0392_ 0
C15935 _0326_ clknet_0__0460_ 0.03931f
C15936 _0697_/a_300_47# _0328_ 0.00119f
C15937 _0519_/a_299_297# net75 0
C15938 _0527_/a_27_297# _0527_/a_109_47# 0.00393f
C15939 _0216_ _1027_/a_193_47# 0.24998f
C15940 VPWR _1019_/a_27_47# 0.42703f
C15941 _0532_/a_81_21# clkbuf_1_1__f__0457_/a_110_47# 0
C15942 _0743_/a_51_297# hold90/a_285_47# 0.00175f
C15943 clknet_0__0463_ _0562_/a_68_297# 0.016f
C15944 net63 VPWR 1.62837f
C15945 acc0.A\[14\] _0996_/a_634_159# 0.00708f
C15946 net45 _1016_/a_891_413# 0.002f
C15947 net101 clknet_1_0__leaf__0457_ 0
C15948 _1067_/a_193_47# _1067_/a_381_47# 0.09503f
C15949 _1067_/a_634_159# _1067_/a_891_413# 0.03684f
C15950 _1067_/a_27_47# _1067_/a_561_413# 0.0027f
C15951 control0.add _0616_/a_78_199# 0.00922f
C15952 _0174_ net180 0.52055f
C15953 _0800_/a_51_297# _0410_ 0
C15954 clknet_1_0__leaf__0459_ _0775_/a_510_47# 0
C15955 _1001_/a_27_47# _0345_ 0.03354f
C15956 _0805_/a_27_47# _0805_/a_181_47# 0.00401f
C15957 _0314_ _0682_/a_150_297# 0
C15958 _0172_ comp0.B\[10\] 0.02571f
C15959 hold35/a_49_47# input2/a_75_212# 0
C15960 _0462_ _0614_/a_29_53# 0.00244f
C15961 _0985_/a_193_47# _0529_/a_27_297# 0
C15962 _0985_/a_27_47# _0529_/a_109_297# 0
C15963 _1000_/a_466_413# _0392_ 0
C15964 _1072_/a_634_159# _1071_/a_891_413# 0
C15965 _1072_/a_466_413# _1071_/a_1059_315# 0
C15966 net199 _0347_ 0.00777f
C15967 VPWR _0324_ 1.86709f
C15968 clknet_1_1__leaf__0460_ _0350_ 0.37178f
C15969 _1004_/a_27_47# _0757_/a_68_297# 0
C15970 VPWR _0581_/a_373_47# 0
C15971 _0620_/a_113_47# _0252_ 0.01006f
C15972 _0183_ _0592_/a_68_297# 0
C15973 net97 _0332_ 0.00847f
C15974 _1009_/a_466_413# _1009_/a_592_47# 0.00553f
C15975 _1009_/a_634_159# _1009_/a_1017_47# 0
C15976 net65 _0989_/a_466_413# 0.01453f
C15977 acc0.A\[7\] _0989_/a_634_159# 0.00324f
C15978 _0252_ _0989_/a_27_47# 0.10333f
C15979 _0252_ hold1/a_49_47# 0
C15980 net36 net147 0
C15981 _0989_/a_634_159# _0989_/a_1059_315# 0
C15982 _0989_/a_27_47# _0989_/a_381_47# 0.06222f
C15983 _0989_/a_193_47# _0989_/a_891_413# 0.1932f
C15984 comp0.B\[13\] hold36/a_391_47# 0
C15985 _0956_/a_304_297# net201 0
C15986 hold16/a_285_47# hold92/a_49_47# 0
C15987 _0348_ _0707_/a_201_297# 0.01548f
C15988 _0717_/a_80_21# _0338_ 0.02615f
C15989 _0717_/a_209_297# _0335_ 0.01182f
C15990 _0982_/a_592_47# VPWR 0
C15991 clknet_0_clk _0160_ 0
C15992 _0476_ _1066_/a_975_413# 0
C15993 _0399_ _0253_ 0.10898f
C15994 _1013_/a_466_413# net43 0
C15995 hold66/a_391_47# _0103_ 0
C15996 _0992_/a_634_159# _0992_/a_1059_315# 0
C15997 _0992_/a_27_47# _0992_/a_381_47# 0.06222f
C15998 _0992_/a_193_47# _0992_/a_891_413# 0.19549f
C15999 _0629_/a_59_75# _0346_ 0
C16000 net24 _0563_/a_512_297# 0
C16001 _0695_/a_217_297# clkbuf_1_0__f__0462_/a_110_47# 0
C16002 net7 net173 0.03208f
C16003 net161 net23 0
C16004 _0606_/a_297_297# VPWR 0
C16005 _1002_/a_27_47# _0603_/a_68_297# 0
C16006 _0166_ _0162_ 0
C16007 VPWR _1053_/a_891_413# 0.18826f
C16008 acc0.A\[16\] _0674_/a_113_47# 0
C16009 _0607_/a_373_47# net43 0.00131f
C16010 _0718_/a_285_47# pp[27] 0.00285f
C16011 _0125_ _1027_/a_1059_315# 0.01636f
C16012 acc0.A\[27\] _1027_/a_561_413# 0
C16013 net54 _0739_/a_79_21# 0.01176f
C16014 _0338_ _0339_ 0
C16015 _0280_ _0655_/a_369_297# 0.00292f
C16016 hold10/a_49_47# control0.reset 0
C16017 _0355_ _1029_/a_193_47# 0
C16018 _0274_ clkbuf_0__0458_/a_110_47# 0.00151f
C16019 _0470_ _0955_/a_32_297# 0.0088f
C16020 _0959_/a_80_21# comp0.B\[5\] 0
C16021 _1014_/a_891_413# acc0.A\[0\] 0.02742f
C16022 _0996_/a_561_413# _0410_ 0
C16023 _0996_/a_975_413# net238 0
C16024 _1045_/a_1059_315# _1043_/a_193_47# 0
C16025 _1045_/a_891_413# _1043_/a_27_47# 0
C16026 _0835_/a_215_47# _0218_ 0.00262f
C16027 hold75/a_285_47# _0267_ 0.0351f
C16028 clknet_0__0458_ _0846_/a_51_297# 0.01368f
C16029 _0957_/a_32_297# net26 0.00444f
C16030 _0481_ _0976_/a_76_199# 0
C16031 _0935_/a_27_47# _1061_/a_193_47# 0.00716f
C16032 hold76/a_49_47# _0461_ 0.0081f
C16033 hold10/a_285_47# _1061_/a_1059_315# 0
C16034 _0983_/a_193_47# net206 0
C16035 _1061_/a_27_47# _1061_/a_634_159# 0.14145f
C16036 net187 hold40/a_391_47# 0.13331f
C16037 _0429_ _0437_ 0.09919f
C16038 _0251_ _0087_ 0.01194f
C16039 _0458_ _0147_ 0
C16040 _0343_ _0408_ 0.02426f
C16041 _0659_/a_68_297# _0990_/a_634_159# 0
C16042 _0626_/a_68_297# _0257_ 0.10424f
C16043 _0124_ _1026_/a_634_159# 0.00122f
C16044 _0572_/a_27_297# net112 0
C16045 net155 _1026_/a_891_413# 0.00143f
C16046 _0216_ _1026_/a_1059_315# 0.0866f
C16047 net23 net26 0.0288f
C16048 _1007_/a_1059_315# _0345_ 0
C16049 _1007_/a_27_47# _0219_ 0.0012f
C16050 A[10] input16/a_75_212# 0.00355f
C16051 _0553_/a_240_47# comp0.B\[6\] 0.00126f
C16052 clknet_1_1__leaf__0459_ net41 0.02016f
C16053 _0689_/a_68_297# _0360_ 0
C16054 _0319_ _0737_/a_35_297# 0.00297f
C16055 clkbuf_0__0459_/a_110_47# _0507_/a_27_297# 0.00339f
C16056 _0795_/a_81_21# net6 0
C16057 _0313_ _0570_/a_27_297# 0
C16058 _0176_ B[11] 0.00541f
C16059 _0817_/a_266_47# acc0.A\[9\] 0.00757f
C16060 _0817_/a_266_297# _0288_ 0
C16061 _0549_/a_150_297# _0207_ 0
C16062 _0420_ _0345_ 0.01897f
C16063 A[14] pp[14] 0.17233f
C16064 _0305_ _0157_ 0
C16065 _0190_ _0988_/a_634_159# 0
C16066 net16 _0988_/a_1059_315# 0
C16067 _0343_ _0291_ 0.02123f
C16068 _0186_ _0150_ 0.05277f
C16069 _0804_/a_79_21# _0414_ 0.0021f
C16070 clkbuf_1_0__f__0459_/a_110_47# _1016_/a_466_413# 0
C16071 hold2/a_285_47# _1047_/a_27_47# 0
C16072 hold2/a_49_47# _1047_/a_193_47# 0
C16073 _0243_ _1019_/a_193_47# 0
C16074 _1020_/a_381_47# acc0.A\[20\] 0
C16075 net36 net125 0.21395f
C16076 _0183_ _1014_/a_27_47# 0
C16077 _0217_ _1014_/a_634_159# 0.04126f
C16078 _1042_/a_891_413# _0203_ 0
C16079 _0977_/a_75_212# _1069_/a_27_47# 0.01019f
C16080 _1065_/a_27_47# clknet_1_0__leaf__0457_ 0
C16081 _0464_ _0536_/a_51_297# 0
C16082 acc0.A\[1\] _0530_/a_81_21# 0
C16083 _0459_ _0345_ 0.00558f
C16084 clknet_1_1__leaf__0463_ _0163_ 0
C16085 _0805_/a_27_47# _0993_/a_27_47# 0
C16086 _0343_ net166 0.02168f
C16087 _0984_/a_381_47# acc0.A\[15\] 0.00169f
C16088 clknet_1_1__leaf__0459_ net217 0.09033f
C16089 _0569_/a_109_297# _1029_/a_27_47# 0
C16090 _0569_/a_27_297# _1029_/a_193_47# 0
C16091 net67 acc0.A\[10\] 0.3848f
C16092 VPWR _1028_/a_1059_315# 0.39842f
C16093 _1069_/a_634_159# _1069_/a_381_47# 0
C16094 hold4/a_285_47# net177 0
C16095 hold4/a_391_47# net109 0.01926f
C16096 _0996_/a_27_47# net228 0
C16097 VPWR _0812_/a_79_21# 0.46673f
C16098 _1059_/a_27_47# acc0.A\[13\] 0.00299f
C16099 _0673_/a_103_199# _0218_ 0
C16100 net56 _0220_ 0.00147f
C16101 _0954_/a_32_297# comp0.B\[11\] 0.11555f
C16102 _0433_ _0431_ 0.00198f
C16103 _1037_/a_1059_315# comp0.B\[4\] 0
C16104 _1041_/a_634_159# _1040_/a_27_47# 0
C16105 _1041_/a_193_47# _1040_/a_193_47# 0
C16106 _1041_/a_27_47# _1040_/a_634_159# 0
C16107 _1031_/a_634_159# _0220_ 0.02213f
C16108 _1031_/a_193_47# _0336_ 0
C16109 _0536_/a_149_47# _0172_ 0.00356f
C16110 input31/a_75_212# net22 0.00523f
C16111 hold66/a_49_47# _0369_ 0.04352f
C16112 _0399_ _1017_/a_27_47# 0
C16113 _0571_/a_109_297# acc0.A\[26\] 0
C16114 pp[15] output43/a_27_47# 0.01068f
C16115 _0199_ _0181_ 0.02087f
C16116 pp[20] output49/a_27_47# 0.00337f
C16117 hold85/a_49_47# _0466_ 0
C16118 _0495_/a_68_297# clknet_1_1__leaf__0457_ 0
C16119 comp0.B\[2\] _0956_/a_304_297# 0.00106f
C16120 _1059_/a_891_413# hold82/a_49_47# 0.00267f
C16121 _1059_/a_466_413# hold82/a_391_47# 0
C16122 input20/a_75_212# hold51/a_49_47# 0
C16123 _1030_/a_634_159# net209 0
C16124 input24/a_75_212# net24 0.10858f
C16125 _0596_/a_59_75# _0217_ 0
C16126 _1051_/a_193_47# net9 0
C16127 _1018_/a_193_47# clknet_0__0461_ 0.00109f
C16128 net99 _0339_ 0
C16129 _0337_ output56/a_27_47# 0
C16130 clknet_1_1__leaf__0459_ _0744_/a_27_47# 0.0024f
C16131 _1002_/a_634_159# _0181_ 0
C16132 _0480_ _0978_/a_27_297# 0
C16133 _0592_/a_150_297# _0379_ 0
C16134 net172 _0136_ 0
C16135 _0743_/a_149_47# clkbuf_1_0__f__0462_/a_110_47# 0
C16136 _0258_ _0434_ 0
C16137 _1034_/a_466_413# _0176_ 0
C16138 _0172_ _0218_ 0.01367f
C16139 _0312_ _0460_ 0.01638f
C16140 _0233_ _0350_ 0.0303f
C16141 clknet_1_1__leaf__0462_ _1008_/a_1017_47# 0
C16142 comp0.B\[5\] _0173_ 0.10584f
C16143 _1032_/a_1059_315# net201 0
C16144 comp0.B\[6\] _0213_ 0.17624f
C16145 _0216_ _0367_ 0
C16146 hold43/a_391_47# clknet_1_1__leaf__0462_ 0.00256f
C16147 pp[9] net189 0
C16148 clknet_1_0__leaf__0463_ input31/a_75_212# 0.00898f
C16149 _0183_ hold18/a_391_47# 0.00155f
C16150 _1014_/a_27_47# acc0.A\[15\] 0
C16151 _1022_/a_1059_315# _1022_/a_1017_47# 0
C16152 _1022_/a_27_47# net151 0.10918f
C16153 hold75/a_391_47# _0218_ 0.02284f
C16154 comp0.B\[7\] _0159_ 0.00286f
C16155 clknet_1_1__leaf__0461_ hold72/a_285_47# 0
C16156 _0645_/a_377_297# _0276_ 0
C16157 _1065_/a_27_47# _1062_/a_466_413# 0
C16158 clknet_1_0__leaf__0459_ _1019_/a_27_47# 0.01817f
C16159 _0119_ _0462_ 0.00165f
C16160 hold2/a_285_47# clknet_1_0__leaf__0461_ 0
C16161 _0174_ _0545_/a_150_297# 0
C16162 clkbuf_1_0__f__0462_/a_110_47# _0345_ 0.11846f
C16163 _0316_ VPWR 1.63391f
C16164 _0265_ _0345_ 0.27843f
C16165 _0456_ clkbuf_0__0457_/a_110_47# 0
C16166 net199 _1025_/a_27_47# 0.00163f
C16167 acc0.A\[16\] _0307_ 0.06258f
C16168 _0994_/a_193_47# _0994_/a_381_47# 0.09972f
C16169 _0994_/a_634_159# _0994_/a_891_413# 0.03684f
C16170 _0994_/a_27_47# _0994_/a_561_413# 0.0027f
C16171 _1020_/a_466_413# clknet_1_0__leaf__0457_ 0.00939f
C16172 _0285_ net79 0.00411f
C16173 _0284_ _0808_/a_266_47# 0
C16174 _0475_ _0474_ 0.17661f
C16175 VPWR hold5/a_49_47# 0.33635f
C16176 _0292_ net217 0.00451f
C16177 B[9] net32 0.00949f
C16178 _1055_/a_1059_315# net179 0.00105f
C16179 _1055_/a_891_413# net141 0
C16180 net247 _0448_ 0
C16181 acc0.A\[24\] _0360_ 0
C16182 VPWR hold3/a_391_47# 0.2183f
C16183 _1023_/a_27_47# net51 0.045f
C16184 _1023_/a_466_413# output51/a_27_47# 0.00198f
C16185 hold5/a_391_47# _1043_/a_891_413# 0
C16186 _0422_ hold81/a_391_47# 0
C16187 hold22/a_49_47# _1053_/a_193_47# 0
C16188 hold22/a_285_47# _1053_/a_27_47# 0
C16189 _0305_ acc0.A\[9\] 0
C16190 _0984_/a_381_47# _0179_ 0
C16191 VPWR _0347_ 6.55966f
C16192 net23 hold84/a_285_47# 0
C16193 _0608_/a_27_47# _0239_ 0.00471f
C16194 _0343_ _0621_/a_285_297# 0.0381f
C16195 _1003_/a_466_413# net89 0
C16196 _1003_/a_634_159# _0101_ 0.04443f
C16197 net36 _1047_/a_1059_315# 0.06673f
C16198 net36 _0473_ 0.02006f
C16199 _0954_/a_32_297# _0202_ 0.01558f
C16200 _0648_/a_27_297# _0404_ 0.01532f
C16201 hold26/a_285_47# _0174_ 0.04955f
C16202 _0217_ _0216_ 0.43105f
C16203 _0183_ _0195_ 0.1893f
C16204 comp0.B\[1\] _0584_/a_109_297# 0
C16205 _1039_/a_27_47# _1039_/a_634_159# 0.13601f
C16206 _0967_/a_487_297# VPWR 0.00443f
C16207 comp0.B\[11\] net173 0
C16208 _0836_/a_150_297# clknet_1_1__leaf__0458_ 0
C16209 hold56/a_285_47# clknet_1_1__leaf_clk 0
C16210 _1020_/a_193_47# _0457_ 0.00991f
C16211 _0197_ _0529_/a_109_297# 0.00353f
C16212 _0343_ _0290_ 0
C16213 _0212_ comp0.B\[6\] 0
C16214 _1015_/a_27_47# _0352_ 0
C16215 comp0.B\[13\] net180 0.00226f
C16216 VPWR _0104_ 0.43349f
C16217 _0985_/a_27_47# net170 0
C16218 _0437_ clknet_1_1__leaf__0458_ 0.00202f
C16219 _0257_ _0252_ 0
C16220 _1010_/a_27_47# _0332_ 0
C16221 _1004_/a_975_413# _0102_ 0
C16222 _0729_/a_68_297# clknet_1_1__leaf__0462_ 0.00995f
C16223 _0518_/a_109_297# _0399_ 0
C16224 net33 _1062_/a_634_159# 0
C16225 _1026_/a_27_47# _1026_/a_193_47# 0.97453f
C16226 _0733_/a_448_47# _0737_/a_35_297# 0
C16227 hold41/a_391_47# net37 0
C16228 _0534_/a_384_47# net175 0
C16229 clknet_0__0458_ hold31/a_285_47# 0
C16230 _0983_/a_381_47# _0347_ 0.00583f
C16231 _0752_/a_27_413# _1005_/a_1059_315# 0.00174f
C16232 _1055_/a_193_47# clknet_1_1__leaf__0458_ 0
C16233 hold18/a_391_47# acc0.A\[15\] 0.0036f
C16234 net229 _0184_ 0.08935f
C16235 net140 _1053_/a_634_159# 0.02239f
C16236 net169 _1053_/a_193_47# 0
C16237 _0982_/a_27_47# _0399_ 0
C16238 _0222_ _0618_/a_297_297# 0.00379f
C16239 _0793_/a_512_297# net41 0
C16240 _0284_ _0345_ 0.01556f
C16241 _0500_/a_27_47# _0146_ 0
C16242 VPWR _0792_/a_209_297# 0.19447f
C16243 VPWR _0987_/a_1017_47# 0
C16244 _1024_/a_1059_315# _1024_/a_891_413# 0.31086f
C16245 _1024_/a_193_47# _1024_/a_975_413# 0
C16246 _1024_/a_466_413# _1024_/a_381_47# 0.03733f
C16247 hold23/a_285_47# net9 0
C16248 _0217_ _1067_/a_27_47# 0
C16249 net86 hold72/a_391_47# 0
C16250 _0502_/a_27_47# _0499_/a_59_75# 0
C16251 net150 _0383_ 0.01911f
C16252 _0348_ pp[30] 0.00214f
C16253 net48 hold3/a_391_47# 0
C16254 VPWR _0745_/a_109_47# 0
C16255 _0718_/a_47_47# _0338_ 0.00624f
C16256 _1021_/a_1059_315# _1020_/a_27_47# 0
C16257 hold56/a_391_47# clkbuf_1_1__f_clk/a_110_47# 0
C16258 clknet_1_1__leaf__0464_ _0542_/a_51_297# 0
C16259 _1011_/a_891_413# _0333_ 0
C16260 _0234_ _0600_/a_103_199# 0.00152f
C16261 _1036_/a_193_47# input25/a_75_212# 0
C16262 net61 _0835_/a_78_199# 0
C16263 _0220_ _0345_ 0.00266f
C16264 hold36/a_285_47# _1045_/a_27_47# 0.01222f
C16265 _0157_ _0181_ 0
C16266 _1000_/a_1017_47# _0244_ 0
C16267 VPWR _1029_/a_1017_47# 0
C16268 net46 _0238_ 0.08003f
C16269 _0514_/a_109_297# clknet_1_1__leaf__0465_ 0.00198f
C16270 _0644_/a_377_297# acc0.A\[13\] 0.00124f
C16271 _0180_ _1049_/a_193_47# 0
C16272 comp0.B\[2\] _1032_/a_1059_315# 0.01785f
C16273 _0982_/a_592_47# _0453_ 0
C16274 clk _1064_/a_1059_315# 0.00296f
C16275 hold96/a_391_47# _0217_ 0.05593f
C16276 _1048_/a_891_413# _1048_/a_975_413# 0.00851f
C16277 _1048_/a_27_47# net134 0.23149f
C16278 _1048_/a_381_47# _1048_/a_561_413# 0.00123f
C16279 hold42/a_285_47# A[10] 0
C16280 net47 _0611_/a_68_297# 0
C16281 clkbuf_1_1__f__0460_/a_110_47# _1010_/a_381_47# 0
C16282 _0712_/a_381_47# _0220_ 0
C16283 _1034_/a_561_413# clknet_1_1__leaf__0463_ 0
C16284 _0195_ acc0.A\[15\] 0.08939f
C16285 hold34/a_391_47# acc0.A\[9\] 0.00137f
C16286 _0831_/a_285_297# _0826_/a_27_53# 0
C16287 _0113_ _0178_ 0.00678f
C16288 clknet_1_1__leaf__0464_ _0142_ 0.0563f
C16289 net173 _0202_ 0
C16290 _0399_ net238 0.34815f
C16291 VPWR _0956_/a_114_297# 0.00671f
C16292 B[9] net10 0.03424f
C16293 VPWR _1016_/a_891_413# 0.17551f
C16294 _0339_ _0396_ 0
C16295 _0981_/a_27_297# clkbuf_0_clk/a_110_47# 0
C16296 _0600_/a_253_47# clkbuf_1_0__f__0460_/a_110_47# 0
C16297 _0490_ clknet_1_0__leaf_clk 0.00672f
C16298 _0734_/a_47_47# _0322_ 0
C16299 _0399_ _0446_ 0
C16300 VPWR comp0.B\[1\] 0.54901f
C16301 _0311_ clkbuf_0__0460_/a_110_47# 0
C16302 _1016_/a_466_413# clkbuf_0__0461_/a_110_47# 0
C16303 _1060_/a_634_159# _0219_ 0
C16304 net76 _0832_/a_113_47# 0
C16305 _0804_/a_79_21# _0404_ 0.0135f
C16306 _0232_ _0618_/a_510_47# 0.00331f
C16307 hold23/a_391_47# acc0.A\[3\] 0.00707f
C16308 _0172_ _0177_ 0.05711f
C16309 _0183_ _0081_ 0
C16310 _0569_/a_109_297# _1028_/a_891_413# 0
C16311 net152 _0204_ 0.14814f
C16312 hold27/a_391_47# VPWR 0.1661f
C16313 _0139_ _0544_/a_149_47# 0
C16314 _0349_ _0110_ 0
C16315 _0729_/a_68_297# net242 0.10246f
C16316 _0310_ _0678_/a_68_297# 0.10708f
C16317 clknet_1_1__leaf__0460_ _0731_/a_299_297# 0
C16318 pp[30] acc0.A\[31\] 0.00737f
C16319 net59 net162 0
C16320 _0217_ net247 0
C16321 _1051_/a_27_47# _0522_/a_27_297# 0
C16322 hold16/a_49_47# _0220_ 0.01364f
C16323 _0766_/a_109_297# _0310_ 0
C16324 _0179_ hold18/a_391_47# 0
C16325 clkbuf_1_0__f__0460_/a_110_47# _1006_/a_27_47# 0
C16326 VPWR clkbuf_0__0465_/a_110_47# 1.46352f
C16327 hold69/a_285_47# net216 0.01036f
C16328 _1056_/a_1059_315# net2 0
C16329 _1056_/a_634_159# _0189_ 0.00182f
C16330 _0130_ _1015_/a_975_413# 0
C16331 hold69/a_49_47# _0371_ 0.12103f
C16332 hold6/a_285_47# net32 0.02832f
C16333 hold6/a_391_47# net152 0
C16334 _1040_/a_1059_315# net174 0.05327f
C16335 _1053_/a_466_413# acc0.A\[6\] 0.00163f
C16336 _1053_/a_27_47# net13 0.00239f
C16337 clknet_1_0__leaf__0465_ _1054_/a_1059_315# 0
C16338 _0410_ _0277_ 0
C16339 _0433_ _0269_ 0
C16340 hold79/a_391_47# _0488_ 0.00337f
C16341 hold79/a_285_47# _0466_ 0.0045f
C16342 _1017_/a_381_47# acc0.A\[18\] 0
C16343 _0292_ net66 0
C16344 net63 _0523_/a_81_21# 0
C16345 _0250_ _1006_/a_27_47# 0
C16346 _0249_ _1006_/a_193_47# 0
C16347 _0256_ _0840_/a_68_297# 0
C16348 hold33/a_285_47# comp0.B\[7\] 0.01281f
C16349 _0111_ clknet_1_1__leaf__0459_ 0
C16350 _1072_/a_1059_315# _1072_/a_891_413# 0.31086f
C16351 _1072_/a_193_47# _1072_/a_975_413# 0
C16352 _1072_/a_466_413# _1072_/a_381_47# 0.03733f
C16353 _0195_ net156 0.04723f
C16354 _0841_/a_79_21# _0444_ 0.13864f
C16355 _0183_ _0505_/a_373_47# 0
C16356 net180 comp0.B\[9\] 0.0251f
C16357 _0216_ _0248_ 0.00116f
C16358 _0640_/a_215_297# _0640_/a_109_53# 0.08065f
C16359 _0852_/a_35_297# acc0.A\[15\] 0
C16360 _0554_/a_68_297# _0554_/a_150_297# 0.00477f
C16361 net237 hold90/a_391_47# 0.13409f
C16362 _0267_ _0345_ 0.03104f
C16363 hold68/a_285_47# _0758_/a_215_47# 0
C16364 VPWR _1025_/a_27_47# 0.63544f
C16365 _0466_ net17 0
C16366 _1067_/a_193_47# control0.add 0
C16367 _0286_ net228 0.00208f
C16368 _0462_ _0373_ 0.02769f
C16369 net82 _0219_ 0
C16370 _0429_ _0252_ 0.08049f
C16371 _0772_/a_79_21# _0345_ 0.01115f
C16372 _0388_ _0397_ 0
C16373 clknet_1_0__leaf__0460_ net107 0.01508f
C16374 _0422_ _0281_ 0
C16375 comp0.B\[4\] _0561_/a_240_47# 0.00278f
C16376 _0251_ _0989_/a_975_413# 0.00268f
C16377 hold31/a_285_47# net178 0.0102f
C16378 _0179_ _0195_ 0.02638f
C16379 _0188_ net67 0.10992f
C16380 net105 _1015_/a_193_47# 0
C16381 net207 _1015_/a_27_47# 0
C16382 _1019_/a_27_47# _0113_ 0
C16383 _1012_/a_27_47# _0722_/a_79_21# 0.00999f
C16384 _0538_/a_149_47# clkbuf_0__0464_/a_110_47# 0
C16385 clknet_1_1__leaf__0459_ net80 0.10355f
C16386 net32 _1041_/a_1017_47# 0
C16387 _0098_ _0392_ 0.00212f
C16388 VPWR hold95/a_49_47# 0.31243f
C16389 _0985_/a_466_413# net10 0
C16390 _0515_/a_81_21# _0186_ 0
C16391 _0343_ _0388_ 0.02907f
C16392 _0217_ _1024_/a_193_47# 0
C16393 acc0.A\[9\] _0181_ 0.13176f
C16394 _0572_/a_27_297# net111 0
C16395 _1004_/a_1059_315# _0380_ 0.0119f
C16396 _1004_/a_891_413# _0350_ 0.04995f
C16397 _0693_/a_68_297# _0352_ 0.00188f
C16398 _0717_/a_80_21# _0348_ 0.07761f
C16399 clknet_1_0__leaf__0462_ output50/a_27_47# 0.00148f
C16400 clknet_1_0__leaf__0459_ _0347_ 0.04071f
C16401 _0997_/a_1059_315# _0997_/a_891_413# 0.31086f
C16402 _0997_/a_193_47# _0997_/a_975_413# 0
C16403 _0997_/a_466_413# _0997_/a_381_47# 0.03733f
C16404 _1049_/a_27_47# net10 0
C16405 _0640_/a_109_53# _0465_ 0.00231f
C16406 hold56/a_391_47# VPWR 0.18816f
C16407 _0081_ acc0.A\[15\] 0.00113f
C16408 net78 _0287_ 0
C16409 _0181_ _0986_/a_592_47# 0
C16410 net18 _1042_/a_27_47# 0.02147f
C16411 net198 _1042_/a_193_47# 0.02699f
C16412 _0372_ _0240_ 0
C16413 hold36/a_285_47# net132 0
C16414 _0534_/a_81_21# net157 0
C16415 _0348_ _0339_ 0.00777f
C16416 _0372_ _0369_ 0.2945f
C16417 VPWR _1051_/a_561_413# 0.00302f
C16418 _0349_ _1010_/a_193_47# 0.01605f
C16419 net26 _0213_ 0
C16420 _0569_/a_109_47# _0347_ 0
C16421 hold39/a_391_47# _0951_/a_109_93# 0
C16422 acc0.A\[12\] _0993_/a_27_47# 0
C16423 net39 _0993_/a_193_47# 0
C16424 _0278_ _0399_ 0
C16425 hold7/a_49_47# net154 0
C16426 clknet_1_0__leaf__0465_ net157 0.10081f
C16427 hold6/a_49_47# _1042_/a_891_413# 0
C16428 hold6/a_391_47# _1042_/a_466_413# 0
C16429 net197 acc0.A\[25\] 0
C16430 _0402_ _0417_ 0.13775f
C16431 _0959_/a_80_21# hold84/a_49_47# 0.01001f
C16432 _0783_/a_79_21# _0347_ 0.10802f
C16433 net36 _0497_/a_68_297# 0.01689f
C16434 _0292_ _0350_ 0
C16435 _0470_ _0474_ 0
C16436 _0463_ _0171_ 0
C16437 _0151_ acc0.A\[6\] 0
C16438 _0192_ net13 0
C16439 _0793_/a_51_297# _0408_ 0.09404f
C16440 _0283_ _0347_ 0
C16441 _0793_/a_240_47# _0405_ 0
C16442 net243 _0756_/a_285_47# 0
C16443 _1027_/a_634_159# _1027_/a_1059_315# 0
C16444 _1027_/a_27_47# _1027_/a_381_47# 0.06222f
C16445 _1027_/a_193_47# _1027_/a_891_413# 0.19489f
C16446 clknet_0__0459_ _0400_ 0
C16447 clknet_1_0__leaf__0463_ _0548_/a_51_297# 0.00151f
C16448 comp0.B\[13\] hold26/a_285_47# 0.0021f
C16449 _0197_ net170 0.02933f
C16450 _0481_ _0488_ 0.07479f
C16451 acc0.A\[15\] _0505_/a_373_47# 0
C16452 _0996_/a_466_413# net41 0
C16453 VPWR _1032_/a_634_159# 0.18525f
C16454 _1061_/a_381_47# _1061_/a_561_413# 0.00123f
C16455 _1061_/a_891_413# _1061_/a_975_413# 0.00851f
C16456 _1061_/a_27_47# net147 0.23024f
C16457 _0753_/a_381_47# _0222_ 0
C16458 _0311_ _1009_/a_27_47# 0
C16459 _0305_ _1009_/a_634_159# 0
C16460 VPWR _0824_/a_59_75# 0.21262f
C16461 net51 _0345_ 0.00349f
C16462 acc0.A\[8\] _0990_/a_561_413# 0
C16463 hold6/a_285_47# net10 0.0396f
C16464 _0581_/a_27_297# acc0.A\[18\] 0.01917f
C16465 _0143_ _0527_/a_109_47# 0
C16466 clknet_0__0457_ hold40/a_49_47# 0.00852f
C16467 hold101/a_49_47# _0442_ 0.02656f
C16468 hold101/a_285_47# _0441_ 0
C16469 net58 _0465_ 0.03705f
C16470 _0124_ net112 0.00191f
C16471 _0195_ acc0.A\[26\] 0.53574f
C16472 _0197_ _0845_/a_109_297# 0
C16473 _0984_/a_891_413# net165 0
C16474 _0341_ _1030_/a_27_47# 0
C16475 _0746_/a_299_297# _0460_ 0
C16476 _0453_ _0347_ 0
C16477 clkbuf_0__0459_/a_110_47# _0185_ 0
C16478 _0977_/a_75_212# _0489_ 0.19636f
C16479 _1032_/a_193_47# _1015_/a_1059_315# 0
C16480 _1032_/a_27_47# _1015_/a_891_413# 0
C16481 hold85/a_285_47# net33 0
C16482 _1035_/a_634_159# _1035_/a_381_47# 0
C16483 acc0.A\[2\] net58 0.18922f
C16484 _0280_ _0300_ 0
C16485 _0298_ _0410_ 0
C16486 _0212_ net26 0.02552f
C16487 _0770_/a_382_297# _0350_ 0
C16488 comp0.B\[15\] _0175_ 0
C16489 clkbuf_1_0__f__0459_/a_110_47# net166 0.00427f
C16490 _1000_/a_193_47# _0247_ 0.18004f
C16491 net145 _0816_/a_68_297# 0
C16492 _0217_ net100 0.1338f
C16493 _0331_ _0690_/a_68_297# 0
C16494 _0489_ _1069_/a_975_413# 0.00192f
C16495 acc0.A\[31\] _0339_ 0.01005f
C16496 _0559_/a_149_47# net204 0
C16497 _1013_/a_1059_315# clknet_1_1__leaf__0461_ 0
C16498 _1048_/a_193_47# acc0.A\[15\] 0
C16499 net205 net160 0
C16500 _1010_/a_193_47# _0701_/a_209_297# 0
C16501 _0764_/a_81_21# _0764_/a_384_47# 0.00138f
C16502 _0343_ net77 0.00744f
C16503 _0127_ _1029_/a_193_47# 0.00378f
C16504 acc0.A\[29\] _1029_/a_1059_315# 0.10003f
C16505 _1011_/a_27_47# _0726_/a_51_297# 0.00112f
C16506 clknet_1_0__leaf__0459_ _1016_/a_891_413# 0.00635f
C16507 _1069_/a_891_413# _0167_ 0
C16508 _1069_/a_381_47# clknet_1_0__leaf_clk 0.00231f
C16509 _1069_/a_634_159# control0.count\[0\] 0
C16510 pp[17] net209 0
C16511 _0993_/a_27_47# _0650_/a_68_297# 0
C16512 _0767_/a_59_75# clkbuf_0__0461_/a_110_47# 0
C16513 _0461_ net23 0
C16514 VPWR net2 0.28744f
C16515 _0621_/a_35_297# _0435_ 0
C16516 _1052_/a_27_47# _0524_/a_27_297# 0
C16517 _1059_/a_381_47# _0185_ 0.00695f
C16518 _0259_ _0346_ 0.52389f
C16519 _0343_ _0223_ 0.60815f
C16520 hold33/a_49_47# hold33/a_285_47# 0.22264f
C16521 hold25/a_49_47# clknet_1_0__leaf__0463_ 0
C16522 net125 _1061_/a_27_47# 0.03956f
C16523 _1039_/a_27_47# net147 0
C16524 net58 net179 0
C16525 _0157_ hold82/a_391_47# 0
C16526 _0608_/a_27_47# _0309_ 0.00464f
C16527 _0239_ _0678_/a_68_297# 0.00398f
C16528 hold64/a_285_47# _0217_ 0.01386f
C16529 _0577_/a_109_297# net150 0.0015f
C16530 _0577_/a_27_297# _0217_ 0.15404f
C16531 _0953_/a_220_297# _1061_/a_27_47# 0
C16532 _0846_/a_149_47# acc0.A\[15\] 0
C16533 _0176_ _0140_ 0
C16534 _0374_ _0103_ 0.20828f
C16535 net88 _0181_ 0.26745f
C16536 net243 _0122_ 0.00554f
C16537 _0120_ _1022_/a_891_413# 0
C16538 acc0.A\[22\] _1022_/a_975_413# 0
C16539 _0577_/a_109_47# net151 0
C16540 _0816_/a_68_297# net67 0.10124f
C16541 _0221_ _0336_ 0
C16542 _0252_ clknet_1_1__leaf__0458_ 0.01924f
C16543 _0785_/a_299_297# net66 0
C16544 clknet_1_1__leaf__0458_ _0989_/a_381_47# 0
C16545 _0538_/a_240_47# _0143_ 0.00117f
C16546 net106 _1015_/a_27_47# 0
C16547 net61 _0399_ 0.02723f
C16548 _0411_ _0668_/a_297_47# 0
C16549 hold37/a_49_47# _0464_ 0
C16550 _0524_/a_109_47# net148 0
C16551 _0673_/a_103_199# net228 0.01363f
C16552 pp[11] _0993_/a_27_47# 0
C16553 output53/a_27_47# _0124_ 0
C16554 net53 net155 0
C16555 _1065_/a_27_47# _0160_ 0
C16556 net36 hold100/a_49_47# 0
C16557 _0343_ _0986_/a_1059_315# 0.02047f
C16558 hold16/a_285_47# _0218_ 0
C16559 _0475_ _0563_/a_51_297# 0.06841f
C16560 _0504_/a_27_47# _0350_ 0
C16561 _1003_/a_193_47# net159 0
C16562 _0575_/a_109_47# acc0.A\[25\] 0
C16563 _0328_ _0318_ 0.0182f
C16564 _0550_/a_512_297# B[7] 0
C16565 _0118_ clknet_1_0__leaf__0457_ 0.03102f
C16566 _0982_/a_193_47# net36 0.03092f
C16567 net45 _1013_/a_193_47# 0.0414f
C16568 hold26/a_285_47# comp0.B\[9\] 0.07322f
C16569 _0236_ _0617_/a_68_297# 0
C16570 _0260_ _0272_ 0
C16571 _0179_ _1048_/a_193_47# 0.03702f
C16572 _0500_/a_27_47# _1048_/a_381_47# 0
C16573 VPWR _0106_ 0.50488f
C16574 _0705_/a_59_75# hold61/a_285_47# 0.00353f
C16575 net177 output51/a_27_47# 0
C16576 net203 _0175_ 0.003f
C16577 net239 clknet_1_1__leaf__0462_ 0.11131f
C16578 _0255_ _0256_ 0.07335f
C16579 net45 _0607_/a_109_297# 0.00167f
C16580 _0456_ _0350_ 0.00121f
C16581 net89 _0101_ 0.0104f
C16582 clkbuf_1_0__f__0458_/a_110_47# acc0.A\[15\] 0.01327f
C16583 net70 _0181_ 0.17702f
C16584 _0255_ _0987_/a_1059_315# 0.00141f
C16585 _0280_ _0404_ 0.02049f
C16586 _0993_/a_1059_315# _0993_/a_891_413# 0.31086f
C16587 _0993_/a_193_47# _0993_/a_975_413# 0
C16588 _0993_/a_466_413# _0993_/a_381_47# 0.03733f
C16589 _1058_/a_381_47# _0156_ 0.11467f
C16590 hold33/a_49_47# net20 0
C16591 hold48/a_391_47# comp0.B\[12\] 0.01086f
C16592 clknet_0__0463_ net247 0
C16593 hold18/a_285_47# net165 0.00793f
C16594 _1039_/a_891_413# _1039_/a_975_413# 0.00851f
C16595 _1039_/a_27_47# net125 0.22166f
C16596 _1039_/a_381_47# _1039_/a_561_413# 0.00123f
C16597 _0346_ net221 0
C16598 net185 hold84/a_391_47# 0
C16599 _0180_ _0531_/a_373_47# 0.00226f
C16600 _0199_ _0531_/a_27_297# 0.00117f
C16601 net46 clkbuf_1_0__f__0461_/a_110_47# 0.01225f
C16602 net187 net1 0
C16603 net178 output47/a_27_47# 0
C16604 _0663_/a_297_47# _0287_ 0
C16605 _0663_/a_207_413# _0293_ 0
C16606 _0580_/a_27_297# _0580_/a_109_297# 0.17136f
C16607 output56/a_27_47# _0333_ 0
C16608 _0996_/a_1059_315# _0400_ 0
C16609 net7 clknet_1_1__leaf__0457_ 0.04098f
C16610 _1032_/a_891_413# _0215_ 0.00272f
C16611 _0179_ _0846_/a_149_47# 0.02771f
C16612 _0465_ _0262_ 0.00296f
C16613 _1026_/a_466_413# _1026_/a_592_47# 0.00553f
C16614 _1026_/a_634_159# _1026_/a_1017_47# 0
C16615 _1059_/a_27_47# VPWR 0.63769f
C16616 _0361_ _0360_ 0.13841f
C16617 _0985_/a_193_47# _0449_ 0.0025f
C16618 clknet_1_0__leaf__0461_ hold93/a_285_47# 0.01917f
C16619 _0985_/a_1017_47# clknet_1_0__leaf__0458_ 0
C16620 _0752_/a_300_297# _0103_ 0
C16621 net36 _0450_ 0
C16622 hold10/a_285_47# _0472_ 0
C16623 _0473_ _1061_/a_27_47# 0
C16624 _0697_/a_80_21# _0324_ 0.1384f
C16625 net36 comp0.B\[8\] 0
C16626 net140 net139 0.0042f
C16627 _0476_ clknet_0_clk 0
C16628 acc0.A\[2\] _0262_ 0.19533f
C16629 _0718_/a_47_47# _0348_ 0.37574f
C16630 _0181_ _1009_/a_634_159# 0.00168f
C16631 _0095_ net41 0.04406f
C16632 _0695_/a_217_297# _0324_ 0.04094f
C16633 _1024_/a_466_413# acc0.A\[24\] 0
C16634 _1024_/a_381_47# _0122_ 0.13795f
C16635 _0313_ net54 0.09569f
C16636 _0355_ acc0.A\[28\] 0
C16637 hold27/a_285_47# _0913_/a_27_47# 0
C16638 net51 net52 0
C16639 _0119_ _1020_/a_193_47# 0
C16640 hold66/a_49_47# hold66/a_391_47# 0.00188f
C16641 _0527_/a_27_297# _0186_ 0.15206f
C16642 _0121_ net176 0
C16643 _0376_ _0223_ 0.00314f
C16644 _0642_/a_27_413# _0437_ 0
C16645 _0662_/a_81_21# _0662_/a_299_297# 0.08213f
C16646 _0343_ _0854_/a_297_297# 0
C16647 hold75/a_285_47# _0347_ 0
C16648 _1057_/a_891_413# net143 0
C16649 net33 _0132_ 0
C16650 _1037_/a_27_47# _1037_/a_634_159# 0.14145f
C16651 pp[16] _0997_/a_1059_315# 0
C16652 _0276_ net5 0
C16653 hold4/a_49_47# hold4/a_285_47# 0.22264f
C16654 acc0.A\[22\] _0756_/a_47_47# 0.0021f
C16655 comp0.B\[10\] _1040_/a_193_47# 0.00584f
C16656 acc0.A\[3\] hold71/a_391_47# 0
C16657 _0972_/a_93_21# _0951_/a_109_93# 0
C16658 hold48/a_49_47# net20 0
C16659 _0186_ _0989_/a_634_159# 0
C16660 hold1/a_391_47# _0186_ 0
C16661 net159 _0471_ 0
C16662 _0957_/a_304_297# net24 0.00153f
C16663 hold48/a_49_47# hold48/a_285_47# 0.22264f
C16664 _0988_/a_1059_315# net142 0
C16665 _0785_/a_81_21# _0423_ 0
C16666 clkbuf_1_0__f__0458_/a_110_47# _0179_ 0.16039f
C16667 net242 net239 0.00255f
C16668 control0.state\[1\] _1067_/a_193_47# 0
C16669 net158 _0142_ 0
C16670 _1068_/a_1017_47# _0468_ 0
C16671 _0790_/a_35_297# _0790_/a_285_47# 0.00723f
C16672 _0538_/a_512_297# _0473_ 0.00128f
C16673 _1041_/a_634_159# _1041_/a_381_47# 0
C16674 _0343_ _1013_/a_1017_47# 0
C16675 _1048_/a_1059_315# clknet_1_1__leaf__0457_ 0
C16676 net121 net24 0
C16677 VPWR _0991_/a_1059_315# 0.4675f
C16678 hold99/a_391_47# _0993_/a_1059_315# 0.01554f
C16679 _0663_/a_27_413# clknet_1_1__leaf__0465_ 0
C16680 _0389_ _0769_/a_81_21# 0.11464f
C16681 VPWR _0496_/a_27_47# 0.2233f
C16682 net166 clkbuf_0__0461_/a_110_47# 0
C16683 _1015_/a_592_47# comp0.B\[15\] 0
C16684 hold89/a_285_47# clknet_0_clk 0
C16685 net146 _0219_ 0.37972f
C16686 _0342_ net60 0
C16687 net106 _0215_ 0
C16688 _1002_/a_891_413# net1 0.02088f
C16689 _0415_ _0345_ 0
C16690 _0409_ net42 0
C16691 _0176_ _1043_/a_634_159# 0
C16692 net201 _0560_/a_68_297# 0
C16693 _1039_/a_27_47# _0473_ 0.03f
C16694 _0569_/a_27_297# acc0.A\[28\] 0.01396f
C16695 _0428_ _0186_ 0
C16696 acc0.A\[29\] _0723_/a_297_47# 0.00155f
C16697 _0274_ _0447_ 0
C16698 comp0.B\[1\] _0113_ 0.05171f
C16699 _1051_/a_27_47# _0193_ 0
C16700 _0707_/a_315_47# _0333_ 0.0107f
C16701 net202 _0584_/a_27_297# 0
C16702 clkbuf_1_1__f__0458_/a_110_47# acc0.A\[6\] 0.02795f
C16703 _0399_ _0812_/a_215_47# 0
C16704 _0741_/a_109_297# acc0.A\[24\] 0.00181f
C16705 net232 hold84/a_49_47# 0
C16706 VPWR _1011_/a_27_47# 0.48688f
C16707 _0195_ _0530_/a_384_47# 0
C16708 _0234_ _0762_/a_79_21# 0.01593f
C16709 _0476_ _0955_/a_220_297# 0
C16710 _0445_ _0084_ 0
C16711 _0266_ _0269_ 0
C16712 _0251_ _0254_ 0.10623f
C16713 clknet_0__0459_ clkbuf_0__0459_/a_110_47# 1.69985f
C16714 _0640_/a_109_53# _0254_ 0
C16715 net65 _0253_ 0.0322f
C16716 _0357_ clknet_1_1__leaf__0462_ 0.01834f
C16717 input2/a_75_212# _0515_/a_299_297# 0.00154f
C16718 _0661_/a_205_297# net67 0
C16719 _1019_/a_27_47# _0345_ 0.44913f
C16720 _0985_/a_27_47# _0846_/a_51_297# 0
C16721 _0574_/a_27_297# net50 0.0054f
C16722 hold69/a_285_47# _0370_ 0
C16723 _0343_ pp[27] 0.0337f
C16724 _0743_/a_240_47# _0359_ 0.00486f
C16725 _1012_/a_193_47# _0110_ 0.2288f
C16726 net183 clknet_0__0464_ 0.00332f
C16727 _0713_/a_27_47# net105 0.03509f
C16728 net89 net35 0.07608f
C16729 clknet_1_1__leaf__0460_ _0195_ 0.02354f
C16730 clkbuf_1_0__f__0457_/a_110_47# net118 0
C16731 _0108_ _0318_ 0
C16732 clknet_1_1__leaf__0460_ net92 0
C16733 _0083_ net10 0
C16734 hold27/a_285_47# _0172_ 0.06923f
C16735 _0124_ net111 0.04468f
C16736 _0216_ _0570_/a_373_47# 0
C16737 _0578_/a_27_297# VPWR 0.28448f
C16738 _0644_/a_377_297# VPWR 0.00418f
C16739 _0567_/a_109_297# net209 0
C16740 _0579_/a_27_297# _0352_ 0
C16741 _0740_/a_113_47# _0219_ 0
C16742 _0324_ _0345_ 0.02272f
C16743 hold99/a_285_47# hold99/a_391_47# 0.41909f
C16744 VPWR _1044_/a_975_413# 0.00477f
C16745 _0146_ _1049_/a_27_47# 0
C16746 clknet_1_0__leaf__0464_ net154 0.00408f
C16747 _0519_/a_299_297# _0436_ 0
C16748 _0152_ _0828_/a_113_297# 0
C16749 VPWR _0425_ 0.42399f
C16750 _0161_ hold84/a_285_47# 0.00102f
C16751 _0314_ VPWR 0.2648f
C16752 net58 _0254_ 0.1161f
C16753 hold35/a_49_47# _0189_ 0.0062f
C16754 hold35/a_391_47# net2 0
C16755 _0316_ _0697_/a_80_21# 0
C16756 _0631_/a_109_297# _0263_ 0.01129f
C16757 clkload4/a_268_47# clkload4/Y 0.00587f
C16758 _0398_ _0352_ 0.0254f
C16759 _0316_ net56 0
C16760 _0756_/a_47_47# _0379_ 0.14637f
C16761 _0756_/a_285_47# _0378_ 0.06696f
C16762 _0684_/a_59_75# _0323_ 0
C16763 _1001_/a_975_413# _0461_ 0
C16764 clkbuf_1_1__f__0465_/a_110_47# net217 0.01201f
C16765 _0983_/a_634_159# _0264_ 0
C16766 _1027_/a_466_413# net156 0.00296f
C16767 _0643_/a_103_199# _0272_ 0.113f
C16768 net44 _0341_ 0.00372f
C16769 _0606_/a_215_297# _0377_ 0
C16770 _0606_/a_297_297# _0345_ 0.00124f
C16771 _0181_ _1067_/a_891_413# 0.00483f
C16772 net141 net47 0.17909f
C16773 _1030_/a_466_413# _0707_/a_75_199# 0
C16774 net239 hold92/a_49_47# 0
C16775 VPWR _0528_/a_384_47# 0
C16776 comp0.B\[2\] _0560_/a_68_297# 0.17282f
C16777 clknet_1_0__leaf__0465_ net13 0.18184f
C16778 _0710_/a_109_47# VPWR 0
C16779 net61 _0619_/a_68_297# 0
C16780 clknet_0__0465_ _0840_/a_68_297# 0.00132f
C16781 clknet_1_0__leaf__0462_ _1023_/a_381_47# 0.00124f
C16782 net204 comp0.B\[5\] 0.03341f
C16783 net56 _0347_ 0
C16784 _0116_ acc0.A\[18\] 0.30224f
C16785 clknet_1_0__leaf__0464_ _0465_ 0.00619f
C16786 _0131_ comp0.B\[6\] 0
C16787 _0582_/a_27_297# _0582_/a_109_297# 0.17136f
C16788 _0751_/a_111_297# _0225_ 0.0024f
C16789 net133 _1061_/a_1059_315# 0
C16790 clknet_1_0__leaf__0464_ _1061_/a_381_47# 0
C16791 _0757_/a_150_297# net50 0
C16792 _0343_ net83 0.00768f
C16793 net176 _0380_ 0.00393f
C16794 _0678_/a_68_297# _0309_ 0.12275f
C16795 _1052_/a_27_47# _1052_/a_466_413# 0.25987f
C16796 _1052_/a_193_47# _1052_/a_634_159# 0.11072f
C16797 net202 _1015_/a_634_159# 0
C16798 _0478_ _1071_/a_193_47# 0.00162f
C16799 _1007_/a_27_47# _1007_/a_193_47# 0.96985f
C16800 _0125_ net197 0.08117f
C16801 _1035_/a_891_413# _0133_ 0.05682f
C16802 _1035_/a_381_47# net121 0.00201f
C16803 _1012_/a_193_47# _1010_/a_193_47# 0
C16804 _0497_/a_68_297# _1061_/a_27_47# 0
C16805 hold87/a_49_47# _0266_ 0
C16806 _1012_/a_27_47# acc0.A\[30\] 0
C16807 _0357_ net242 0
C16808 _1058_/a_27_47# _1058_/a_891_413# 0.03224f
C16809 _1058_/a_193_47# _1058_/a_1059_315# 0.03405f
C16810 _1058_/a_634_159# _1058_/a_466_413# 0.23992f
C16811 net139 input14/a_75_212# 0.00183f
C16812 clkload4/a_110_47# _0459_ 0
C16813 B[15] net23 0.00264f
C16814 hold69/a_391_47# _0350_ 0.04221f
C16815 hold10/a_391_47# _0499_/a_59_75# 0
C16816 _0343_ _0781_/a_68_297# 0.00427f
C16817 hold14/a_49_47# B[1] 0
C16818 _0747_/a_79_21# clknet_1_0__leaf__0460_ 0
C16819 _1051_/a_381_47# _0172_ 0.02688f
C16820 _0110_ clknet_1_1__leaf__0461_ 0
C16821 _0353_ _0723_/a_27_413# 0.00142f
C16822 VPWR _0180_ 2.51112f
C16823 _0558_/a_68_297# _1035_/a_891_413# 0.00141f
C16824 VPWR net218 0.18292f
C16825 _1050_/a_634_159# _0527_/a_27_297# 0
C16826 _1050_/a_193_47# _0527_/a_109_297# 0
C16827 _0356_ acc0.A\[29\] 0.02589f
C16828 _0399_ _0431_ 0
C16829 _0310_ _0780_/a_285_47# 0
C16830 _0176_ _0175_ 0.01669f
C16831 VPWR net152 0.24627f
C16832 _0718_/a_377_297# _0349_ 0.00188f
C16833 _0718_/a_285_47# _0337_ 0.03978f
C16834 _1011_/a_193_47# net227 0
C16835 _1011_/a_466_413# _0354_ 0.01228f
C16836 _1011_/a_634_159# _0355_ 0.0238f
C16837 _0462_ _0773_/a_117_297# 0
C16838 VPWR _1013_/a_193_47# 0.29863f
C16839 net182 net2 0.00181f
C16840 _0626_/a_68_297# _0218_ 0
C16841 clknet_1_0__leaf_clk control0.count\[0\] 0.37093f
C16842 _1033_/a_381_47# _1065_/a_1059_315# 0
C16843 _0983_/a_193_47# clknet_1_0__leaf__0458_ 0.00199f
C16844 _0607_/a_109_297# VPWR 0.19046f
C16845 _0399_ _0659_/a_68_297# 0
C16846 _1052_/a_891_413# net148 0.0026f
C16847 _1052_/a_27_47# _0194_ 0.00126f
C16848 _0258_ _0186_ 0.02803f
C16849 net117 _0568_/a_27_297# 0
C16850 _0642_/a_298_297# _0434_ 0
C16851 _0328_ _1007_/a_27_47# 0
C16852 _0812_/a_79_21# _0345_ 0.00312f
C16853 _0477_ _1065_/a_193_47# 0
C16854 _0432_ VPWR 0.72619f
C16855 net21 B[12] 0.0052f
C16856 acc0.A\[9\] _0990_/a_193_47# 0
C16857 net149 hold60/a_49_47# 0
C16858 _0310_ _0677_/a_47_47# 0
C16859 _0217_ _0120_ 0.37718f
C16860 _0953_/a_32_297# net147 0.01657f
C16861 comp0.B\[10\] _1061_/a_1059_315# 0
C16862 _0195_ _1018_/a_561_413# 0.00124f
C16863 net156 _1026_/a_381_47# 0
C16864 _1027_/a_466_413# acc0.A\[26\] 0
C16865 net65 output61/a_27_47# 0.02129f
C16866 _0346_ _0772_/a_215_47# 0
C16867 hold68/a_49_47# _0380_ 0
C16868 net58 _0988_/a_561_413# 0
C16869 _0136_ _0549_/a_68_297# 0
C16870 _0467_ _1067_/a_975_413# 0
C16871 _0297_ _0400_ 0
C16872 _0195_ _1049_/a_891_413# 0.00112f
C16873 pp[30] _0708_/a_68_297# 0
C16874 _0786_/a_80_21# _0786_/a_217_297# 0.12661f
C16875 _0685_/a_68_297# _0685_/a_150_297# 0.00477f
C16876 _1038_/a_1059_315# _0176_ 0.00218f
C16877 _0343_ _0216_ 0.06417f
C16878 _1021_/a_27_47# acc0.A\[20\] 0
C16879 _1039_/a_27_47# _0497_/a_68_297# 0.01167f
C16880 hold59/a_49_47# _0116_ 0
C16881 net205 _1034_/a_193_47# 0
C16882 net33 net25 0
C16883 _0985_/a_193_47# _0260_ 0
C16884 net59 _1012_/a_1059_315# 0.08631f
C16885 _0994_/a_193_47# _0218_ 0.03964f
C16886 _0403_ _0993_/a_466_413# 0
C16887 comp0.B\[12\] net195 0.01295f
C16888 comp0.B\[11\] net19 0.08529f
C16889 net67 _0806_/a_113_297# 0
C16890 _0995_/a_1059_315# pp[14] 0.02522f
C16891 hold13/a_285_47# _1039_/a_27_47# 0
C16892 _0579_/a_109_297# net105 0
C16893 _0413_ _0405_ 0
C16894 _0412_ _0400_ 0
C16895 _0137_ B[7] 0
C16896 _0798_/a_113_297# _0219_ 0.00173f
C16897 _0538_/a_240_47# _0174_ 0.01466f
C16898 VPWR _1042_/a_466_413# 0.24345f
C16899 _1056_/a_193_47# acc0.A\[9\] 0.01502f
C16900 _0982_/a_27_47# _0346_ 0.03225f
C16901 output35/a_27_47# done 0.15955f
C16902 _0316_ _0345_ 0
C16903 _0518_/a_27_297# acc0.A\[7\] 0
C16904 _1043_/a_1059_315# _1042_/a_381_47# 0
C16905 _1043_/a_381_47# _1042_/a_1059_315# 0
C16906 clknet_1_1__leaf__0464_ net198 0.02465f
C16907 _1030_/a_27_47# acc0.A\[30\] 0.1535f
C16908 _1030_/a_381_47# _0704_/a_68_297# 0.00136f
C16909 _0477_ net33 0
C16910 net105 _0399_ 0.10634f
C16911 _0642_/a_27_413# _0252_ 0.0906f
C16912 hold89/a_49_47# _0488_ 0
C16913 _0988_/a_27_47# _0988_/a_1059_315# 0.04875f
C16914 _0988_/a_193_47# _0988_/a_466_413# 0.07855f
C16915 clkbuf_1_1__f__0465_/a_110_47# net66 0.00503f
C16916 control0.reset _0173_ 0.09274f
C16917 net232 _0471_ 0
C16918 _1039_/a_634_159# _0174_ 0
C16919 _0352_ _0754_/a_240_47# 0
C16920 _0814_/a_27_47# _0347_ 0
C16921 _0347_ _0345_ 0.14718f
C16922 _0984_/a_891_413# _0983_/a_27_47# 0
C16923 _0869_/a_27_47# net47 0
C16924 _0998_/a_193_47# _0781_/a_68_297# 0.00156f
C16925 _0388_ clkbuf_0__0461_/a_110_47# 0
C16926 _0730_/a_79_21# _0358_ 0.20617f
C16927 _0183_ acc0.A\[15\] 0.10145f
C16928 comp0.B\[14\] _1040_/a_1059_315# 0
C16929 acc0.A\[17\] _0240_ 0.0542f
C16930 _0580_/a_109_297# _0117_ 0.00413f
C16931 _0324_ net52 0.17248f
C16932 net63 _0836_/a_68_297# 0.02166f
C16933 hold20/a_391_47# _0490_ 0
C16934 _0953_/a_32_297# _0953_/a_220_297# 0.00132f
C16935 hold20/a_285_47# net167 0.00974f
C16936 acc0.A\[17\] _0369_ 0.02729f
C16937 hold28/a_49_47# _0465_ 0
C16938 _0367_ _0319_ 0
C16939 hold21/a_391_47# hold22/a_391_47# 0
C16940 _0542_/a_51_297# _0542_/a_240_47# 0.03076f
C16941 net63 net212 0.00353f
C16942 _0346_ net238 0.00763f
C16943 hold96/a_285_47# _0575_/a_27_297# 0
C16944 hold96/a_49_47# _0575_/a_109_297# 0
C16945 _0162_ _1064_/a_891_413# 0.00172f
C16946 _0485_ _1064_/a_975_413# 0
C16947 _0559_/a_51_297# clknet_1_1__leaf__0463_ 0.0019f
C16948 hold52/a_391_47# net200 0
C16949 _1026_/a_381_47# acc0.A\[26\] 0
C16950 hold94/a_391_47# net51 0
C16951 _1001_/a_27_47# clknet_1_0__leaf__0457_ 0.01435f
C16952 acc0.A\[2\] hold28/a_49_47# 0.29357f
C16953 _0465_ _1047_/a_592_47# 0
C16954 net77 _0842_/a_59_75# 0
C16955 _0999_/a_193_47# _0396_ 0.00106f
C16956 _0472_ _1061_/a_592_47# 0
C16957 _0346_ _0446_ 0
C16958 clknet_1_1__leaf__0460_ _1009_/a_381_47# 0.00682f
C16959 _0817_/a_266_297# _0424_ 0.01101f
C16960 _0242_ _0771_/a_382_47# 0
C16961 net56 hold95/a_49_47# 0.34754f
C16962 acc0.A\[3\] _0845_/a_109_47# 0
C16963 _1035_/a_27_47# net27 0.01157f
C16964 _0853_/a_68_297# _0218_ 0.18675f
C16965 _0981_/a_109_47# _0484_ 0
C16966 clknet_1_1__leaf__0458_ _0988_/a_891_413# 0
C16967 net46 _0616_/a_78_199# 0.068f
C16968 _0122_ acc0.A\[24\] 0
C16969 net19 _0202_ 0.00116f
C16970 _0141_ _0540_/a_240_47# 0
C16971 _0203_ net20 0.0478f
C16972 net15 _0437_ 0
C16973 _0982_/a_466_413# hold60/a_49_47# 0.00133f
C16974 _0982_/a_193_47# hold60/a_391_47# 0
C16975 _0982_/a_634_159# hold60/a_285_47# 0
C16976 _0787_/a_209_297# _0787_/a_209_47# 0
C16977 _0787_/a_80_21# _0787_/a_303_47# 0.01146f
C16978 hold47/a_391_47# net154 0
C16979 _0461_ _0614_/a_183_297# 0
C16980 _0230_ net241 0.06894f
C16981 _0226_ _0219_ 0.49971f
C16982 _0792_/a_209_297# _0345_ 0.00749f
C16983 _0252_ _0218_ 0
C16984 _0174_ _1040_/a_1017_47# 0
C16985 _1037_/a_891_413# _1037_/a_975_413# 0.00851f
C16986 _1037_/a_381_47# _1037_/a_561_413# 0.00123f
C16987 A[8] net12 0
C16988 _0218_ _0989_/a_381_47# 0
C16989 _0997_/a_634_159# _0218_ 0.00109f
C16990 VPWR hold70/a_285_47# 0.27585f
C16991 _0195_ _0998_/a_466_413# 0.02348f
C16992 clkbuf_1_1__f__0465_/a_110_47# _0350_ 0
C16993 _0369_ net5 0.02158f
C16994 net231 _0951_/a_109_93# 0.02804f
C16995 _0255_ clknet_0__0465_ 0.09575f
C16996 pp[30] _1030_/a_634_159# 0.00803f
C16997 net59 _1030_/a_1059_315# 0
C16998 comp0.B\[8\] _1061_/a_27_47# 0
C16999 _0708_/a_68_297# _0339_ 0.00114f
C17000 VPWR _1005_/a_975_413# 0.00546f
C17001 _0463_ _0494_/a_27_47# 0.00488f
C17002 hold89/a_49_47# _1064_/a_27_47# 0
C17003 _0143_ _0473_ 0.00135f
C17004 _0629_/a_59_75# _0446_ 0
C17005 _0428_ net62 0.00153f
C17006 _0985_/a_891_413# _0844_/a_297_47# 0
C17007 net54 _0321_ 0.00259f
C17008 _1054_/a_1017_47# _0180_ 0.00208f
C17009 _0183_ _0179_ 0
C17010 pp[7] VPWR 0.57512f
C17011 _0251_ _0625_/a_59_75# 0
C17012 _1001_/a_193_47# _1001_/a_466_413# 0.07593f
C17013 _1001_/a_27_47# _1001_/a_1059_315# 0.04875f
C17014 net49 clknet_1_0__leaf__0460_ 0.16653f
C17015 clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ 1.65028f
C17016 _0621_/a_285_297# acc0.A\[6\] 0.0114f
C17017 _0343_ _0825_/a_68_297# 0
C17018 net233 _0843_/a_150_297# 0
C17019 hold76/a_49_47# net223 0
C17020 _0176_ net129 0.06276f
C17021 _1062_/a_27_47# _1062_/a_634_159# 0.14145f
C17022 _0717_/a_303_47# _0333_ 0.0041f
C17023 _0399_ _0269_ 0
C17024 _0239_ _0677_/a_47_47# 0.02327f
C17025 _0183_ hold40/a_285_47# 0.00719f
C17026 _0670_/a_79_21# clkbuf_1_1__f__0459_/a_110_47# 0
C17027 net81 acc0.A\[13\] 0
C17028 _0143_ clkbuf_1_1__f__0464_/a_110_47# 0
C17029 _0127_ acc0.A\[28\] 0
C17030 _0473_ _0953_/a_32_297# 0.03512f
C17031 hold38/a_285_47# _0951_/a_109_93# 0
C17032 net137 net13 0
C17033 _0831_/a_35_297# _0831_/a_285_47# 0.00723f
C17034 output44/a_27_47# _0195_ 0
C17035 _0575_/a_27_297# _1024_/a_27_47# 0.00892f
C17036 _0963_/a_117_297# _0489_ 0.00181f
C17037 net35 clkbuf_0_clk/a_110_47# 0.00248f
C17038 _0822_/a_109_297# _0255_ 0
C17039 clknet_1_1__leaf__0459_ _0195_ 0.17598f
C17040 _0146_ _0531_/a_109_47# 0
C17041 acc0.A\[21\] hold94/a_49_47# 0
C17042 _0459_ clknet_1_0__leaf__0457_ 0.00343f
C17043 _1049_/a_891_413# _1048_/a_193_47# 0.00726f
C17044 _1049_/a_1059_315# _1048_/a_634_159# 0
C17045 _0758_/a_79_21# acc0.A\[23\] 0.01956f
C17046 clknet_1_0__leaf__0464_ clknet_0__0464_ 0.08112f
C17047 _1058_/a_193_47# pp[10] 0
C17048 net248 _0828_/a_113_297# 0
C17049 hold14/a_285_47# _1037_/a_193_47# 0
C17050 hold14/a_49_47# _1037_/a_634_159# 0
C17051 hold14/a_391_47# _1037_/a_27_47# 0
C17052 _0572_/a_27_297# VPWR 0.27472f
C17053 net45 net59 0
C17054 _0967_/a_109_93# hold84/a_391_47# 0
C17055 VPWR _1006_/a_381_47# 0.07567f
C17056 clkbuf_0__0465_/a_110_47# _0345_ 0
C17057 _0278_ _0346_ 0
C17058 _0222_ hold29/a_285_47# 0
C17059 _0546_/a_51_297# _0545_/a_68_297# 0
C17060 _1000_/a_193_47# _0217_ 0
C17061 hold43/a_49_47# _1029_/a_27_47# 0
C17062 clkload1/Y _0271_ 0
C17063 net194 _0538_/a_149_47# 0
C17064 acc0.A\[5\] _0835_/a_215_47# 0
C17065 _0143_ _0186_ 0
C17066 _0195_ _1030_/a_975_413# 0
C17067 _0216_ _1030_/a_381_47# 0
C17068 _0346_ _0245_ 0
C17069 net48 _1005_/a_975_413# 0
C17070 VPWR _0986_/a_381_47# 0.07545f
C17071 _1039_/a_27_47# comp0.B\[8\] 0
C17072 _0715_/a_27_47# net62 0.16873f
C17073 _0714_/a_512_297# _0219_ 0
C17074 pp[9] _1058_/a_1059_315# 0
C17075 _0694_/a_113_47# _0219_ 0
C17076 VPWR _0495_/a_150_297# 0.00191f
C17077 _1070_/a_27_47# _0978_/a_27_297# 0
C17078 hold55/a_285_47# _0891_/a_27_47# 0
C17079 _1031_/a_27_47# net209 0
C17080 _1031_/a_381_47# hold62/a_285_47# 0
C17081 _0701_/a_303_47# _0332_ 0
C17082 _0186_ _0988_/a_193_47# 0
C17083 net34 rst 0.00326f
C17084 _1004_/a_466_413# _0216_ 0.01921f
C17085 _0179_ acc0.A\[15\] 0.07071f
C17086 net126 pp[0] 0
C17087 hold78/a_285_47# _0714_/a_51_297# 0
C17088 _0225_ _0103_ 0.00541f
C17089 _0561_/a_51_297# _0561_/a_512_297# 0.0116f
C17090 VPWR _0616_/a_292_297# 0.00977f
C17091 _0157_ clknet_1_1__leaf__0465_ 0.17656f
C17092 _0195_ _0171_ 0
C17093 _1072_/a_27_47# _1068_/a_1059_315# 0
C17094 _1072_/a_466_413# _1068_/a_193_47# 0
C17095 _1072_/a_193_47# _1068_/a_466_413# 0.00177f
C17096 _0476_ _1065_/a_27_47# 0
C17097 _0345_ hold95/a_49_47# 0.00123f
C17098 _0515_/a_81_21# _0514_/a_109_297# 0
C17099 _0515_/a_299_297# _0514_/a_27_297# 0
C17100 _0464_ _0463_ 0
C17101 _0198_ _0147_ 0
C17102 _0347_ net52 0.10373f
C17103 pp[0] input8/a_75_212# 0.00281f
C17104 comp0.B\[13\] _0538_/a_240_47# 0.00428f
C17105 _1001_/a_1059_315# _0459_ 0
C17106 _0317_ clkbuf_1_1__f__0460_/a_110_47# 0.0407f
C17107 _0287_ _0288_ 0.13792f
C17108 _0738_/a_68_297# _0738_/a_150_297# 0.00477f
C17109 _1003_/a_975_413# acc0.A\[21\] 0
C17110 acc0.A\[12\] _0716_/a_27_47# 0.01464f
C17111 _0265_ clknet_1_0__leaf__0457_ 0
C17112 output67/a_27_47# _0186_ 0
C17113 _0538_/a_51_297# _1046_/a_891_413# 0
C17114 net59 _0587_/a_27_47# 0
C17115 _0461_ _0391_ 0.00216f
C17116 _1035_/a_891_413# _0208_ 0
C17117 net69 _0264_ 0
C17118 _0274_ _0275_ 0.11396f
C17119 hold87/a_49_47# _0399_ 0.0127f
C17120 _1047_/a_634_159# _1047_/a_1059_315# 0
C17121 _1047_/a_27_47# _1047_/a_381_47# 0.06222f
C17122 _1047_/a_193_47# _1047_/a_891_413# 0.19489f
C17123 net47 _1060_/a_193_47# 0
C17124 _1030_/a_634_159# _0339_ 0.01332f
C17125 _1030_/a_1059_315# _0335_ 0
C17126 _0547_/a_68_297# net174 0
C17127 _0206_ _1040_/a_561_413# 0.00204f
C17128 hold97/a_391_47# _0330_ 0
C17129 _0504_/a_27_47# _1014_/a_27_47# 0
C17130 _0957_/a_220_297# _0472_ 0.00864f
C17131 hold1/a_49_47# _0987_/a_1059_315# 0.01071f
C17132 _0401_ _0673_/a_103_199# 0.00109f
C17133 net83 _0793_/a_51_297# 0.00754f
C17134 _0957_/a_114_297# _0475_ 0.00172f
C17135 _0104_ net52 0
C17136 _0331_ _0365_ 0.00523f
C17137 net46 _0384_ 0
C17138 clknet_1_0__leaf__0462_ acc0.A\[23\] 0.05707f
C17139 _0664_/a_79_21# _0285_ 0.20409f
C17140 _1041_/a_891_413# _0174_ 0.02152f
C17141 hold5/a_391_47# hold51/a_285_47# 0
C17142 net245 net81 0.02439f
C17143 _0133_ _0473_ 0
C17144 _0582_/a_109_297# _0115_ 0.00169f
C17145 net234 _1014_/a_466_413# 0
C17146 _0456_ _1014_/a_27_47# 0
C17147 _0797_/a_207_413# acc0.A\[13\] 0.00172f
C17148 net178 _0517_/a_384_47# 0.01006f
C17149 _1007_/a_466_413# _1007_/a_592_47# 0.00553f
C17150 _1007_/a_634_159# _1007_/a_1017_47# 0
C17151 _1052_/a_1059_315# _1052_/a_1017_47# 0
C17152 _1001_/a_891_413# clknet_1_0__leaf__0461_ 0
C17153 _0180_ _0523_/a_81_21# 0
C17154 hold96/a_391_47# _1004_/a_466_413# 0.00868f
C17155 VPWR _0360_ 0.41049f
C17156 _1012_/a_27_47# net96 0
C17157 VPWR _0854_/a_510_47# 0
C17158 _0525_/a_81_21# _0522_/a_27_297# 0
C17159 net240 hold93/a_285_47# 0.02563f
C17160 _0837_/a_266_47# _0837_/a_585_47# 0.0013f
C17161 _1058_/a_466_413# net144 0
C17162 _0172_ _1044_/a_561_413# 0.00163f
C17163 _0179_ _1052_/a_561_413# 0.00226f
C17164 _0502_/a_27_47# _0533_/a_109_297# 0
C17165 net185 _0957_/a_32_297# 0
C17166 _1020_/a_1059_315# _0352_ 0.03913f
C17167 net190 _1027_/a_27_47# 0
C17168 _1021_/a_27_47# net107 0.22772f
C17169 _1021_/a_634_159# clknet_1_0__leaf__0461_ 0
C17170 A[8] pp[5] 0.16337f
C17171 VPWR _0498_/a_51_297# 0.4682f
C17172 acc0.A\[5\] _0172_ 0.47481f
C17173 _0986_/a_27_47# _0840_/a_68_297# 0
C17174 _0557_/a_245_297# VPWR 0.00505f
C17175 net248 _0433_ 0.07236f
C17176 _0219_ net41 0.29155f
C17177 _0731_/a_81_21# _0462_ 0.00168f
C17178 pp[9] net47 0
C17179 _0258_ net62 0.06393f
C17180 hold74/a_285_47# _0305_ 0.00861f
C17181 _0635_/a_27_47# _0265_ 0.03921f
C17182 net185 net23 0
C17183 net61 _0346_ 0.0276f
C17184 _1003_/a_466_413# _0487_ 0
C17185 control0.state\[0\] _0951_/a_209_311# 0
C17186 control0.state\[1\] _0951_/a_109_93# 0.14593f
C17187 _0669_/a_111_297# net41 0
C17188 _1011_/a_592_47# _0109_ 0.00188f
C17189 net97 _0355_ 0
C17190 _0216_ _0726_/a_512_297# 0
C17191 _1018_/a_193_47# _0580_/a_109_297# 0
C17192 _1033_/a_1059_315# control0.reset 0
C17193 _1002_/a_1017_47# VPWR 0
C17194 net40 net6 0.16866f
C17195 hold21/a_391_47# A[7] 0
C17196 _1061_/a_634_159# comp0.B\[9\] 0
C17197 _0139_ net196 0
C17198 net61 net65 0.31109f
C17199 clkbuf_0_clk/a_110_47# _1063_/a_466_413# 0
C17200 net61 _0989_/a_466_413# 0
C17201 _1000_/a_27_47# _0372_ 0
C17202 _0924_/a_27_47# net8 0
C17203 hold59/a_285_47# _0350_ 0
C17204 _0243_ _0616_/a_493_297# 0
C17205 clkbuf_1_0__f__0462_/a_110_47# hold90/a_391_47# 0.00514f
C17206 hold75/a_391_47# net222 0.13101f
C17207 hold40/a_49_47# hold40/a_391_47# 0.00188f
C17208 _0983_/a_193_47# _0455_ 0
C17209 _0983_/a_634_159# _0454_ 0
C17210 acc0.A\[9\] clknet_1_1__leaf__0465_ 0.39385f
C17211 _0286_ hold70/a_49_47# 0
C17212 _0283_ hold70/a_285_47# 0
C17213 _0251_ pp[3] 0
C17214 net183 comp0.B\[14\] 0.20355f
C17215 output58/a_27_47# _0434_ 0.00825f
C17216 _1063_/a_634_159# _1063_/a_466_413# 0.23992f
C17217 _1063_/a_193_47# _1063_/a_1059_315# 0.03405f
C17218 _1063_/a_27_47# _1063_/a_891_413# 0.03089f
C17219 _0645_/a_129_47# acc0.A\[15\] 0
C17220 _0645_/a_285_47# net42 0
C17221 _0174_ net147 0
C17222 acc0.A\[22\] _0374_ 0.00198f
C17223 _0555_/a_51_297# net171 0
C17224 net45 net81 0
C17225 net36 net207 0
C17226 _0975_/a_145_75# control0.state\[2\] 0
C17227 _0975_/a_59_75# _0486_ 0.1711f
C17228 _0658_/a_113_47# _0181_ 0
C17229 clkbuf_1_1__f__0458_/a_110_47# _0826_/a_219_297# 0.0068f
C17230 hold86/a_49_47# _0465_ 0.00353f
C17231 _1019_/a_634_159# _0346_ 0
C17232 _0219_ hold62/a_285_47# 0
C17233 net156 acc0.A\[26\] 0.0307f
C17234 _0179_ _0513_/a_81_21# 0.04103f
C17235 _1037_/a_634_159# _0208_ 0
C17236 net159 _1063_/a_193_47# 0
C17237 _0786_/a_472_297# _0402_ 0
C17238 _1063_/a_1059_315# _0460_ 0.00984f
C17239 _0821_/a_113_47# net63 0
C17240 _0462_ _1006_/a_193_47# 0.00634f
C17241 input32/a_75_212# input22/a_75_212# 0.00122f
C17242 net61 _0629_/a_59_75# 0
C17243 hold86/a_49_47# acc0.A\[2\] 0
C17244 net180 net8 0
C17245 hold58/a_391_47# comp0.B\[2\] 0
C17246 hold52/a_285_47# _1025_/a_27_47# 0
C17247 net158 _1049_/a_466_413# 0
C17248 net89 _0161_ 0
C17249 control0.state\[2\] _0164_ 0
C17250 _0984_/a_1017_47# VPWR 0
C17251 hold74/a_49_47# net43 0.02096f
C17252 _0504_/a_27_47# _0195_ 0
C17253 net44 acc0.A\[30\] 0.16259f
C17254 _0760_/a_47_47# _0219_ 0
C17255 _0819_/a_81_21# clkbuf_0__0465_/a_110_47# 0.01624f
C17256 _0135_ net121 0
C17257 net58 pp[3] 0
C17258 clkbuf_1_0__f__0464_/a_110_47# net154 0
C17259 _1004_/a_891_413# net90 0
C17260 net227 _0707_/a_75_199# 0
C17261 _1011_/a_891_413# acc0.A\[29\] 0.01305f
C17262 _0718_/a_285_47# _0333_ 0
C17263 net197 _1026_/a_891_413# 0.0023f
C17264 _1004_/a_466_413# _1024_/a_193_47# 0
C17265 _1004_/a_27_47# _1024_/a_1059_315# 0
C17266 _1004_/a_193_47# _1024_/a_466_413# 0
C17267 _0732_/a_80_21# _0367_ 0
C17268 _0251_ _0273_ 0.0235f
C17269 _0394_ _0347_ 0.00682f
C17270 _0308_ _0352_ 0
C17271 _1060_/a_634_159# _1060_/a_466_413# 0.23992f
C17272 _1060_/a_193_47# _1060_/a_1059_315# 0.03405f
C17273 _1060_/a_27_47# _1060_/a_891_413# 0.03224f
C17274 _1028_/a_27_47# net94 0
C17275 net114 _1008_/a_27_47# 0.00127f
C17276 _0510_/a_109_47# acc0.A\[10\] 0.00348f
C17277 hold43/a_285_47# _1028_/a_1059_315# 0.0054f
C17278 _0191_ acc0.A\[7\] 0.25144f
C17279 net15 _0252_ 0
C17280 net245 _0797_/a_207_413# 0
C17281 _0195_ _0456_ 0
C17282 _0399_ clknet_0__0461_ 0.00163f
C17283 net187 _0462_ 0.00111f
C17284 _0143_ _1050_/a_634_159# 0
C17285 _0850_/a_68_297# _0265_ 0.00115f
C17286 _1012_/a_193_47# _0097_ 0
C17287 _1012_/a_466_413# _0396_ 0
C17288 hold47/a_391_47# clknet_0__0464_ 0
C17289 net194 clkbuf_0__0464_/a_110_47# 0
C17290 _0805_/a_109_47# clknet_1_1__leaf__0459_ 0
C17291 hold56/a_391_47# _1065_/a_1059_315# 0
C17292 hold56/a_285_47# _1065_/a_891_413# 0
C17293 _1025_/a_27_47# net52 0
C17294 net36 _0551_/a_27_47# 0
C17295 _0218_ net239 0
C17296 _0106_ _0345_ 0
C17297 _0988_/a_891_413# _0988_/a_1017_47# 0.00617f
C17298 _0467_ _0971_/a_299_297# 0.01924f
C17299 _0856_/a_510_47# _0456_ 0.00384f
C17300 _0988_/a_634_159# net74 0
C17301 _0568_/a_27_297# _0704_/a_68_297# 0
C17302 _0553_/a_149_47# _0553_/a_240_47# 0.06872f
C17303 _1067_/a_193_47# clknet_1_1__leaf_clk 0.00976f
C17304 pp[29] _0354_ 0
C17305 output57/a_27_47# _0109_ 0
C17306 net125 _0174_ 0.03139f
C17307 net120 clknet_0__0463_ 0
C17308 _0968_/a_193_297# control0.state\[0\] 0
C17309 _0968_/a_109_297# control0.state\[1\] 0.01243f
C17310 net56 _1011_/a_27_47# 0
C17311 pp[27] _0568_/a_27_297# 0
C17312 _1053_/a_1059_315# _0252_ 0
C17313 _1053_/a_381_47# acc0.A\[7\] 0
C17314 acc0.A\[14\] _0465_ 0.00543f
C17315 _0320_ _0687_/a_145_75# 0
C17316 clknet_1_0__leaf__0460_ _0757_/a_68_297# 0.00224f
C17317 _1041_/a_634_159# _0206_ 0
C17318 _1041_/a_466_413# comp0.B\[8\] 0
C17319 _0982_/a_381_47# _0465_ 0
C17320 _0753_/a_381_47# _0378_ 0
C17321 VPWR _1014_/a_1059_315# 0.3792f
C17322 _1071_/a_193_47# VPWR 0.32489f
C17323 _0327_ _0326_ 0
C17324 _0309_ _0780_/a_285_47# 0
C17325 _0367_ _0250_ 0
C17326 _0542_/a_512_297# _0141_ 0
C17327 acc0.A\[2\] clkbuf_1_0__f__0464_/a_110_47# 0
C17328 _0369_ _0303_ 0
C17329 _0588_/a_113_47# _0220_ 0.00961f
C17330 net58 _0273_ 0
C17331 clknet_1_0__leaf__0457_ _0772_/a_79_21# 0.02117f
C17332 _0984_/a_27_47# hold75/a_49_47# 0
C17333 clkload1/Y clknet_1_0__leaf__0465_ 0.25445f
C17334 _0172_ _1042_/a_634_159# 0.00167f
C17335 _1021_/a_381_47# _0460_ 0.00253f
C17336 _1021_/a_975_413# clknet_1_0__leaf__0457_ 0
C17337 pp[9] pp[10] 0.10265f
C17338 hold46/a_285_47# clknet_0__0464_ 0
C17339 net133 _1047_/a_381_47# 0
C17340 _0386_ acc0.A\[18\] 0
C17341 _0680_/a_80_21# _0250_ 0
C17342 _0716_/a_27_47# net42 0.01009f
C17343 net127 net174 0
C17344 VPWR output40/a_27_47# 0.29616f
C17345 net46 _0383_ 0
C17346 _0257_ _0256_ 0.3615f
C17347 _0992_/a_193_47# net143 0
C17348 clkbuf_0__0464_/a_110_47# _1046_/a_634_159# 0.01021f
C17349 pp[17] pp[30] 0.15535f
C17350 _0309_ _0677_/a_47_47# 0.14426f
C17351 hold73/a_285_47# hold73/a_391_47# 0.41909f
C17352 _0409_ net5 0.09571f
C17353 _0535_/a_68_297# _0473_ 0
C17354 hold79/a_391_47# _0167_ 0
C17355 output54/a_27_47# _1027_/a_27_47# 0
C17356 _1008_/a_27_47# _0365_ 0.03997f
C17357 _0994_/a_27_47# _0347_ 0
C17358 _0144_ _1061_/a_891_413# 0
C17359 _0347_ _1008_/a_592_47# 0.00107f
C17360 net59 VPWR 1.17038f
C17361 _0399_ _0082_ 0
C17362 _0999_/a_193_47# net43 0.00105f
C17363 _1037_/a_1017_47# _0135_ 0.00109f
C17364 net180 net10 0
C17365 _0369_ _0281_ 0
C17366 net175 _1048_/a_634_159# 0.00166f
C17367 _0996_/a_1059_315# hold91/a_391_47# 0.01554f
C17368 _0313_ _0695_/a_80_21# 0
C17369 hold25/a_391_47# _1038_/a_193_47# 0
C17370 hold25/a_285_47# _1038_/a_634_159# 0.00537f
C17371 _0517_/a_81_21# acc0.A\[10\] 0
C17372 _0573_/a_27_47# _0171_ 0
C17373 clknet_1_0__leaf__0464_ _0536_/a_51_297# 0
C17374 _0958_/a_27_47# _1062_/a_27_47# 0
C17375 clkbuf_1_0__f__0465_/a_110_47# _0434_ 0.00122f
C17376 _0097_ clknet_1_1__leaf__0461_ 0.00339f
C17377 _0538_/a_149_47# _1045_/a_27_47# 0
C17378 _0538_/a_51_297# _1045_/a_466_413# 0
C17379 net44 _0779_/a_79_21# 0.08877f
C17380 _0635_/a_27_47# _0267_ 0.05639f
C17381 net149 _1047_/a_27_47# 0.0131f
C17382 hold74/a_285_47# _0181_ 0
C17383 VPWR _1022_/a_27_47# 0.70843f
C17384 output59/a_27_47# _0568_/a_109_297# 0
C17385 hold45/a_285_47# net3 0
C17386 hold9/a_391_47# net113 0
C17387 net44 _0310_ 0
C17388 _0993_/a_193_47# net38 0.00505f
C17389 _0999_/a_27_47# _0999_/a_193_47# 0.96647f
C17390 hold13/a_285_47# _0133_ 0
C17391 _1017_/a_27_47# net221 0
C17392 _0172_ _0562_/a_150_297# 0
C17393 _0121_ net177 0
C17394 hold30/a_391_47# acc0.A\[23\] 0
C17395 VPWR _0679_/a_150_297# 0.00357f
C17396 _1001_/a_634_159# _0772_/a_215_47# 0
C17397 _1001_/a_891_413# _1001_/a_1017_47# 0.00617f
C17398 _0457_ _0173_ 0.00254f
C17399 _0991_/a_1059_315# _0345_ 0.00146f
C17400 hold58/a_49_47# VPWR 0.28222f
C17401 hold47/a_285_47# clknet_1_0__leaf__0464_ 0.01785f
C17402 _0115_ _1060_/a_466_413# 0
C17403 _1035_/a_466_413# net25 0
C17404 _0174_ _0473_ 0.13383f
C17405 net70 clknet_1_1__leaf__0465_ 0
C17406 net60 pp[31] 0.13483f
C17407 _1062_/a_891_413# _1062_/a_975_413# 0.00851f
C17408 _1062_/a_381_47# _1062_/a_561_413# 0.00123f
C17409 net55 _0729_/a_68_297# 0.03047f
C17410 net132 _0527_/a_109_297# 0
C17411 _1011_/a_466_413# _0353_ 0
C17412 net39 _0647_/a_47_47# 0.40026f
C17413 _0472_ comp0.B\[10\] 0.02626f
C17414 net84 _0369_ 0
C17415 _1021_/a_466_413# _1021_/a_381_47# 0.03733f
C17416 _1021_/a_193_47# _1021_/a_975_413# 0
C17417 _1021_/a_1059_315# _1021_/a_891_413# 0.31086f
C17418 _1033_/a_634_159# net23 0
C17419 pp[27] _0109_ 0
C17420 control0.add _0242_ 0.33835f
C17421 net199 _1024_/a_466_413# 0
C17422 hold41/a_391_47# net188 0.13551f
C17423 _0854_/a_510_47# _0453_ 0
C17424 _1017_/a_634_159# _0459_ 0.00641f
C17425 _0147_ _1048_/a_466_413# 0
C17426 _1049_/a_1059_315# net134 0
C17427 _0607_/a_373_47# _0399_ 0
C17428 _0985_/a_27_47# clknet_1_1__leaf__0457_ 0
C17429 clknet_1_0__leaf__0462_ clknet_1_1__leaf__0462_ 0.00361f
C17430 _0732_/a_80_21# _0742_/a_299_297# 0.04251f
C17431 _0124_ VPWR 0.54778f
C17432 _0510_/a_27_297# _0510_/a_373_47# 0.01338f
C17433 _0996_/a_891_413# _0670_/a_215_47# 0
C17434 control0.state\[0\] _0181_ 0
C17435 _0174_ clkbuf_1_1__f__0464_/a_110_47# 0
C17436 acc0.A\[31\] _0708_/a_150_297# 0
C17437 hold15/a_285_47# net60 0
C17438 _0459_ _1060_/a_1017_47# 0
C17439 _0322_ acc0.A\[28\] 0
C17440 _0733_/a_79_199# _0733_/a_544_297# 0.00594f
C17441 _0200_ _0953_/a_32_297# 0.00253f
C17442 _0963_/a_35_297# clk 0.00135f
C17443 hold65/a_49_47# _0274_ 0.00362f
C17444 _0481_ _0167_ 0
C17445 net62 _0988_/a_193_47# 0.01132f
C17446 hold98/a_285_47# net42 0.00451f
C17447 _0327_ acc0.A\[28\] 0
C17448 _1011_/a_27_47# _0345_ 0.03776f
C17449 hold87/a_285_47# net36 0.09277f
C17450 clkbuf_1_0__f__0465_/a_110_47# _0989_/a_1059_315# 0
C17451 net48 _1022_/a_27_47# 0.03212f
C17452 _0294_ _1060_/a_193_47# 0.0016f
C17453 _1031_/a_634_159# _1013_/a_193_47# 0
C17454 _1031_/a_193_47# _1013_/a_634_159# 0
C17455 _1031_/a_466_413# _1013_/a_27_47# 0
C17456 _1031_/a_27_47# _1013_/a_466_413# 0
C17457 control0.state\[1\] _0486_ 0.3849f
C17458 net34 control0.state\[2\] 0.76563f
C17459 clknet_1_1__leaf__0464_ _1043_/a_592_47# 0.00164f
C17460 _0350_ _0219_ 0.6711f
C17461 _0195_ _0568_/a_109_47# 0.00524f
C17462 _0216_ _0568_/a_27_297# 0.20968f
C17463 net132 _1061_/a_193_47# 0
C17464 _1046_/a_193_47# net147 0
C17465 _0372_ acc0.A\[19\] 0.0035f
C17466 _0111_ _0219_ 0.00815f
C17467 _0953_/a_32_297# comp0.B\[8\] 0.16441f
C17468 net149 clknet_1_0__leaf__0461_ 0.24871f
C17469 _1034_/a_466_413# clknet_0__0463_ 0
C17470 _1034_/a_381_47# clkbuf_1_1__f__0463_/a_110_47# 0.00126f
C17471 _0799_/a_209_297# net41 0
C17472 hold26/a_391_47# net152 0
C17473 hold26/a_285_47# net32 0
C17474 _0503_/a_109_297# _0217_ 0
C17475 hold38/a_391_47# _1034_/a_466_413# 0
C17476 acc0.A\[8\] _0826_/a_27_53# 0
C17477 _0260_ _0636_/a_59_75# 0.03806f
C17478 hold17/a_391_47# _1071_/a_27_47# 0.00285f
C17479 hold17/a_285_47# _1071_/a_193_47# 0.00241f
C17480 hold17/a_49_47# _1071_/a_634_159# 0.00168f
C17481 hold78/a_285_47# net225 0.00999f
C17482 _0984_/a_193_47# _0399_ 0
C17483 comp0.B\[5\] _0562_/a_68_297# 0
C17484 _0750_/a_109_47# _0460_ 0
C17485 hold31/a_49_47# _0438_ 0
C17486 _0561_/a_51_297# _0132_ 0.22637f
C17487 _0717_/a_80_21# pp[17] 0
C17488 VPWR _1067_/a_634_159# 0.20206f
C17489 hold29/a_49_47# _1022_/a_1059_315# 0
C17490 _1050_/a_27_47# _0186_ 0.02936f
C17491 hold100/a_391_47# _0263_ 0.0503f
C17492 _0251_ _0086_ 0.00232f
C17493 _0466_ _0468_ 0.63101f
C17494 net17 _1062_/a_193_47# 0
C17495 _0313_ _0743_/a_512_297# 0
C17496 _0515_/a_299_297# _0189_ 0.00955f
C17497 _1033_/a_27_47# clknet_1_0__leaf__0461_ 0
C17498 _0228_ _1005_/a_193_47# 0
C17499 _0982_/a_466_413# _0263_ 0
C17500 pp[17] _0339_ 0.00741f
C17501 net62 net72 0.32981f
C17502 hold88/a_285_47# net58 0
C17503 _0640_/a_297_297# _0271_ 0
C17504 _1020_/a_1059_315# net106 0
C17505 _0450_ net72 0
C17506 _0691_/a_68_297# _0181_ 0
C17507 _0248_ clkbuf_1_0__f__0460_/a_110_47# 0
C17508 _0473_ _0208_ 0
C17509 _0618_/a_215_47# _0618_/a_510_47# 0.00529f
C17510 _0475_ _0173_ 0.06328f
C17511 hold14/a_49_47# hold14/a_391_47# 0.00188f
C17512 _1036_/a_1017_47# clknet_1_1__leaf__0463_ 0
C17513 VPWR _0335_ 0.46315f
C17514 _0389_ _0771_/a_215_297# 0.10343f
C17515 _0243_ _0771_/a_27_413# 0.09158f
C17516 acc0.A\[7\] input11/a_75_212# 0
C17517 _0226_ _0594_/a_113_47# 0.00951f
C17518 _0348_ _1030_/a_466_413# 0.00106f
C17519 _0510_/a_373_47# _0181_ 0.00259f
C17520 _0644_/a_129_47# _0304_ 0
C17521 _0461_ _1019_/a_975_413# 0
C17522 _0346_ _0431_ 0.24338f
C17523 _0425_ _0345_ 0.05376f
C17524 _0314_ _0345_ 0.04965f
C17525 _0401_ _0814_/a_109_47# 0.00151f
C17526 _1001_/a_891_413# _0218_ 0.00276f
C17527 _0343_ pp[1] 0
C17528 _0179_ hold83/a_49_47# 0
C17529 _0956_/a_32_297# _0214_ 0.02854f
C17530 _0133_ _0132_ 0.07206f
C17531 _0372_ _0249_ 0
C17532 _1041_/a_891_413# comp0.B\[9\] 0.00304f
C17533 _1047_/a_466_413# _0145_ 0.03715f
C17534 net45 _0790_/a_35_297# 0
C17535 hold12/a_391_47# _0237_ 0
C17536 hold12/a_49_47# _0382_ 0
C17537 hold1/a_285_47# _0085_ 0
C17538 hold1/a_391_47# net73 0
C17539 _0346_ _0659_/a_68_297# 0.0138f
C17540 net65 _0431_ 0
C17541 net81 VPWR 0.3443f
C17542 hold61/a_285_47# hold62/a_49_47# 0
C17543 net157 _1048_/a_27_47# 0
C17544 net185 _0213_ 0
C17545 _0973_/a_109_297# net107 0
C17546 net53 pp[25] 0.00955f
C17547 _0399_ clkbuf_0__0458_/a_110_47# 0.00556f
C17548 net125 _1046_/a_193_47# 0
C17549 _0725_/a_209_297# _0334_ 0
C17550 _0343_ _0337_ 0.02179f
C17551 net58 _0086_ 0.17551f
C17552 _0710_/a_109_47# _0345_ 0
C17553 hold41/a_391_47# _0155_ 0
C17554 _0183_ _1018_/a_561_413# 0
C17555 net28 _0175_ 0.00388f
C17556 _1004_/a_1059_315# _0756_/a_47_47# 0
C17557 net236 _0468_ 0.05648f
C17558 _0536_/a_149_47# _0472_ 0
C17559 _0465_ _0823_/a_109_297# 0
C17560 net243 _1004_/a_592_47# 0
C17561 _0253_ net74 0.009f
C17562 _0525_/a_81_21# _0193_ 0
C17563 output44/a_27_47# hold15/a_49_47# 0.008f
C17564 _0123_ _1007_/a_27_47# 0
C17565 _0328_ _0740_/a_113_47# 0
C17566 _0440_ _0442_ 0.10005f
C17567 _0233_ _0183_ 0
C17568 _0518_/a_27_297# _0186_ 0.1367f
C17569 _0805_/a_27_47# _0418_ 0
C17570 hold69/a_391_47# net92 0
C17571 _0217_ _0575_/a_373_47# 0.00365f
C17572 hold42/a_391_47# net37 0.01054f
C17573 _0733_/a_79_199# _0317_ 0
C17574 _1057_/a_891_413# net37 0.0038f
C17575 _0234_ net213 0.01623f
C17576 _0514_/a_109_47# net142 0
C17577 _1034_/a_27_47# _1034_/a_634_159# 0.13601f
C17578 _0536_/a_51_297# _0536_/a_245_297# 0.01218f
C17579 _0101_ _0487_ 0.00166f
C17580 _0796_/a_79_21# _0796_/a_510_47# 0.00844f
C17581 _0796_/a_297_297# _0796_/a_215_47# 0
C17582 net44 _0239_ 0.17727f
C17583 net162 _1030_/a_193_47# 0
C17584 net168 _1053_/a_193_47# 0
C17585 _0559_/a_51_297# hold58/a_285_47# 0.0017f
C17586 _0216_ _0109_ 0.00822f
C17587 hold10/a_285_47# comp0.B\[15\] 0.00799f
C17588 _0993_/a_193_47# _0282_ 0
C17589 net104 _0580_/a_27_297# 0
C17590 clknet_0__0464_ clkbuf_1_0__f__0464_/a_110_47# 0.31134f
C17591 net64 _0826_/a_27_53# 0
C17592 _0253_ output61/a_27_47# 0
C17593 _0626_/a_68_297# _0268_ 0
C17594 net133 net149 0
C17595 net185 _0212_ 0.08166f
C17596 net147 comp0.B\[9\] 0
C17597 _1057_/a_561_413# net67 0
C17598 hold25/a_49_47# _0550_/a_240_47# 0
C17599 _0982_/a_466_413# clknet_1_0__leaf__0461_ 0.00116f
C17600 clkbuf_0_clk/a_110_47# _0161_ 0.00275f
C17601 _1038_/a_1059_315# net28 0
C17602 _1013_/a_193_47# _0345_ 0.00234f
C17603 _0983_/a_1017_47# _0081_ 0
C17604 net69 _0454_ 0.06806f
C17605 hold69/a_285_47# _0240_ 0
C17606 VPWR A[15] 0.33854f
C17607 clkbuf_0__0464_/a_110_47# _1045_/a_27_47# 0.00212f
C17608 _0517_/a_299_297# _0181_ 0
C17609 _1063_/a_634_159# _0161_ 0.04087f
C17610 net235 _0988_/a_27_47# 0.00217f
C17611 _0746_/a_81_21# _0350_ 0.04856f
C17612 _0195_ _0095_ 0
C17613 _0854_/a_79_21# acc0.A\[18\] 0
C17614 control0.count\[3\] _1072_/a_27_47# 0.43185f
C17615 output56/a_27_47# acc0.A\[29\] 0
C17616 net105 _0346_ 0.02177f
C17617 net78 _0992_/a_27_47# 0.22901f
C17618 _0305_ acc0.A\[13\] 0
C17619 acc0.A\[8\] _0087_ 0.14513f
C17620 acc0.A\[1\] hold2/a_391_47# 0.06769f
C17621 _0326_ _0346_ 0
C17622 _0399_ net67 0.05041f
C17623 hold96/a_285_47# net176 0
C17624 _0226_ _0101_ 0
C17625 VPWR _1024_/a_466_413# 0.25501f
C17626 _0959_/a_80_21# _0470_ 0.11005f
C17627 _0432_ _0345_ 0.06941f
C17628 _0585_/a_27_297# net149 0.07258f
C17629 net203 _0563_/a_245_297# 0.00225f
C17630 _0550_/a_51_297# net7 0
C17631 _0982_/a_1059_315# net47 0
C17632 _0172_ net31 0.15135f
C17633 clknet_1_0__leaf__0464_ _1050_/a_381_47# 0
C17634 _1049_/a_891_413# acc0.A\[15\] 0
C17635 _0586_/a_27_47# _0218_ 0.1767f
C17636 _0677_/a_285_47# net43 0
C17637 VPWR _1048_/a_891_413# 0.19525f
C17638 net18 _0542_/a_149_47# 0.00363f
C17639 _0343_ _0406_ 0.26373f
C17640 acc0.A\[4\] hold7/a_49_47# 0.29428f
C17641 _1028_/a_592_47# clknet_1_1__leaf__0462_ 0.00168f
C17642 _0731_/a_81_21# _0312_ 0.01226f
C17643 net158 _0147_ 0
C17644 _1055_/a_1059_315# net66 0
C17645 _1055_/a_466_413# acc0.A\[8\] 0
C17646 _0795_/a_81_21# _0407_ 0
C17647 comp0.B\[13\] _0473_ 0.3223f
C17648 _0601_/a_150_297# _0223_ 0
C17649 _0642_/a_382_47# _0253_ 0
C17650 comp0.B\[1\] net24 0.00175f
C17651 pp[27] _0725_/a_80_21# 0
C17652 hold47/a_285_47# hold47/a_391_47# 0.41909f
C17653 _0809_/a_384_47# net228 0
C17654 _0197_ clknet_1_1__leaf__0457_ 0
C17655 hold13/a_285_47# _0174_ 0
C17656 _0473_ _1046_/a_193_47# 0.01618f
C17657 _0355_ _0339_ 0
C17658 net227 _0338_ 0.00282f
C17659 net178 _0990_/a_891_413# 0
C17660 _1004_/a_193_47# _0122_ 0
C17661 VPWR _1010_/a_592_47# 0
C17662 _1000_/a_466_413# _1000_/a_381_47# 0.03733f
C17663 _1000_/a_193_47# _1000_/a_975_413# 0
C17664 _1000_/a_1059_315# _1000_/a_891_413# 0.31086f
C17665 _0993_/a_27_47# _0281_ 0
C17666 _1060_/a_466_413# net146 0.00156f
C17667 _1060_/a_634_159# _0158_ 0.00401f
C17668 VPWR _0797_/a_207_413# 0.16762f
C17669 _1051_/a_1059_315# net154 0
C17670 _1051_/a_193_47# net11 0.00219f
C17671 _0256_ clknet_1_1__leaf__0458_ 0
C17672 control0.count\[1\] _0979_/a_27_297# 0.0013f
C17673 net230 net168 0.11668f
C17674 _0459_ _0508_/a_81_21# 0
C17675 _1072_/a_466_413# VPWR 0.24813f
C17676 VPWR _0841_/a_215_47# 0.00128f
C17677 _1053_/a_1017_47# net11 0
C17678 net125 comp0.B\[9\] 0
C17679 _0143_ net136 0
C17680 _0300_ hold91/a_49_47# 0
C17681 comp0.B\[13\] clkbuf_1_1__f__0464_/a_110_47# 0
C17682 _0555_/a_51_297# _0553_/a_51_297# 0
C17683 _0953_/a_220_297# comp0.B\[9\] 0.0073f
C17684 hold56/a_49_47# control0.reset 0.02015f
C17685 _0329_ _1011_/a_193_47# 0
C17686 acc0.A\[12\] _0289_ 0
C17687 _0128_ _0704_/a_68_297# 0
C17688 _0399_ _0986_/a_975_413# 0
C17689 net240 _1063_/a_27_47# 0
C17690 net207 hold60/a_391_47# 0.15273f
C17691 pp[27] _0128_ 0.00328f
C17692 VPWR _1009_/a_1017_47# 0
C17693 clknet_1_1__leaf__0459_ _0650_/a_150_297# 0
C17694 hold14/a_391_47# _0208_ 0
C17695 _0698_/a_199_47# _0330_ 0.00151f
C17696 _0451_ net47 0
C17697 net27 _0173_ 0.0151f
C17698 _0457_ _1033_/a_1059_315# 0.01715f
C17699 _0280_ _0420_ 0.0093f
C17700 _0537_/a_150_297# comp0.B\[12\] 0
C17701 _0231_ _0379_ 0
C17702 _0979_/a_109_297# clkbuf_1_0__f_clk/a_110_47# 0
C17703 _0361_ _0181_ 0
C17704 _1050_/a_27_47# _1050_/a_634_159# 0.14145f
C17705 hold59/a_49_47# _0854_/a_79_21# 0
C17706 VPWR _0741_/a_109_297# 0.00597f
C17707 hold37/a_285_47# clknet_0__0464_ 0.02356f
C17708 _0959_/a_472_297# _0160_ 0.00467f
C17709 _1019_/a_27_47# clknet_1_0__leaf__0457_ 0
C17710 comp0.B\[13\] hold49/a_49_47# 0
C17711 net23 _0487_ 0
C17712 _1032_/a_27_47# control0.reset 0
C17713 hold85/a_49_47# net17 0.04854f
C17714 hold74/a_285_47# clknet_1_1__leaf__0461_ 0.10501f
C17715 clkload1/a_268_47# _0432_ 0
C17716 _0221_ _1011_/a_193_47# 0.02039f
C17717 _0311_ clknet_0__0460_ 0
C17718 clknet_1_1__leaf__0460_ _0780_/a_35_297# 0
C17719 _0271_ _0261_ 0
C17720 _1018_/a_466_413# _0181_ 0
C17721 clknet_1_1__leaf__0463_ _1065_/a_466_413# 0
C17722 _0179_ _1049_/a_891_413# 0.05112f
C17723 net113 _0352_ 0
C17724 _0819_/a_299_297# _0401_ 0.06521f
C17725 _0427_ _0815_/a_113_297# 0
C17726 _0430_ _0437_ 0
C17727 net36 _0199_ 0.01559f
C17728 _0621_/a_285_47# _0437_ 0
C17729 _0999_/a_634_159# _1012_/a_193_47# 0
C17730 _0999_/a_466_413# _1012_/a_27_47# 0
C17731 _0999_/a_27_47# _1012_/a_466_413# 0
C17732 _0625_/a_59_75# _0625_/a_145_75# 0.00658f
C17733 _0222_ _0754_/a_240_47# 0.02994f
C17734 _0346_ _0269_ 0
C17735 clkbuf_0__0464_/a_110_47# net132 0.04547f
C17736 _0997_/a_466_413# pp[14] 0
C17737 _0997_/a_891_413# net41 0.0337f
C17738 clkbuf_1_1__f__0463_/a_110_47# net201 0
C17739 _1071_/a_891_413# clknet_0_clk 0.00239f
C17740 _1008_/a_592_47# _0106_ 0.00164f
C17741 _0313_ _0329_ 0.00866f
C17742 _0670_/a_79_21# _0277_ 0.00116f
C17743 _0559_/a_51_297# _0134_ 0
C17744 VPWR comp0.B\[12\] 1.0848f
C17745 hold13/a_285_47# _0208_ 0.0022f
C17746 _0397_ _0307_ 0.14502f
C17747 net224 _1009_/a_27_47# 0.0085f
C17748 _0472_ _0177_ 0
C17749 clknet_1_0__leaf__0461_ _0393_ 0
C17750 acc0.A\[5\] _0437_ 0
C17751 net175 net134 0.00208f
C17752 _0313_ clknet_1_0__leaf__0460_ 0
C17753 _0577_/a_109_47# VPWR 0.00392f
C17754 hold25/a_49_47# net172 0
C17755 hold25/a_285_47# net124 0
C17756 net46 _0756_/a_129_47# 0
C17757 control0.state\[2\] _1066_/a_466_413# 0
C17758 acc0.A\[14\] _1060_/a_634_159# 0.00166f
C17759 _0343_ _0307_ 0
C17760 _0477_ _1062_/a_27_47# 0.03721f
C17761 _1020_/a_193_47# net187 0
C17762 comp0.B\[4\] _0176_ 0
C17763 net25 _0561_/a_51_297# 0.12659f
C17764 hold46/a_49_47# hold46/a_285_47# 0.22264f
C17765 _1000_/a_193_47# _1018_/a_891_413# 0
C17766 control0.state\[2\] _1068_/a_466_413# 0
C17767 _0486_ _1068_/a_634_159# 0.01692f
C17768 _0143_ _1045_/a_193_47# 0.00198f
C17769 net183 _1045_/a_891_413# 0
C17770 _0998_/a_1059_315# net42 0.00227f
C17771 net35 _0487_ 0.52752f
C17772 _0200_ _0535_/a_68_297# 0.10555f
C17773 hold58/a_49_47# _1036_/a_27_47# 0
C17774 net22 net18 0
C17775 _0606_/a_215_297# _0460_ 0.00355f
C17776 hold70/a_285_47# _0345_ 0.00628f
C17777 _1055_/a_634_159# _0290_ 0
C17778 _0343_ _1000_/a_193_47# 0.02321f
C17779 _0308_ _0392_ 0
C17780 _0610_/a_145_75# _0242_ 0
C17781 net202 clknet_1_0__leaf__0460_ 0
C17782 _0999_/a_466_413# _0999_/a_592_47# 0.00553f
C17783 _0999_/a_634_159# _0999_/a_1017_47# 0
C17784 net17 _1063_/a_975_413# 0
C17785 _0339_ _0567_/a_109_297# 0.00585f
C17786 _0992_/a_381_47# _0090_ 0.11467f
C17787 hold48/a_49_47# _0537_/a_68_297# 0
C17788 _0473_ comp0.B\[9\] 0.28037f
C17789 _1001_/a_27_47# _1019_/a_1059_315# 0.00319f
C17790 _1001_/a_466_413# _1019_/a_193_47# 0
C17791 _1001_/a_193_47# _1019_/a_466_413# 0
C17792 _1017_/a_381_47# _0115_ 0.12032f
C17793 _0754_/a_245_297# _0103_ 0
C17794 _0731_/a_299_297# _0219_ 0
C17795 _0583_/a_109_297# clknet_1_1__leaf__0461_ 0
C17796 VPWR _0993_/a_466_413# 0.26095f
C17797 _1001_/a_891_413# _0099_ 0
C17798 _0629_/a_59_75# _0269_ 0
C17799 _0565_/a_149_47# comp0.B\[0\] 0.00253f
C17800 clknet_1_0__leaf__0462_ _1007_/a_466_413# 0.01645f
C17801 _0404_ hold91/a_49_47# 0
C17802 hold24/a_285_47# net29 0.00147f
C17803 _0697_/a_80_21# _0360_ 0
C17804 _0356_ clknet_1_1__leaf__0462_ 0
C17805 _0639_/a_109_297# _0186_ 0
C17806 _0133_ net25 0.19467f
C17807 _0534_/a_384_47# _0465_ 0
C17808 _0983_/a_193_47# _0217_ 0
C17809 hold88/a_49_47# net47 0.0027f
C17810 hold47/a_391_47# comp0.B\[14\] 0
C17811 _1020_/a_381_47# net202 0.00194f
C17812 _0186_ _0987_/a_27_47# 0.00953f
C17813 net67 _0295_ 0
C17814 _0216_ _0725_/a_80_21# 0
C17815 _0370_ _0318_ 0
C17816 _1043_/a_634_159# _0542_/a_51_297# 0.00163f
C17817 _0695_/a_80_21# clkbuf_0__0460_/a_110_47# 0.01002f
C17818 hold100/a_285_47# _0267_ 0
C17819 _0305_ net45 0.04634f
C17820 _1021_/a_381_47# _0119_ 0.13132f
C17821 net119 net23 0
C17822 _0181_ acc0.A\[13\] 0
C17823 net199 _0122_ 0
C17824 _0558_/a_68_297# net25 0.01144f
C17825 _0558_/a_150_297# B[2] 0
C17826 net82 acc0.A\[14\] 0
C17827 clknet_0__0461_ _0306_ 0
C17828 net103 _0459_ 0.01706f
C17829 _0218_ net149 0
C17830 _0174_ _0200_ 0.12866f
C17831 clknet_1_1__leaf__0459_ acc0.A\[15\] 0.03489f
C17832 _0510_/a_373_47# _0187_ 0
C17833 control0.count\[2\] _0979_/a_109_297# 0.00236f
C17834 _0133_ _0477_ 0.00226f
C17835 clknet_1_0__leaf__0465_ hold7/a_285_47# 0.02183f
C17836 _1017_/a_466_413# _0218_ 0
C17837 _0257_ clknet_0__0465_ 0.00631f
C17838 _1051_/a_193_47# clknet_1_1__leaf__0458_ 0
C17839 VPWR _0790_/a_35_297# 0.31745f
C17840 _1043_/a_891_413# net20 0
C17841 hold77/a_49_47# acc0.A\[27\] 0
C17842 _1002_/a_27_47# clknet_1_0__leaf__0460_ 0.0259f
C17843 acc0.A\[20\] _0352_ 0.53326f
C17844 _1006_/a_634_159# _0219_ 0
C17845 _0174_ comp0.B\[8\] 0.02708f
C17846 _0482_ clknet_1_0__leaf_clk 0
C17847 acc0.A\[12\] _0655_/a_109_93# 0.00667f
C17848 hold87/a_49_47# _0346_ 0
C17849 _0800_/a_149_47# net81 0
C17850 _0751_/a_183_297# _0219_ 0
C17851 _0216_ _0128_ 0.03839f
C17852 hold41/a_49_47# acc0.A\[11\] 0.04619f
C17853 _1050_/a_27_47# net62 0
C17854 _0467_ _1068_/a_1059_315# 0.00154f
C17855 _0518_/a_27_297# _0518_/a_109_47# 0.00393f
C17856 _0120_ _0224_ 0.00228f
C17857 acc0.A\[22\] _0225_ 0.07882f
C17858 _0461_ _0773_/a_285_47# 0
C17859 _0985_/a_27_47# _0985_/a_891_413# 0.03224f
C17860 _0985_/a_193_47# _0985_/a_1059_315# 0.03405f
C17861 _0985_/a_634_159# _0985_/a_466_413# 0.23992f
C17862 comp0.B\[2\] clkbuf_1_1__f__0463_/a_110_47# 0.02216f
C17863 _0217_ _0526_/a_27_47# 0
C17864 hold46/a_285_47# comp0.B\[14\] 0.06228f
C17865 net193 _0535_/a_68_297# 0.00242f
C17866 _0973_/a_27_297# net17 0.00623f
C17867 _0780_/a_285_297# _0397_ 0.07186f
C17868 _1018_/a_27_47# _1018_/a_466_413# 0.26005f
C17869 _1018_/a_193_47# _1018_/a_634_159# 0.11072f
C17870 clknet_1_0__leaf__0465_ net21 0.00426f
C17871 control0.count\[2\] _1071_/a_975_413# 0
C17872 _0985_/a_193_47# _1049_/a_193_47# 0.00131f
C17873 net46 net110 0.00763f
C17874 net50 _1022_/a_634_159# 0
C17875 net194 _1050_/a_193_47# 0
C17876 _0208_ _0132_ 0.0165f
C17877 _0818_/a_109_47# clknet_0__0465_ 0
C17878 hold29/a_285_47# net151 0
C17879 _0590_/a_113_47# net177 0
C17880 acc0.A\[12\] _0418_ 0.00461f
C17881 _0785_/a_81_21# _0817_/a_81_21# 0
C17882 _0171_ acc0.A\[15\] 0.23874f
C17883 clknet_1_1__leaf_clk _0951_/a_109_93# 0.01228f
C17884 _0080_ _0263_ 0
C17885 _0651_/a_113_47# acc0.A\[10\] 0
C17886 _0296_ _0670_/a_79_21# 0
C17887 _1019_/a_1059_315# _0459_ 0.00134f
C17888 hold99/a_49_47# VPWR 0.31375f
C17889 _0753_/a_79_21# _0343_ 0.1703f
C17890 net68 _1047_/a_193_47# 0
C17891 _0152_ _0619_/a_68_297# 0
C17892 hold44/a_285_47# _0195_ 0
C17893 _0330_ hold50/a_391_47# 0
C17894 VPWR _0756_/a_285_47# 0.00344f
C17895 _0172_ _0548_/a_240_47# 0.04791f
C17896 _0276_ _0669_/a_29_53# 0.30566f
C17897 _1054_/a_27_47# input15/a_75_212# 0
C17898 _0644_/a_47_47# _0301_ 0.00157f
C17899 _0734_/a_285_47# _0359_ 0
C17900 VPWR _1027_/a_561_413# 0.00306f
C17901 _0555_/a_51_297# _0135_ 0.10689f
C17902 hold79/a_49_47# hold79/a_391_47# 0.00188f
C17903 _0586_/a_27_47# _0099_ 0.0526f
C17904 net44 _0309_ 0.04067f
C17905 VPWR _0749_/a_299_297# 0.28279f
C17906 _0693_/a_68_297# _0366_ 0.00322f
C17907 _0350_ net94 0.01611f
C17908 _0101_ _0760_/a_47_47# 0
C17909 _0997_/a_466_413# _0408_ 0
C17910 VPWR _0678_/a_150_297# 0.00228f
C17911 VPWR _1052_/a_27_47# 0.47958f
C17912 net193 _0174_ 0.14801f
C17913 _0179_ clknet_1_1__leaf__0459_ 0
C17914 _0338_ net208 0.00981f
C17915 _1023_/a_27_47# _1022_/a_27_47# 0.0011f
C17916 _0328_ _0694_/a_113_47# 0
C17917 _0317_ clkbuf_1_1__f__0462_/a_110_47# 0.00966f
C17918 _1056_/a_466_413# acc0.A\[10\] 0.00731f
C17919 clk _0484_ 0.06549f
C17920 net45 _0675_/a_150_297# 0
C17921 _0240_ acc0.A\[18\] 0
C17922 hold3/a_49_47# _0460_ 0
C17923 net233 _0265_ 0
C17924 _0743_/a_149_47# _0360_ 0.02871f
C17925 _0487_ _1063_/a_466_413# 0.00443f
C17926 net152 _1040_/a_27_47# 0
C17927 _0655_/a_109_93# _0650_/a_68_297# 0
C17928 _1019_/a_891_413# clknet_1_0__leaf__0461_ 0
C17929 comp0.B\[10\] _1046_/a_891_413# 0
C17930 net248 _0399_ 0
C17931 _1004_/a_381_47# _0379_ 0
C17932 clknet_0__0457_ acc0.A\[18\] 0
C17933 net55 _0357_ 0.04697f
C17934 _0415_ _0648_/a_27_297# 0
C17935 _0346_ _0991_/a_381_47# 0.00674f
C17936 _0600_/a_253_47# acc0.A\[23\] 0
C17937 net9 _0142_ 0
C17938 _0191_ _0186_ 0.00311f
C17939 _0994_/a_1059_315# net80 0
C17940 _0176_ _0541_/a_150_297# 0
C17941 hold78/a_391_47# _0341_ 0.05507f
C17942 hold78/a_285_47# _0340_ 0
C17943 _0544_/a_240_47# _0204_ 0
C17944 net61 _0253_ 0.00112f
C17945 _0544_/a_512_297# net198 0.00173f
C17946 _0345_ _0360_ 0.05523f
C17947 net10 hold51/a_391_47# 0.01981f
C17948 _0121_ hold4/a_49_47# 0
C17949 _0371_ _0460_ 0.02877f
C17950 _0637_/a_139_47# _0263_ 0.01023f
C17951 _1034_/a_891_413# _1034_/a_975_413# 0.00851f
C17952 _1034_/a_381_47# _1034_/a_561_413# 0.00123f
C17953 _0504_/a_27_47# _0183_ 0.33356f
C17954 net206 clknet_1_0__leaf__0461_ 0.27713f
C17955 _0343_ _0507_/a_109_297# 0.00102f
C17956 output64/a_27_47# pp[8] 0
C17957 _1021_/a_1017_47# acc0.A\[21\] 0
C17958 B[2] input27/a_75_212# 0.07726f
C17959 input25/a_75_212# B[4] 0.0033f
C17960 hold6/a_49_47# hold6/a_285_47# 0.22264f
C17961 _0480_ _0976_/a_505_21# 0.0013f
C17962 net67 _0811_/a_299_297# 0.0027f
C17963 acc0.A\[23\] _1006_/a_27_47# 0
C17964 net48 _0749_/a_299_297# 0
C17965 hold59/a_285_47# _0195_ 0
C17966 _0080_ clknet_1_0__leaf__0461_ 0.00188f
C17967 _0816_/a_68_297# _0816_/a_150_297# 0.00477f
C17968 _0640_/a_392_297# clknet_0__0465_ 0
C17969 _0627_/a_297_297# VPWR 0
C17970 _0183_ _0456_ 0.42423f
C17971 _0499_/a_59_75# _0178_ 0.11057f
C17972 clknet_0__0464_ _1045_/a_381_47# 0.00108f
C17973 hold10/a_285_47# _0176_ 0
C17974 hold54/a_285_47# control0.reset 0
C17975 _0481_ hold79/a_49_47# 0.05773f
C17976 _0218_ _0094_ 0.00202f
C17977 _0225_ _0379_ 0.00737f
C17978 _0179_ _0292_ 0.12231f
C17979 _0483_ _0169_ 0
C17980 net58 _0991_/a_27_47# 0
C17981 VPWR _1026_/a_1017_47# 0
C17982 net59 net56 0
C17983 _0848_/a_109_297# _0451_ 0
C17984 _0225_ _0372_ 0.0024f
C17985 hold78/a_391_47# _1013_/a_891_413# 0
C17986 _0343_ _0333_ 0.04395f
C17987 VPWR _0817_/a_266_47# 0.00645f
C17988 pp[16] net41 0.0574f
C17989 acc0.A\[20\] net207 0
C17990 _0549_/a_150_297# _0176_ 0
C17991 _1001_/a_193_47# _0352_ 0
C17992 _0793_/a_149_47# net42 0.00413f
C17993 _0793_/a_51_297# _0406_ 0
C17994 pp[30] _1031_/a_27_47# 0.00246f
C17995 VPWR _0122_ 0.22871f
C17996 net45 _0181_ 0.035f
C17997 clknet_0__0459_ net42 0
C17998 _0626_/a_68_297# _0443_ 0.00142f
C17999 pp[15] _1013_/a_1059_315# 0.00108f
C18000 clknet_0_clk _0972_/a_93_21# 0
C18001 net149 _0112_ 0.01962f
C18002 _0172_ net7 0.43488f
C18003 _0559_/a_240_47# _0211_ 0
C18004 _1071_/a_1059_315# _0488_ 0
C18005 _1071_/a_466_413# _0466_ 0.00854f
C18006 _1018_/a_1059_315# _0242_ 0
C18007 clknet_1_0__leaf__0464_ acc0.A\[4\] 0.11188f
C18008 hold76/a_49_47# _0244_ 0.00243f
C18009 _0993_/a_634_159# _0286_ 0
C18010 net81 _0995_/a_634_159# 0
C18011 hold77/a_391_47# _1009_/a_27_47# 0
C18012 hold77/a_285_47# _1009_/a_193_47# 0
C18013 hold8/a_285_47# _0352_ 0
C18014 clknet_1_0__leaf__0460_ _1005_/a_592_47# 0
C18015 _1017_/a_634_159# _1017_/a_592_47# 0
C18016 net179 acc0.A\[8\] 0
C18017 _0708_/a_68_297# _0708_/a_150_297# 0.00477f
C18018 hold13/a_391_47# _0555_/a_51_297# 0
C18019 _1058_/a_27_47# net3 0
C18020 _0753_/a_381_47# _0375_ 0.00264f
C18021 _0753_/a_79_21# _0376_ 0.04733f
C18022 _0233_ _0752_/a_27_413# 0
C18023 _0723_/a_27_413# hold80/a_391_47# 0.00266f
C18024 clknet_1_0__leaf__0459_ _0790_/a_35_297# 0
C18025 _1052_/a_891_413# net9 0.03228f
C18026 _0343_ _0732_/a_80_21# 0
C18027 _0251_ _0621_/a_35_297# 0
C18028 _0786_/a_80_21# _0422_ 0.00308f
C18029 net24 _0496_/a_27_47# 0.0536f
C18030 _0644_/a_285_47# _0346_ 0
C18031 comp0.B\[7\] net180 0.23584f
C18032 hold24/a_285_47# _0137_ 0
C18033 _0984_/a_381_47# _0219_ 0
C18034 _0504_/a_27_47# acc0.A\[15\] 0.07277f
C18035 net190 hold50/a_391_47# 0
C18036 _0831_/a_35_297# clkbuf_1_1__f__0458_/a_110_47# 0.0081f
C18037 _1006_/a_381_47# net52 0
C18038 _1000_/a_381_47# _0098_ 0.11464f
C18039 _0507_/a_27_297# net5 0.19659f
C18040 _1000_/a_466_413# net45 0.01988f
C18041 _0232_ clknet_1_0__leaf__0460_ 0.01377f
C18042 net58 _0350_ 0.07992f
C18043 _0464_ _1048_/a_193_47# 0
C18044 comp0.B\[1\] clknet_1_0__leaf__0457_ 0
C18045 _1056_/a_1059_315# hold34/a_391_47# 0
C18046 _1056_/a_891_413# hold34/a_285_47# 0
C18047 _0430_ _0252_ 0.02268f
C18048 net146 _0158_ 0.01766f
C18049 _0259_ _0431_ 0
C18050 _0543_/a_68_297# _0543_/a_150_297# 0.00477f
C18051 comp0.B\[13\] _0200_ 0.00674f
C18052 pp[18] acc0.A\[31\] 0.2223f
C18053 _0804_/a_79_21# _0415_ 0.0963f
C18054 hold82/a_391_47# acc0.A\[13\] 0
C18055 _0456_ acc0.A\[15\] 0
C18056 _0216_ _0601_/a_150_297# 0
C18057 _0521_/a_81_21# _0521_/a_384_47# 0.00138f
C18058 _0200_ _1046_/a_193_47# 0
C18059 _1033_/a_634_159# _1033_/a_466_413# 0.23992f
C18060 _1033_/a_193_47# _1033_/a_1059_315# 0.03405f
C18061 _1033_/a_27_47# _1033_/a_891_413# 0.03224f
C18062 _0655_/a_109_93# net42 0
C18063 hold36/a_285_47# net20 0
C18064 _0259_ _0659_/a_68_297# 0.04891f
C18065 VPWR _0951_/a_209_311# 0.19687f
C18066 _0343_ clkbuf_1_0__f__0460_/a_110_47# 0.02191f
C18067 acc0.A\[5\] _0252_ 0
C18068 net64 _0465_ 0.00256f
C18069 net55 _0734_/a_285_47# 0
C18070 clknet_0__0458_ _0835_/a_215_47# 0
C18071 _1012_/a_634_159# _1012_/a_466_413# 0.23992f
C18072 _1012_/a_193_47# _1012_/a_1059_315# 0.03405f
C18073 _1012_/a_27_47# _1012_/a_891_413# 0.03224f
C18074 _0853_/a_68_297# net222 0
C18075 _0196_ _0527_/a_27_297# 0.12497f
C18076 _0287_ _0424_ 0
C18077 _0216_ _0331_ 0
C18078 _0346_ _0082_ 0.0033f
C18079 _0758_/a_79_21# _0105_ 0
C18080 _0352_ _1007_/a_891_413# 0
C18081 _1056_/a_1059_315# _0510_/a_27_297# 0.00101f
C18082 _0512_/a_27_297# _0186_ 0.09525f
C18083 _0399_ _0302_ 0
C18084 _0107_ _1009_/a_193_47# 0.21404f
C18085 _0195_ _1031_/a_381_47# 0.00492f
C18086 _0216_ _1031_/a_1059_315# 0
C18087 _0363_ _1009_/a_1059_315# 0
C18088 net211 _0369_ 0.00556f
C18089 _0343_ _0250_ 0.05128f
C18090 _0476_ _0957_/a_304_297# 0
C18091 net37 _0419_ 0
C18092 clknet_0__0457_ net211 0.32126f
C18093 net227 _0332_ 0
C18094 net58 _0621_/a_35_297# 0.01139f
C18095 _0343_ hold98/a_391_47# 0.03807f
C18096 _1072_/a_561_413# clknet_0_clk 0.00112f
C18097 _1050_/a_891_413# _1050_/a_975_413# 0.00851f
C18098 _1050_/a_27_47# net136 0.2266f
C18099 _1050_/a_381_47# _1050_/a_561_413# 0.00123f
C18100 _0272_ VPWR 0.37086f
C18101 _0990_/a_1059_315# _0181_ 0.0058f
C18102 net35 _0760_/a_47_47# 0
C18103 _1041_/a_1059_315# _0546_/a_51_297# 0.00134f
C18104 _1041_/a_27_47# _0546_/a_240_47# 0
C18105 _0218_ _0393_ 0.11251f
C18106 _1024_/a_891_413# net50 0.00132f
C18107 clknet_1_0__leaf__0464_ _1051_/a_466_413# 0
C18108 hold74/a_391_47# net44 0
C18109 _0195_ _0589_/a_113_47# 0
C18110 VPWR _0837_/a_368_297# 0.00925f
C18111 _0764_/a_81_21# _0462_ 0.02419f
C18112 net61 output61/a_27_47# 0.2423f
C18113 _0515_/a_81_21# acc0.A\[9\] 0
C18114 _0241_ _1019_/a_193_47# 0
C18115 hold24/a_285_47# comp0.B\[6\] 0.0012f
C18116 clkbuf_1_0__f__0465_/a_110_47# _0186_ 0
C18117 _0180_ _0527_/a_373_47# 0.00267f
C18118 control0.state\[1\] _0965_/a_47_47# 0.00108f
C18119 net233 _0267_ 0
C18120 _0305_ VPWR 1.65042f
C18121 _0349_ VPWR 0.37211f
C18122 _0544_/a_51_297# _1043_/a_27_47# 0
C18123 _0461_ _0386_ 0.00606f
C18124 _0998_/a_592_47# net43 0
C18125 hold16/a_391_47# _0704_/a_68_297# 0.01241f
C18126 _1054_/a_381_47# _1052_/a_1059_315# 0
C18127 _0802_/a_145_75# _0403_ 0
C18128 _0504_/a_27_47# _0179_ 0
C18129 _0176_ _1040_/a_381_47# 0.01948f
C18130 _1014_/a_466_413# hold2/a_285_47# 0
C18131 _1014_/a_1059_315# hold2/a_49_47# 0
C18132 _1014_/a_634_159# hold2/a_391_47# 0
C18133 _0179_ _1054_/a_466_413# 0.00837f
C18134 net46 _0618_/a_79_21# 0
C18135 net21 _1044_/a_466_413# 0.0105f
C18136 _0143_ _1044_/a_27_47# 0
C18137 _0566_/a_27_47# clknet_1_1__leaf__0457_ 0
C18138 clknet_0__0465_ clknet_1_1__leaf__0458_ 0.06305f
C18139 acc0.A\[14\] net146 0.09752f
C18140 net21 net137 0
C18141 _0337_ _0568_/a_27_297# 0
C18142 net45 _1018_/a_27_47# 0
C18143 net25 _0208_ 0.13144f
C18144 comp0.B\[13\] net193 0.17849f
C18145 _0995_/a_466_413# _0797_/a_27_413# 0.00154f
C18146 net59 _0345_ 0.01712f
C18147 _1056_/a_1059_315# _0181_ 0.01152f
C18148 control0.state\[2\] _0166_ 0.02046f
C18149 _1031_/a_27_47# _0339_ 0.0364f
C18150 _0750_/a_109_47# _0373_ 0
C18151 net205 _1036_/a_1059_315# 0
C18152 _0973_/a_27_297# _0165_ 0.11038f
C18153 _0973_/a_373_47# net240 0.00122f
C18154 _0555_/a_149_47# _0208_ 0.03196f
C18155 _0820_/a_79_21# _0369_ 0.15099f
C18156 _0270_ _0638_/a_109_297# 0.01253f
C18157 net193 _1046_/a_193_47# 0
C18158 comp0.B\[13\] _1046_/a_466_413# 0
C18159 _0360_ net52 0
C18160 hold98/a_285_47# net60 0
C18161 _0459_ _0774_/a_68_297# 0.00461f
C18162 comp0.B\[2\] _0163_ 0
C18163 _0574_/a_27_297# _1007_/a_381_47# 0
C18164 _1054_/a_634_159# net75 0
C18165 _0182_ _1061_/a_1059_315# 0
C18166 _0444_ _0840_/a_68_297# 0
C18167 comp0.B\[15\] _1047_/a_27_47# 0
C18168 _1012_/a_634_159# net98 0
C18169 _1012_/a_1059_315# clknet_1_1__leaf__0461_ 0
C18170 _1046_/a_27_47# _1046_/a_1059_315# 0.04672f
C18171 _1046_/a_193_47# _1046_/a_466_413# 0.07855f
C18172 pp[30] _0712_/a_79_21# 0
C18173 _0978_/a_109_297# _0466_ 0.05817f
C18174 _0978_/a_109_47# _0488_ 0
C18175 _0999_/a_1017_47# net85 0
C18176 _1019_/a_1059_315# _0772_/a_79_21# 0
C18177 clknet_1_1__leaf__0463_ B[1] 0.02439f
C18178 _0130_ _0173_ 0
C18179 hold55/a_391_47# _0208_ 0.00984f
C18180 acc0.A\[20\] net106 0
C18181 _0256_ _0218_ 0.12905f
C18182 net223 _0391_ 0.30104f
C18183 _1056_/a_193_47# _0517_/a_299_297# 0.00112f
C18184 _1056_/a_27_47# _0517_/a_384_47# 0
C18185 _1032_/a_634_159# clknet_1_0__leaf__0457_ 0.00205f
C18186 _1016_/a_561_413# net221 0.00197f
C18187 _1016_/a_634_159# _0115_ 0.0014f
C18188 _0968_/a_193_297# VPWR 0.00131f
C18189 _0221_ _0707_/a_75_199# 0.10691f
C18190 _0752_/a_384_47# _0376_ 0.00124f
C18191 clknet_1_0__leaf__0462_ _0105_ 0.19176f
C18192 net45 _0677_/a_377_297# 0
C18193 _0329_ _0321_ 0.08127f
C18194 _0181_ clkbuf_1_1__f_clk/a_110_47# 0.00589f
C18195 hold18/a_391_47# _0219_ 0
C18196 _1050_/a_27_47# _1045_/a_193_47# 0
C18197 _1050_/a_193_47# _1045_/a_27_47# 0
C18198 _0775_/a_215_47# _0393_ 0.00622f
C18199 _0996_/a_466_413# acc0.A\[15\] 0.00538f
C18200 _0996_/a_1059_315# net42 0.01385f
C18201 _0984_/a_193_47# _0346_ 0.01486f
C18202 clknet_0__0463_ _0175_ 0.19474f
C18203 clknet_1_0__leaf__0463_ _1038_/a_193_47# 0.03845f
C18204 _0200_ comp0.B\[9\] 0.08264f
C18205 _0172_ comp0.B\[11\] 0
C18206 hold64/a_49_47# acc0.A\[18\] 0
C18207 _0211_ _1036_/a_466_413# 0
C18208 net129 _0542_/a_51_297# 0.00523f
C18209 _1043_/a_466_413# net19 0
C18210 clkbuf_0__0460_/a_110_47# clknet_1_0__leaf__0460_ 0
C18211 _0822_/a_109_297# clknet_1_1__leaf__0458_ 0
C18212 hold38/a_49_47# _0215_ 0
C18213 hold38/a_391_47# _0175_ 0.01984f
C18214 acc0.A\[12\] _1057_/a_466_413# 0
C18215 VPWR _0701_/a_209_297# 0.19563f
C18216 _0399_ net6 0.02206f
C18217 _0662_/a_81_21# _0423_ 0.05193f
C18218 hold27/a_285_47# _0472_ 0
C18219 _0723_/a_27_413# _0336_ 0
C18220 _0723_/a_207_413# _0220_ 0
C18221 VPWR hold73/a_49_47# 0.27439f
C18222 _1033_/a_975_413# net17 0
C18223 _0479_ _0486_ 0
C18224 _0693_/a_68_297# acc0.A\[24\] 0.18992f
C18225 _0457_ _1032_/a_27_47# 0.0167f
C18226 _0857_/a_27_47# _1032_/a_891_413# 0.00936f
C18227 net85 clknet_1_1__leaf__0461_ 0.15919f
C18228 pp[8] net3 0
C18229 net58 _0839_/a_109_297# 0
C18230 net44 _0999_/a_466_413# 0
C18231 comp0.B\[8\] comp0.B\[9\] 0.31016f
C18232 net59 hold16/a_49_47# 0
C18233 _0229_ _0750_/a_181_47# 0
C18234 _0226_ _0750_/a_27_47# 0.19748f
C18235 _0648_/a_27_297# _0347_ 0
C18236 _0262_ _0350_ 0
C18237 _0181_ _0584_/a_109_297# 0.01788f
C18238 hold34/a_391_47# VPWR 0.1592f
C18239 _1000_/a_634_159# net46 0
C18240 _0294_ _1016_/a_27_47# 0.005f
C18241 hold37/a_285_47# comp0.B\[14\] 0.00146f
C18242 _1052_/a_466_413# _0522_/a_109_297# 0
C18243 _0195_ _0219_ 0.52483f
C18244 hold20/a_285_47# _0484_ 0
C18245 net162 _0567_/a_27_297# 0.12101f
C18246 net92 _0219_ 0
C18247 clknet_0__0459_ _0645_/a_377_297# 0
C18248 _0598_/a_297_47# acc0.A\[21\] 0.0016f
C18249 _0598_/a_382_297# _0227_ 0.01509f
C18250 _0518_/a_109_47# _0191_ 0
C18251 VPWR _0675_/a_150_297# 0.00135f
C18252 net61 _0446_ 0.19286f
C18253 _0217_ output50/a_27_47# 0
C18254 _1039_/a_634_159# net8 0.03522f
C18255 _1038_/a_1059_315# clknet_0__0463_ 0
C18256 _0985_/a_634_159# _0083_ 0.0392f
C18257 _0195_ _0728_/a_59_75# 0
C18258 _0214_ _0562_/a_150_297# 0
C18259 clkbuf_1_0__f__0463_/a_110_47# _1040_/a_1059_315# 0.022f
C18260 pp[28] hold16/a_285_47# 0
C18261 hold10/a_391_47# _0501_/a_27_47# 0
C18262 VPWR _0510_/a_27_297# 0.18833f
C18263 _0326_ _1007_/a_381_47# 0
C18264 _0165_ net17 0.30317f
C18265 _1018_/a_193_47# net104 0.00747f
C18266 _1018_/a_1059_315# _1018_/a_1017_47# 0
C18267 hold67/a_49_47# clknet_1_1__leaf__0465_ 0.01965f
C18268 _0463_ _0957_/a_32_297# 0
C18269 comp0.B\[15\] clknet_1_0__leaf__0461_ 0.03852f
C18270 net232 _0485_ 0
C18271 _0789_/a_208_47# _0409_ 0
C18272 _0299_ _0795_/a_299_297# 0
C18273 hold47/a_391_47# acc0.A\[4\] 0.00117f
C18274 _0734_/a_47_47# _0326_ 0
C18275 _0982_/a_634_159# _0982_/a_592_47# 0
C18276 hold88/a_285_47# _0833_/a_79_21# 0
C18277 _1011_/a_891_413# clknet_1_1__leaf__0462_ 0
C18278 _1049_/a_466_413# _1049_/a_561_413# 0.00772f
C18279 _1049_/a_634_159# _1049_/a_975_413# 0
C18280 net145 _0346_ 0
C18281 _0983_/a_1017_47# acc0.A\[15\] 0
C18282 hold65/a_49_47# _0433_ 0.00202f
C18283 _0210_ net29 0
C18284 net148 acc0.A\[6\] 0
C18285 net12 _0522_/a_373_47# 0
C18286 _0194_ _0522_/a_109_297# 0
C18287 _0115_ _0116_ 0
C18288 hold56/a_49_47# _0475_ 0
C18289 _0172_ _0202_ 0.02699f
C18290 _0747_/a_79_21# _0747_/a_215_47# 0.04584f
C18291 net48 hold73/a_49_47# 0.32234f
C18292 _0552_/a_150_297# _0209_ 0
C18293 VPWR _0618_/a_297_297# 0.01069f
C18294 net40 input6/a_75_212# 0.00797f
C18295 _1052_/a_27_47# _0523_/a_81_21# 0.00185f
C18296 _1053_/a_27_47# _1053_/a_466_413# 0.27314f
C18297 _1053_/a_193_47# _1053_/a_634_159# 0.12729f
C18298 _0575_/a_27_297# _0575_/a_109_47# 0.00393f
C18299 _0137_ _0138_ 0
C18300 _0714_/a_51_297# _0218_ 0.04958f
C18301 _1019_/a_891_413# _0218_ 0
C18302 net193 comp0.B\[9\] 0
C18303 _0195_ _1008_/a_634_159# 0
C18304 hold39/a_391_47# _1065_/a_27_47# 0
C18305 _0348_ net208 0
C18306 _1066_/a_193_47# _1066_/a_592_47# 0
C18307 _1066_/a_466_413# _1066_/a_561_413# 0.00772f
C18308 _1066_/a_634_159# _1066_/a_975_413# 0
C18309 _0627_/a_215_53# acc0.A\[6\] 0.00103f
C18310 _0328_ _0350_ 0
C18311 _0831_/a_117_297# acc0.A\[8\] 0
C18312 _0327_ _1010_/a_27_47# 0
C18313 _0849_/a_215_47# _0263_ 0
C18314 control0.reset _0562_/a_68_297# 0
C18315 net45 _0999_/a_1017_47# 0
C18316 _0678_/a_68_297# _0777_/a_47_47# 0.00204f
C18317 pp[0] input28/a_75_212# 0
C18318 _0201_ _1042_/a_193_47# 0
C18319 net31 _1040_/a_193_47# 0
C18320 _1023_/a_381_47# _1022_/a_891_413# 0
C18321 _0833_/a_79_21# _0086_ 0.05058f
C18322 _0833_/a_510_47# net235 0.00455f
C18323 _0680_/a_217_297# _0462_ 0.00601f
C18324 _1068_/a_466_413# _1068_/a_561_413# 0.00772f
C18325 _1068_/a_634_159# _1068_/a_975_413# 0
C18326 _0401_ _0809_/a_384_47# 0
C18327 A[0] net1 0.00739f
C18328 _1030_/a_634_159# _1030_/a_466_413# 0.23992f
C18329 _1030_/a_193_47# _1030_/a_1059_315# 0.03405f
C18330 _1030_/a_27_47# _1030_/a_891_413# 0.03089f
C18331 _1041_/a_193_47# _0176_ 0
C18332 _0350_ _0599_/a_113_47# 0
C18333 _0254_ acc0.A\[8\] 0.05041f
C18334 _0439_ _0181_ 0
C18335 _0712_/a_79_21# _0339_ 0.04697f
C18336 acc0.A\[22\] hold68/a_391_47# 0
C18337 net105 _0782_/a_27_47# 0
C18338 _0399_ acc0.A\[0\] 0
C18339 _0946_/a_30_53# net226 0
C18340 _0487_ _0161_ 0.1656f
C18341 _0218_ net206 0.03935f
C18342 VPWR _0181_ 6.88618f
C18343 net76 net47 0.01809f
C18344 net81 _0345_ 0
C18345 _1034_/a_27_47# control0.sh 0
C18346 hold41/a_49_47# A[12] 0
C18347 _0305_ clknet_1_0__leaf__0459_ 0.05138f
C18348 _0330_ _0726_/a_245_297# 0
C18349 hold9/a_49_47# hold9/a_391_47# 0.00188f
C18350 _0429_ _0519_/a_81_21# 0.00165f
C18351 _0092_ _0279_ 0.14209f
C18352 clkbuf_1_1__f__0461_/a_110_47# acc0.A\[17\] 0.06659f
C18353 net148 _0523_/a_384_47# 0.01035f
C18354 _0524_/a_27_297# _0150_ 0
C18355 _0346_ net67 0.01836f
C18356 _1035_/a_891_413# clknet_1_1__leaf__0463_ 0.00685f
C18357 _1035_/a_466_413# net122 0
C18358 _0753_/a_297_297# net46 0.00283f
C18359 _0992_/a_193_47# net37 0
C18360 _0804_/a_79_21# _0347_ 0.11911f
C18361 _0786_/a_80_21# _0423_ 0
C18362 _0216_ _0611_/a_68_297# 0.02202f
C18363 _0770_/a_79_21# acc0.A\[19\] 0
C18364 hold53/a_391_47# net200 0.14498f
C18365 net198 _0140_ 0.11568f
C18366 _0110_ _0308_ 0
C18367 clkbuf_1_0__f__0459_/a_110_47# _0507_/a_109_297# 0.0012f
C18368 _1015_/a_466_413# _0181_ 0.00536f
C18369 _0987_/a_27_47# _0987_/a_634_159# 0.14145f
C18370 _0081_ _0219_ 0
C18371 _0152_ net65 0.00118f
C18372 hold64/a_49_47# net211 0.00115f
C18373 _0182_ _0631_/a_109_297# 0
C18374 net45 clknet_1_1__leaf__0461_ 0.23811f
C18375 _0946_/a_30_53# _0946_/a_112_297# 0.00501f
C18376 _1051_/a_975_413# _0186_ 0.00107f
C18377 _1034_/a_561_413# comp0.B\[2\] 0.00227f
C18378 net194 _1045_/a_27_47# 0
C18379 _0313_ _0696_/a_109_297# 0.00482f
C18380 _0125_ _1008_/a_466_413# 0
C18381 acc0.A\[27\] _1008_/a_381_47# 0
C18382 _0992_/a_466_413# net67 0
C18383 _0340_ clknet_1_1__leaf__0462_ 0.00103f
C18384 _1000_/a_466_413# VPWR 0.24856f
C18385 _0307_ clkbuf_0__0461_/a_110_47# 0.00312f
C18386 control0.count\[3\] _0467_ 0
C18387 net164 _0488_ 0.14046f
C18388 _0480_ _0466_ 0.04413f
C18389 _1072_/a_891_413# _0466_ 0
C18390 _0151_ _1053_/a_27_47# 0.14345f
C18391 net43 _0407_ 0.00246f
C18392 _0369_ _0826_/a_27_53# 0
C18393 hold89/a_391_47# clk 0.01358f
C18394 _0299_ net6 0.18583f
C18395 net133 comp0.B\[15\] 0.02673f
C18396 clknet_1_1__leaf__0462_ _0737_/a_35_297# 0.00126f
C18397 _0232_ hold94/a_285_47# 0
C18398 _0346_ _1006_/a_975_413# 0
C18399 _1029_/a_27_47# _1029_/a_634_159# 0.14145f
C18400 hold2/a_391_47# net247 0
C18401 net14 hold21/a_285_47# 0
C18402 net48 _0181_ 0
C18403 _0255_ _0444_ 0
C18404 _0352_ _0772_/a_297_297# 0
C18405 acc0.A\[1\] _0869_/a_27_47# 0
C18406 _1032_/a_561_413# clknet_1_0__leaf__0461_ 0
C18407 hold57/a_391_47# net36 0
C18408 _0703_/a_109_297# _0334_ 0
C18409 clknet_0_clk net231 0.35137f
C18410 _0805_/a_27_47# _0417_ 0.08788f
C18411 _0716_/a_27_47# _0303_ 0
C18412 _0343_ _0998_/a_891_413# 0.00322f
C18413 _0581_/a_109_47# _0393_ 0
C18414 _0722_/a_297_297# clknet_1_1__leaf__0462_ 0
C18415 net90 _0219_ 0
C18416 comp0.B\[13\] _1045_/a_193_47# 0.00164f
C18417 _0399_ _0580_/a_109_297# 0.04086f
C18418 _1050_/a_27_47# net73 0
C18419 net136 _0987_/a_27_47# 0.00144f
C18420 hold33/a_285_47# hold26/a_49_47# 0.03151f
C18421 hold66/a_285_47# _0754_/a_51_297# 0
C18422 _0645_/a_47_47# _0996_/a_891_413# 0
C18423 _1015_/a_27_47# _0565_/a_51_297# 0
C18424 clknet_1_0__leaf__0465_ _0536_/a_512_297# 0
C18425 _1017_/a_592_47# net103 0.00301f
C18426 net119 _0161_ 0.0024f
C18427 clknet_1_0__leaf__0463_ _0550_/a_512_297# 0
C18428 _1017_/a_381_47# _1016_/a_193_47# 0.00117f
C18429 _0520_/a_109_47# _0180_ 0.00302f
C18430 _0587_/a_27_47# clknet_1_1__leaf__0461_ 0.00917f
C18431 net160 _1036_/a_1059_315# 0
C18432 net64 _0254_ 0.24391f
C18433 hold30/a_285_47# net51 0
C18434 net236 _0480_ 0.00214f
C18435 _0094_ net228 0.00174f
C18436 _0227_ net49 0.25928f
C18437 net166 _1060_/a_193_47# 0
C18438 _1037_/a_634_159# clknet_1_1__leaf__0463_ 0
C18439 _0756_/a_47_47# _1023_/a_466_413# 0
C18440 _0756_/a_285_47# _1023_/a_27_47# 0
C18441 _0208_ _0352_ 0.02667f
C18442 net5 _0185_ 0.00277f
C18443 _0098_ net45 0
C18444 _1033_/a_27_47# _0956_/a_32_297# 0.00106f
C18445 _0998_/a_634_159# clkbuf_1_1__f__0461_/a_110_47# 0.00983f
C18446 _0555_/a_51_297# _0555_/a_240_47# 0.03076f
C18447 _1028_/a_27_47# _1028_/a_193_47# 0.96054f
C18448 _0565_/a_240_47# _0171_ 0
C18449 _0428_ acc0.A\[9\] 0.05344f
C18450 _0606_/a_215_297# _0373_ 0.00197f
C18451 A[12] _0513_/a_299_297# 0
C18452 hold41/a_285_47# _1057_/a_27_47# 0
C18453 _0416_ _0092_ 0
C18454 _0660_/a_113_47# acc0.A\[9\] 0
C18455 _1067_/a_381_47# _1065_/a_27_47# 0
C18456 _1067_/a_193_47# _1065_/a_891_413# 0
C18457 _0399_ _0790_/a_285_297# 0
C18458 net204 _0136_ 0
C18459 net58 _0986_/a_634_159# 0
C18460 _0192_ _0151_ 0.09197f
C18461 _1033_/a_634_159# _0131_ 0.00108f
C18462 _0985_/a_193_47# VPWR 0.31889f
C18463 net63 _0987_/a_466_413# 0
C18464 _0102_ net51 0
C18465 clkbuf_0__0462_/a_110_47# _0319_ 0.00537f
C18466 _0965_/a_377_297# _0478_ 0.00581f
C18467 VPWR _1018_/a_27_47# 0.43512f
C18468 _1039_/a_592_47# _0176_ 0.00285f
C18469 _0130_ _1033_/a_1059_315# 0.00479f
C18470 _0722_/a_79_21# _0720_/a_68_297# 0
C18471 _0985_/a_1059_315# _0636_/a_59_75# 0
C18472 _0846_/a_149_47# _0219_ 0
C18473 net226 _0487_ 0
C18474 _0244_ _0582_/a_109_297# 0
C18475 _1056_/a_1059_315# _0187_ 0
C18476 hold55/a_49_47# hold55/a_391_47# 0.00188f
C18477 _0243_ _1000_/a_1059_315# 0
C18478 net46 _0242_ 0.20684f
C18479 _0743_/a_51_297# _0366_ 0
C18480 hold22/a_49_47# _0179_ 0.03899f
C18481 _0372_ _0462_ 0.12368f
C18482 hold4/a_285_47# _1005_/a_1059_315# 0.0013f
C18483 _1009_/a_381_47# _0219_ 0.00253f
C18484 clkbuf_1_0__f__0465_/a_110_47# net62 0
C18485 _0459_ hold72/a_391_47# 0.01133f
C18486 _0664_/a_79_21# _0401_ 0
C18487 _0343_ _1030_/a_1017_47# 0
C18488 hold54/a_285_47# _0457_ 0.00321f
C18489 _1055_/a_975_413# acc0.A\[9\] 0
C18490 net194 net132 0.03878f
C18491 hold26/a_49_47# net20 0.0013f
C18492 _1041_/a_891_413# net32 0.00183f
C18493 _1041_/a_634_159# _0139_ 0.00226f
C18494 VPWR _0677_/a_377_297# 0.00367f
C18495 _0519_/a_81_21# clknet_1_1__leaf__0458_ 0.01417f
C18496 hold37/a_49_47# hold37/a_285_47# 0.22264f
C18497 _0337_ _0725_/a_80_21# 0
C18498 _0967_/a_215_297# _0946_/a_30_53# 0
C18499 _0946_/a_112_297# _0487_ 0
C18500 _0350_ _0988_/a_975_413# 0
C18501 clkbuf_1_1__f__0459_/a_110_47# acc0.A\[13\] 0.00155f
C18502 _0517_/a_299_297# clknet_1_1__leaf__0465_ 0
C18503 _0508_/a_299_297# net228 0.05895f
C18504 comp0.B\[4\] net28 0
C18505 _0229_ _0606_/a_109_53# 0
C18506 VPWR _0544_/a_240_47# 0.00216f
C18507 _0993_/a_634_159# net79 0
C18508 _0108_ _0350_ 0.14497f
C18509 _0983_/a_466_413# _1018_/a_466_413# 0
C18510 hold87/a_391_47# _0459_ 0
C18511 _0828_/a_113_297# _0828_/a_199_47# 0
C18512 VPWR _1034_/a_891_413# 0.17741f
C18513 _0715_/a_27_47# acc0.A\[9\] 0
C18514 clknet_1_0__leaf__0460_ _1067_/a_466_413# 0
C18515 _0462_ hold40/a_49_47# 0
C18516 net18 _1043_/a_193_47# 0.01948f
C18517 net198 _1043_/a_634_159# 0.02128f
C18518 _0369_ _0087_ 0.01074f
C18519 net163 acc0.A\[30\] 0.0908f
C18520 _0960_/a_109_47# control0.count\[1\] 0
C18521 _0343_ _0983_/a_193_47# 0.01849f
C18522 _0531_/a_27_297# _0531_/a_373_47# 0.01338f
C18523 clknet_1_0__leaf__0459_ _0181_ 0.07675f
C18524 clknet_1_0__leaf__0462_ _0359_ 0.00412f
C18525 _0578_/a_27_297# clknet_1_0__leaf__0457_ 0.02213f
C18526 clkbuf_1_0__f__0458_/a_110_47# _0219_ 0
C18527 _0553_/a_240_47# _0463_ 0
C18528 _0179_ net169 0.10045f
C18529 _1053_/a_466_413# A[5] 0.00158f
C18530 _1002_/a_634_159# acc0.A\[20\] 0
C18531 _0998_/a_634_159# _0998_/a_1059_315# 0
C18532 _0998_/a_27_47# _0998_/a_381_47# 0.05761f
C18533 _0998_/a_193_47# _0998_/a_891_413# 0.19421f
C18534 pp[17] _0708_/a_150_297# 0
C18535 _0195_ hold61/a_49_47# 0
C18536 _0337_ _0128_ 0.00898f
C18537 net126 comp0.B\[8\] 0.19257f
C18538 hold41/a_49_47# _0154_ 0
C18539 _1003_/a_634_159# _0369_ 0
C18540 _0343_ _0287_ 0
C18541 _0796_/a_510_47# _0400_ 0
C18542 _0498_/a_149_47# _1061_/a_27_47# 0
C18543 _1024_/a_27_47# net177 0
C18544 _0122_ _1023_/a_27_47# 0
C18545 net110 _1023_/a_193_47# 0
C18546 hold56/a_49_47# _1033_/a_193_47# 0.01265f
C18547 hold56/a_285_47# _1033_/a_27_47# 0.00137f
C18548 net8 net147 0.00226f
C18549 _0396_ _0395_ 0.09259f
C18550 VPWR _0507_/a_373_47# 0
C18551 _0174_ _1044_/a_27_47# 0
C18552 _1001_/a_975_413# _0350_ 0
C18553 net118 _0584_/a_373_47# 0
C18554 _1019_/a_27_47# _1019_/a_1059_315# 0.04875f
C18555 _1019_/a_193_47# _1019_/a_466_413# 0.08301f
C18556 net44 _1012_/a_891_413# 0.00495f
C18557 _1046_/a_891_413# _1046_/a_1017_47# 0.00617f
C18558 _0798_/a_113_297# _0798_/a_199_47# 0
C18559 _0143_ _0196_ 0
C18560 _1019_/a_891_413# _0099_ 0
C18561 net31 _0207_ 0
C18562 acc0.A\[4\] clkbuf_1_0__f__0464_/a_110_47# 0
C18563 pp[26] net190 0
C18564 _1056_/a_891_413# _0153_ 0
C18565 _0809_/a_299_297# hold70/a_285_47# 0
C18566 clknet_1_0__leaf__0463_ net29 0.07178f
C18567 _0341_ net116 0
C18568 clknet_1_1__leaf__0458_ _0986_/a_27_47# 0
C18569 net133 _0533_/a_109_47# 0
C18570 VPWR _1012_/a_193_47# 0.3255f
C18571 VPWR hold82/a_391_47# 0.18531f
C18572 _0221_ _0338_ 0.03988f
C18573 net133 hold71/a_285_47# 0
C18574 _0964_/a_109_297# _0484_ 0.00124f
C18575 _0218_ _0405_ 0
C18576 _1051_/a_1059_315# _1050_/a_381_47# 0
C18577 _1051_/a_381_47# _1050_/a_1059_315# 0
C18578 _0565_/a_51_297# _0215_ 0.12561f
C18579 _0684_/a_59_75# _0316_ 0.11023f
C18580 _0548_/a_51_297# _1040_/a_891_413# 0
C18581 clknet_1_0__leaf__0462_ net200 0.06638f
C18582 _0985_/a_592_47# net175 0
C18583 _0642_/a_27_413# clknet_0__0465_ 0
C18584 _0453_ _0181_ 0.02628f
C18585 net196 net19 0.05006f
C18586 _0211_ net161 0.00331f
C18587 net9 _1049_/a_466_413# 0.00262f
C18588 net175 _1049_/a_381_47# 0
C18589 acc0.A\[12\] net189 0.13243f
C18590 hold54/a_285_47# _0475_ 0
C18591 control0.sh _0565_/a_149_47# 0
C18592 _0210_ comp0.B\[6\] 0.04987f
C18593 _0974_/a_79_199# _0468_ 0.11527f
C18594 acc0.A\[31\] _1031_/a_193_47# 0
C18595 hold15/a_391_47# _1031_/a_1059_315# 0.00145f
C18596 hold15/a_285_47# _1031_/a_891_413# 0
C18597 _1041_/a_891_413# net10 0
C18598 net207 _0208_ 0
C18599 _0340_ hold92/a_49_47# 0
C18600 hold3/a_49_47# _0373_ 0.01021f
C18601 _0585_/a_27_297# hold71/a_285_47# 0
C18602 hold76/a_391_47# _0247_ 0
C18603 control0.state\[1\] clknet_0_clk 0.09496f
C18604 _0280_ _0347_ 0.0273f
C18605 _1021_/a_193_47# _0578_/a_27_297# 0.0018f
C18606 net86 net46 0
C18607 hold88/a_285_47# hold88/a_391_47# 0.41909f
C18608 _0568_/a_27_297# _0333_ 0
C18609 _0722_/a_79_21# net116 0
C18610 _0758_/a_215_47# _0758_/a_510_47# 0.00529f
C18611 _1024_/a_193_47# pp[24] 0
C18612 _1024_/a_466_413# net52 0.00493f
C18613 VPWR _0999_/a_1017_47# 0
C18614 hold32/a_49_47# A[12] 0
C18615 clkload3/a_268_47# net84 0
C18616 _1052_/a_592_47# acc0.A\[6\] 0.00143f
C18617 _1052_/a_1059_315# _0193_ 0.0045f
C18618 _1052_/a_381_47# net13 0
C18619 hold35/a_391_47# _0181_ 0
C18620 _0246_ _0347_ 0
C18621 _0990_/a_634_159# _0990_/a_466_413# 0.23992f
C18622 _0990_/a_193_47# _0990_/a_1059_315# 0.03112f
C18623 _0990_/a_27_47# _0990_/a_891_413# 0.03089f
C18624 _0463_ _0213_ 0.00244f
C18625 _0211_ net26 0.02742f
C18626 _0732_/a_209_47# VPWR 0
C18627 clknet_0__0461_ net221 0
C18628 _0790_/a_35_297# _0345_ 0.00603f
C18629 _0313_ hold90/a_285_47# 0
C18630 net168 _0519_/a_384_47# 0.01008f
C18631 _0218_ _0773_/a_35_297# 0
C18632 _0733_/a_448_47# clkbuf_0__0462_/a_110_47# 0.00159f
C18633 _0179_ clkbuf_1_1__f__0465_/a_110_47# 0.02168f
C18634 net125 net8 0.03549f
C18635 _0984_/a_381_47# net58 0
C18636 VPWR _0187_ 0.23687f
C18637 _0641_/a_113_47# _0435_ 0
C18638 _0464_ acc0.A\[15\] 0.09385f
C18639 _0747_/a_79_21# _0352_ 0.14377f
C18640 _0174_ _0546_/a_245_297# 0.00263f
C18641 net150 _0228_ 0.66518f
C18642 _0985_/a_561_413# acc0.A\[3\] 0
C18643 _0967_/a_109_93# _0967_/a_215_297# 0.15204f
C18644 _0967_/a_215_297# _0487_ 0
C18645 _0967_/a_297_297# _0485_ 0
C18646 acc0.A\[25\] _1007_/a_634_159# 0
C18647 _0485_ _0162_ 0.10961f
C18648 _0343_ _0793_/a_240_47# 0.00174f
C18649 hold97/a_49_47# _0322_ 0.00212f
C18650 pp[18] _0708_/a_68_297# 0.00534f
C18651 output45/a_27_47# net60 0.00763f
C18652 comp0.B\[10\] _0546_/a_149_47# 0.00191f
C18653 net248 _0346_ 0.07829f
C18654 _1021_/a_27_47# net202 0
C18655 hold53/a_285_47# _1025_/a_27_47# 0.00403f
C18656 hold88/a_391_47# _0086_ 0
C18657 _1049_/a_1059_315# acc0.A\[3\] 0.08391f
C18658 clknet_0__0465_ _0218_ 0.00171f
C18659 _1034_/a_27_47# _0955_/a_32_297# 0.00139f
C18660 hold97/a_49_47# _0327_ 0
C18661 _1021_/a_27_47# clknet_1_1__leaf__0463_ 0
C18662 _1011_/a_1059_315# hold80/a_285_47# 0.0054f
C18663 VPWR clknet_1_1__leaf__0461_ 3.32712f
C18664 hold9/a_391_47# _0739_/a_79_21# 0
C18665 _0409_ _0669_/a_29_53# 0
C18666 clknet_1_0__leaf__0459_ _1018_/a_27_47# 0
C18667 _0229_ hold3/a_285_47# 0
C18668 net248 net65 0
C18669 net248 _0989_/a_466_413# 0
C18670 _0551_/a_27_47# _0208_ 0.15369f
C18671 _1070_/a_193_47# _1070_/a_592_47# 0.00135f
C18672 _1070_/a_466_413# _1070_/a_561_413# 0.00772f
C18673 _1070_/a_634_159# _1070_/a_975_413# 0
C18674 net10 net147 0
C18675 _1052_/a_466_413# _0150_ 0.03276f
C18676 clknet_0__0459_ acc0.A\[17\] 0
C18677 _1053_/a_193_47# net139 0.00518f
C18678 _1053_/a_1059_315# _1053_/a_1017_47# 0
C18679 pp[17] _1030_/a_466_413# 0
C18680 net44 _1030_/a_891_413# 0.05074f
C18681 _1015_/a_891_413# net118 0
C18682 net189 _0650_/a_68_297# 0
C18683 clknet_1_0__leaf__0465_ _1050_/a_975_413# 0
C18684 net225 _0218_ 0.09527f
C18685 _0960_/a_181_47# control0.count\[2\] 0.00228f
C18686 net45 _0998_/a_561_413# 0
C18687 acc0.A\[22\] _1023_/a_891_413# 0
C18688 _0183_ _1023_/a_1059_315# 0
C18689 _0577_/a_27_297# net109 0
C18690 _0195_ net94 0
C18691 _0198_ _1061_/a_891_413# 0
C18692 _1032_/a_891_413# _0208_ 0
C18693 _1066_/a_1059_315# control0.sh 0.16384f
C18694 _0584_/a_27_297# net201 0
C18695 _1014_/a_193_47# _0465_ 0
C18696 _1062_/a_193_47# _0468_ 0
C18697 hold37/a_285_47# acc0.A\[4\] 0.00105f
C18698 _0183_ hold59/a_285_47# 0
C18699 _0995_/a_193_47# net43 0
C18700 VPWR _1030_/a_193_47# 0.29108f
C18701 clknet_1_1__leaf__0463_ _0561_/a_512_297# 0
C18702 net7 _1040_/a_193_47# 0
C18703 _0768_/a_109_297# _0308_ 0
C18704 _1061_/a_634_159# _0492_/a_27_47# 0
C18705 _1017_/a_27_47# hold72/a_49_47# 0.00835f
C18706 net109 _1022_/a_592_47# 0.00105f
C18707 _0749_/a_299_297# _0345_ 0.01589f
C18708 net182 _0181_ 0
C18709 output55/a_27_47# net116 0
C18710 acc0.A\[14\] net41 0.5259f
C18711 _0997_/a_466_413# net83 0
C18712 _0261_ _0845_/a_109_47# 0.00828f
C18713 clknet_1_0__leaf__0458_ _0263_ 0.01728f
C18714 net103 _0347_ 0
C18715 clknet_1_1__leaf__0463_ _0473_ 0
C18716 _0275_ _0399_ 0.02557f
C18717 _1021_/a_27_47# _1002_/a_27_47# 0.00132f
C18718 _0517_/a_81_21# A[9] 0
C18719 _0461_ _0240_ 0.00141f
C18720 clknet_1_1__leaf__0465_ acc0.A\[13\] 0
C18721 _0736_/a_311_297# _0181_ 0
C18722 clknet_1_0__leaf__0458_ _1047_/a_27_47# 0
C18723 hold27/a_285_47# _1046_/a_891_413# 0
C18724 _0461_ _0369_ 0.0015f
C18725 input4/a_75_212# _0187_ 0
C18726 _0194_ _0150_ 0
C18727 acc0.A\[12\] _0417_ 0
C18728 clknet_0__0457_ _0461_ 0.03025f
C18729 acc0.A\[27\] net113 0
C18730 _0133_ net122 0
C18731 _1056_/a_634_159# _1056_/a_466_413# 0.23992f
C18732 _1056_/a_193_47# _1056_/a_1059_315# 0.03405f
C18733 _1056_/a_27_47# _1056_/a_891_413# 0.03224f
C18734 _0533_/a_27_297# _0208_ 0
C18735 _1032_/a_1059_315# net17 0.01175f
C18736 _0402_ _0290_ 0
C18737 A[15] _1040_/a_27_47# 0
C18738 _0458_ _0271_ 0
C18739 _0226_ _0230_ 0
C18740 _0179_ _0464_ 0.00476f
C18741 _0113_ _0181_ 0.1707f
C18742 clknet_0__0459_ net5 0.03306f
C18743 net49 pp[21] 0.08461f
C18744 _0987_/a_381_47# _0987_/a_561_413# 0.00123f
C18745 _0987_/a_27_47# net73 0.22928f
C18746 _0987_/a_891_413# _0987_/a_975_413# 0.00851f
C18747 clknet_1_1__leaf__0459_ _0292_ 0
C18748 hold74/a_285_47# _0398_ 0
C18749 input11/a_75_212# input12/a_75_212# 0
C18750 hold47/a_391_47# _0149_ 0
C18751 _0476_ _0555_/a_51_297# 0
C18752 _0109_ _0333_ 0.00397f
C18753 _0323_ _0315_ 0.02736f
C18754 _0855_/a_81_21# net234 0.17823f
C18755 clkload2/a_268_47# clknet_1_0__leaf__0464_ 0.00294f
C18756 _0199_ _1047_/a_634_159# 0
C18757 _0182_ _1047_/a_381_47# 0
C18758 net8 _0473_ 0.02012f
C18759 acc0.A\[20\] net220 0.17065f
C18760 output54/a_27_47# pp[26] 0.15771f
C18761 _1047_/a_891_413# net218 0
C18762 _1041_/a_27_47# _0548_/a_51_297# 0
C18763 _0098_ VPWR 0.35424f
C18764 _1004_/a_634_159# _1004_/a_975_413# 0
C18765 _1004_/a_466_413# _1004_/a_561_413# 0.00772f
C18766 net125 net10 0
C18767 net47 _0986_/a_193_47# 0
C18768 _0557_/a_149_47# _1035_/a_1059_315# 0
C18769 _1027_/a_1059_315# _1008_/a_193_47# 0
C18770 _1027_/a_193_47# _1008_/a_1059_315# 0
C18771 net157 _1049_/a_1059_315# 0
C18772 _0665_/a_109_297# net5 0.00297f
C18773 net230 net139 0.00387f
C18774 clkload4/Y acc0.A\[16\] 0.00127f
C18775 acc0.A\[31\] _0712_/a_297_297# 0
C18776 _1067_/a_193_47# hold93/a_285_47# 0
C18777 _1067_/a_634_159# hold93/a_49_47# 0
C18778 _0680_/a_217_297# _0312_ 0.00271f
C18779 _0349_ net56 0.25455f
C18780 _0265_ _0264_ 0.22919f
C18781 net106 _0208_ 0
C18782 _0448_ _0843_/a_68_297# 0
C18783 clknet_1_0__leaf__0465_ _1053_/a_466_413# 0.00243f
C18784 _1029_/a_891_413# _1029_/a_975_413# 0.00851f
C18785 _1029_/a_27_47# net115 0.23069f
C18786 _1029_/a_381_47# _1029_/a_561_413# 0.00123f
C18787 net58 hold18/a_391_47# 0
C18788 comp0.B\[15\] _0177_ 0
C18789 _1019_/a_193_47# _0352_ 0
C18790 B[1] input28/a_75_212# 0.07599f
C18791 input24/a_75_212# B[5] 0.00144f
C18792 hold87/a_391_47# _0267_ 0
C18793 _0577_/a_373_47# clknet_1_0__leaf__0460_ 0
C18794 hold69/a_49_47# _0250_ 0.00282f
C18795 comp0.B\[13\] _1044_/a_27_47# 0
C18796 _0216_ control0.reset 0
C18797 VPWR _0531_/a_27_297# 0.20429f
C18798 _0269_ _0446_ 0.10573f
C18799 _0328_ _0737_/a_285_297# 0.00183f
C18800 _0817_/a_266_47# _0345_ 0.00408f
C18801 _0817_/a_266_47# _0814_/a_27_47# 0
C18802 _0346_ _0302_ 0
C18803 _0313_ clknet_0__0462_ 0.13177f
C18804 clkload0/X _1072_/a_891_413# 0
C18805 _0346_ _0795_/a_299_297# 0.00863f
C18806 hold66/a_285_47# _0219_ 0
C18807 acc0.A\[4\] _0987_/a_561_413# 0
C18808 _0399_ _0583_/a_27_297# 0
C18809 clknet_1_0__leaf__0458_ clknet_1_0__leaf__0461_ 0.00238f
C18810 _0502_/a_27_47# clknet_1_1__leaf__0457_ 0.10986f
C18811 _1000_/a_27_47# acc0.A\[18\] 0.00896f
C18812 clknet_1_0__leaf__0465_ _0144_ 0.026f
C18813 _1004_/a_1059_315# _0225_ 0
C18814 net61 _0431_ 0
C18815 _1020_/a_27_47# _0183_ 0.02947f
C18816 _1020_/a_466_413# net150 0.00113f
C18817 clknet_1_0__leaf__0463_ _0137_ 0.24726f
C18818 _1046_/a_27_47# net131 0
C18819 _0806_/a_113_297# _0806_/a_199_47# 0
C18820 net103 _1016_/a_891_413# 0.00429f
C18821 _0403_ _0277_ 0
C18822 _0096_ net43 0.0014f
C18823 _1016_/a_27_47# _1016_/a_466_413# 0.26005f
C18824 _1016_/a_193_47# _1016_/a_634_159# 0.11072f
C18825 input2/a_75_212# _0189_ 0
C18826 hold58/a_49_47# net24 0
C18827 net58 _0195_ 0.00245f
C18828 hold11/a_285_47# _1061_/a_27_47# 0
C18829 hold11/a_49_47# _1061_/a_193_47# 0
C18830 _0379_ _1023_/a_891_413# 0
C18831 clknet_1_1__leaf__0460_ hold69/a_391_47# 0.02388f
C18832 net84 clkbuf_1_1__f__0461_/a_110_47# 0.00553f
C18833 _1033_/a_891_413# comp0.B\[15\] 0
C18834 _0478_ _0976_/a_76_199# 0
C18835 _1028_/a_466_413# _1028_/a_592_47# 0.00553f
C18836 _1028_/a_634_159# _1028_/a_1017_47# 0
C18837 _0249_ _0617_/a_68_297# 0.10736f
C18838 net188 hold42/a_391_47# 0.04349f
C18839 net63 A[4] 0
C18840 net188 _1057_/a_891_413# 0
C18841 _0343_ _0996_/a_891_413# 0.00203f
C18842 _0223_ _0460_ 0
C18843 _0473_ _1042_/a_1059_315# 0
C18844 hold87/a_49_47# _0982_/a_27_47# 0
C18845 _1067_/a_27_47# control0.reset 0.01233f
C18846 _0369_ _0989_/a_975_413# 0
C18847 _1057_/a_27_47# net4 0
C18848 _0765_/a_215_47# _0460_ 0.00329f
C18849 VPWR _0990_/a_193_47# 0.31297f
C18850 A[10] net3 0
C18851 _0999_/a_27_47# _0096_ 0
C18852 _0999_/a_193_47# _0399_ 0
C18853 net119 _0131_ 0.01605f
C18854 net63 _0085_ 0.02927f
C18855 _0210_ net26 0.00707f
C18856 acc0.A\[8\] pp[3] 0
C18857 clkbuf_0__0462_/a_110_47# _0250_ 0
C18858 _0557_/a_51_297# _1037_/a_1059_315# 0
C18859 _0151_ clknet_1_0__leaf__0465_ 0.02408f
C18860 comp0.B\[10\] _0176_ 0.48132f
C18861 VPWR _1049_/a_592_47# 0
C18862 clknet_1_0__leaf__0459_ clknet_1_1__leaf__0461_ 0.10469f
C18863 net149 clkbuf_1_0__f__0461_/a_110_47# 0
C18864 clknet_0__0457_ _0465_ 0.01005f
C18865 _0556_/a_68_297# B[1] 0
C18866 net237 _0315_ 0.00151f
C18867 _0403_ _0808_/a_81_21# 0
C18868 net140 hold83/a_285_47# 0.0047f
C18869 net169 hold83/a_49_47# 0
C18870 _0473_ net10 0.04039f
C18871 net49 _0352_ 0.00172f
C18872 net20 hold51/a_285_47# 0.06078f
C18873 _1017_/a_27_47# clknet_0__0461_ 0
C18874 _0647_/a_129_47# VPWR 0.00336f
C18875 _0460_ _1006_/a_1059_315# 0.02243f
C18876 _0201_ clknet_1_1__leaf__0464_ 0.03325f
C18877 _0981_/a_109_297# _0169_ 0
C18878 _1036_/a_1059_315# _1034_/a_193_47# 0
C18879 _1036_/a_193_47# _1034_/a_1059_315# 0
C18880 VPWR _1066_/a_592_47# 0.00158f
C18881 control0.count\[3\] _0961_/a_113_297# 0
C18882 _0965_/a_47_47# _0479_ 0
C18883 net167 _1072_/a_634_159# 0
C18884 _1010_/a_466_413# clknet_1_1__leaf__0462_ 0
C18885 hold37/a_391_47# clknet_1_0__leaf__0465_ 0.00933f
C18886 control0.state\[0\] _0488_ 0.2446f
C18887 _1053_/a_891_413# A[4] 0.01143f
C18888 clkload0/a_27_47# _0183_ 0
C18889 _0271_ clkbuf_1_1__f__0458_/a_110_47# 0
C18890 comp0.B\[14\] _1044_/a_891_413# 0
C18891 _0783_/a_79_21# clknet_1_1__leaf__0461_ 0.00628f
C18892 _0730_/a_79_21# net57 0
C18893 _0517_/a_81_21# _0516_/a_27_297# 0.01185f
C18894 clknet_1_0__leaf__0463_ comp0.B\[6\] 0.00381f
C18895 _1051_/a_1059_315# _0987_/a_381_47# 0
C18896 _1056_/a_193_47# VPWR 0.3212f
C18897 net101 clknet_1_1__leaf__0457_ 0
C18898 hold14/a_391_47# clknet_1_1__leaf__0463_ 0.03064f
C18899 _0229_ _0238_ 0
C18900 _0226_ _0236_ 0.17496f
C18901 _0993_/a_592_47# _0417_ 0
C18902 _0993_/a_891_413# _0091_ 0
C18903 clkbuf_1_0__f__0459_/a_110_47# _0983_/a_193_47# 0
C18904 clknet_1_1__leaf__0459_ _0655_/a_215_53# 0
C18905 _0512_/a_27_297# _0512_/a_109_47# 0.00393f
C18906 _0770_/a_79_21# _0770_/a_297_47# 0.03259f
C18907 net58 _0852_/a_35_297# 0
C18908 _0475_ _0562_/a_68_297# 0
C18909 hold86/a_49_47# _0350_ 0.01844f
C18910 _0855_/a_299_297# VPWR 0.24739f
C18911 hold39/a_49_47# _1035_/a_1059_315# 0
C18912 net198 net129 0
C18913 _0695_/a_80_21# _0368_ 0.00677f
C18914 clknet_1_0__leaf__0465_ _1046_/a_592_47# 0
C18915 _0273_ acc0.A\[8\] 0.00785f
C18916 _0697_/a_472_297# _0319_ 0.0052f
C18917 hold85/a_49_47# _0468_ 0
C18918 _0996_/a_1059_315# net5 0.03457f
C18919 _0305_ _0345_ 0.00724f
C18920 _0346_ net6 0.02342f
C18921 net247 control0.reset 0
C18922 clknet_0_clk _1068_/a_634_159# 0.01333f
C18923 _0331_ _0319_ 0
C18924 _0349_ _0345_ 0.02383f
C18925 acc0.A\[21\] _0381_ 0.4474f
C18926 net88 acc0.A\[20\] 0
C18927 _0341_ _0220_ 0.0056f
C18928 _0998_/a_1059_315# net84 0
C18929 _1020_/a_466_413# control0.add 0
C18930 net178 _1055_/a_193_47# 0.00159f
C18931 acc0.A\[11\] _0418_ 0
C18932 net10 _0186_ 0.0695f
C18933 _0159_ _0935_/a_27_47# 0
C18934 _0097_ _0308_ 0
C18935 net89 _0369_ 0
C18936 _0159_ _1061_/a_193_47# 0.23119f
C18937 net247 _1061_/a_891_413# 0
C18938 _0183_ _0219_ 0.20898f
C18939 _0984_/a_891_413# net47 0
C18940 _0346_ _0447_ 0
C18941 _0799_/a_80_21# _0409_ 0
C18942 net231 _1065_/a_27_47# 0
C18943 _0350_ _0391_ 0.02122f
C18944 _1035_/a_193_47# net28 0
C18945 _1019_/a_891_413# _1019_/a_1017_47# 0.00617f
C18946 _1019_/a_193_47# net207 0.26141f
C18947 _0348_ _0221_ 0.20076f
C18948 _0714_/a_245_297# _0714_/a_240_47# 0
C18949 _1019_/a_634_159# net105 0
C18950 net7 _0207_ 0
C18951 clknet_1_0__leaf__0462_ hold63/a_391_47# 0.01355f
C18952 hold18/a_49_47# _0263_ 0
C18953 net51 _1005_/a_193_47# 0.0011f
C18954 hold42/a_391_47# _0155_ 0
C18955 _0098_ clknet_1_0__leaf__0459_ 0.00369f
C18956 _0467_ comp0.B\[6\] 0.01055f
C18957 _0420_ net37 0.00433f
C18958 _0403_ _0296_ 0
C18959 _0256_ _0268_ 0.00312f
C18960 _0172_ _0544_/a_149_47# 0
C18961 _0553_/a_240_47# clkbuf_1_0__f__0463_/a_110_47# 0
C18962 _0725_/a_80_21# _0333_ 0.05938f
C18963 _1051_/a_1059_315# acc0.A\[4\] 0.00196f
C18964 _0329_ _0332_ 0.32089f
C18965 _0267_ _0264_ 0.02507f
C18966 hold52/a_285_47# _0122_ 0
C18967 _0949_/a_59_75# _0161_ 0
C18968 net64 pp[3] 0
C18969 hold83/a_391_47# acc0.A\[6\] 0
C18970 _0548_/a_512_297# net174 0.00278f
C18971 _0726_/a_51_297# _0354_ 0.10341f
C18972 acc0.A\[4\] _1045_/a_381_47# 0
C18973 net8 _0497_/a_68_297# 0
C18974 hold9/a_285_47# acc0.A\[28\] 0
C18975 _1058_/a_975_413# net67 0
C18976 net43 _0395_ 0
C18977 net242 _1010_/a_466_413# 0
C18978 _0180_ _0499_/a_59_75# 0
C18979 _0533_/a_109_297# _0178_ 0
C18980 _0465_ _0844_/a_79_21# 0.00303f
C18981 net9 _0147_ 0.01989f
C18982 net175 acc0.A\[3\] 0.19705f
C18983 acc0.A\[14\] _0350_ 0.0196f
C18984 control0.state\[0\] _1064_/a_27_47# 0
C18985 hold64/a_49_47# _0461_ 0
C18986 _0130_ _1032_/a_27_47# 0.0029f
C18987 _1015_/a_193_47# _0584_/a_27_297# 0
C18988 _1015_/a_27_47# _0584_/a_109_297# 0
C18989 _0134_ B[1] 0
C18990 hold58/a_391_47# _1035_/a_1059_315# 0
C18991 hold58/a_285_47# _1035_/a_891_413# 0.00153f
C18992 _0655_/a_109_93# hold81/a_391_47# 0
C18993 _1050_/a_27_47# _0196_ 0
C18994 _1070_/a_193_47# _0976_/a_76_199# 0.00386f
C18995 _1070_/a_27_47# _0976_/a_505_21# 0.00208f
C18996 hold38/a_285_47# _1065_/a_27_47# 0.00319f
C18997 hold38/a_49_47# _1065_/a_193_47# 0
C18998 hold13/a_285_47# net8 0
C18999 net245 _0800_/a_51_297# 0.10215f
C19000 _1059_/a_27_47# _0508_/a_81_21# 0.00275f
C19001 _0536_/a_149_47# _0176_ 0
C19002 _0182_ net149 0.04796f
C19003 _0629_/a_59_75# _0447_ 0
C19004 acc0.A\[2\] _0844_/a_79_21# 0.0015f
C19005 _0195_ _0262_ 0
C19006 comp0.B\[6\] comp0.B\[0\] 0
C19007 _0902_/a_27_47# _0242_ 0
C19008 _0739_/a_79_21# _0739_/a_215_47# 0.04584f
C19009 VPWR _0998_/a_561_413# 0.00213f
C19010 _0112_ hold71/a_285_47# 0
C19011 _1020_/a_27_47# hold40/a_285_47# 0
C19012 _1020_/a_193_47# hold40/a_49_47# 0
C19013 _0127_ hold50/a_49_47# 0
C19014 hold99/a_391_47# _0091_ 0
C19015 clknet_1_0__leaf__0465_ _0987_/a_975_413# 0
C19016 _0347_ _0739_/a_510_47# 0.00602f
C19017 _0352_ _0739_/a_79_21# 0.11163f
C19018 _1029_/a_193_47# acc0.A\[28\] 0.00204f
C19019 _0990_/a_1059_315# clknet_1_1__leaf__0465_ 0
C19020 net81 _0411_ 0.00241f
C19021 _0347_ _0102_ 0.02752f
C19022 _0731_/a_81_21# _0294_ 0
C19023 _0221_ _0332_ 0.18409f
C19024 _0465_ _1048_/a_634_159# 0.00167f
C19025 _0999_/a_27_47# _0395_ 0
C19026 _0122_ net52 0.02289f
C19027 _0965_/a_377_297# VPWR 0.00595f
C19028 _1054_/a_193_47# net9 0
C19029 _0292_ _0785_/a_299_297# 0.00912f
C19030 VPWR clkbuf_1_1__f__0459_/a_110_47# 1.28449f
C19031 _0294_ _0991_/a_1017_47# 0
C19032 _0990_/a_634_159# _0088_ 0.03943f
C19033 net125 _0498_/a_245_297# 0.00141f
C19034 _0388_ _0614_/a_29_53# 0
C19035 hold81/a_391_47# _0418_ 0
C19036 acc0.A\[15\] _0219_ 0.17851f
C19037 _1002_/a_975_413# _0460_ 0
C19038 net88 _0880_/a_27_47# 0
C19039 _1002_/a_1017_47# clknet_1_0__leaf__0457_ 0
C19040 acc0.A\[2\] _1048_/a_634_159# 0
C19041 _1032_/a_1059_315# _0165_ 0
C19042 _0807_/a_68_297# _0807_/a_150_297# 0.00477f
C19043 _0793_/a_51_297# _0793_/a_240_47# 0.03076f
C19044 net64 _0273_ 0.06374f
C19045 acc0.A\[27\] hold8/a_285_47# 0
C19046 _0273_ _0621_/a_117_297# 0
C19047 net45 _0567_/a_27_297# 0
C19048 _0367_ acc0.A\[23\] 0
C19049 _0598_/a_382_297# _0237_ 0.00129f
C19050 _0230_ _0760_/a_47_47# 0
C19051 net42 _0669_/a_183_297# 0
C19052 net46 hold29/a_49_47# 0.02798f
C19053 hold65/a_49_47# _0399_ 0.04331f
C19054 _1050_/a_466_413# _0180_ 0
C19055 _0743_/a_512_297# _0368_ 0
C19056 acc0.A\[16\] _1060_/a_891_413# 0
C19057 net61 _0269_ 0
C19058 _0967_/a_487_297# _0476_ 0
C19059 _0346_ acc0.A\[0\] 0.18969f
C19060 _0260_ _0258_ 0.00101f
C19061 comp0.B\[7\] _1039_/a_634_159# 0
C19062 _0110_ hold92/a_391_47# 0
C19063 net200 _1025_/a_891_413# 0.00122f
C19064 _0216_ _0869_/a_27_47# 0
C19065 hold68/a_285_47# _0575_/a_109_297# 0
C19066 hold68/a_391_47# _0575_/a_27_297# 0.01653f
C19067 _1034_/a_634_159# comp0.B\[6\] 0.0177f
C19068 _1034_/a_27_47# _0474_ 0
C19069 _1034_/a_466_413# comp0.B\[5\] 0
C19070 _1034_/a_891_413# comp0.B\[3\] 0
C19071 hold21/a_285_47# net63 0
C19072 _0465_ _0846_/a_240_47# 0.00112f
C19073 _0438_ _0439_ 0.05325f
C19074 _1051_/a_193_47# _1051_/a_381_47# 0.09936f
C19075 _1051_/a_634_159# _1051_/a_891_413# 0.03684f
C19076 _1051_/a_27_47# _1051_/a_561_413# 0.0027f
C19077 comp0.B\[14\] _1042_/a_27_47# 0
C19078 _1056_/a_1059_315# clknet_1_1__leaf__0465_ 0
C19079 _0802_/a_145_75# VPWR 0
C19080 _0347_ _0774_/a_68_297# 0.00769f
C19081 VPWR _0438_ 0.48013f
C19082 hold15/a_49_47# hold61/a_49_47# 0
C19083 net55 _0356_ 0.00294f
C19084 pp[27] _0705_/a_59_75# 0.01046f
C19085 acc0.A\[18\] acc0.A\[19\] 0.0027f
C19086 _1070_/a_592_47# VPWR 0.0032f
C19087 _1070_/a_1059_315# control0.count\[1\] 0.11721f
C19088 _1045_/a_634_159# _1045_/a_592_47# 0
C19089 _0480_ _1069_/a_1059_315# 0
C19090 hold90/a_391_47# _0360_ 0.05353f
C19091 _1003_/a_1059_315# hold66/a_49_47# 0
C19092 hold27/a_49_47# clknet_1_0__leaf__0465_ 0.00134f
C19093 hold55/a_49_47# net106 0.05001f
C19094 net186 control0.reset 0
C19095 _0120_ net109 0.02356f
C19096 VPWR _1043_/a_1059_315# 0.39915f
C19097 VPWR _0636_/a_59_75# 0.20014f
C19098 _0217_ acc0.A\[23\] 0.1742f
C19099 _0146_ net147 0
C19100 _0678_/a_150_297# _0394_ 0
C19101 hold21/a_49_47# _0191_ 0
C19102 hold21/a_391_47# net15 0.00284f
C19103 clknet_0__0459_ _0303_ 0.00109f
C19104 clkbuf_0__0460_/a_110_47# hold90/a_285_47# 0
C19105 _0218_ _0986_/a_27_47# 0
C19106 _1028_/a_193_47# _0350_ 0
C19107 _1038_/a_27_47# _0175_ 0
C19108 clknet_1_1__leaf__0463_ _0132_ 0.00884f
C19109 _1018_/a_634_159# _0399_ 0
C19110 _0559_/a_51_297# comp0.B\[2\] 0
C19111 _1043_/a_634_159# _1043_/a_592_47# 0
C19112 net175 net157 0
C19113 hold18/a_285_47# net47 0.00195f
C19114 _0343_ acc0.A\[29\] 0.03652f
C19115 VPWR _1015_/a_27_47# 0.70931f
C19116 net191 _0347_ 0
C19117 clknet_0__0458_ _0252_ 0.00225f
C19118 acc0.A\[30\] net116 0
C19119 hold88/a_285_47# acc0.A\[8\] 0.08527f
C19120 net78 net228 0.00166f
C19121 _0554_/a_68_297# B[1] 0
C19122 input14/a_75_212# hold83/a_285_47# 0
C19123 _1004_/a_592_47# VPWR 0
C19124 _0518_/a_373_47# _0180_ 0.00112f
C19125 _0786_/a_80_21# _0369_ 0.0051f
C19126 _1054_/a_634_159# _1054_/a_1059_315# 0
C19127 _1054_/a_27_47# _1054_/a_381_47# 0.06222f
C19128 _1054_/a_193_47# _1054_/a_891_413# 0.19468f
C19129 clkbuf_1_1__f_clk/a_110_47# _0215_ 0
C19130 _1016_/a_381_47# _0352_ 0
C19131 _1071_/a_193_47# control0.count\[0\] 0.00249f
C19132 _1071_/a_891_413# clknet_1_0__leaf_clk 0.00956f
C19133 _1015_/a_27_47# _1015_/a_466_413# 0.27314f
C19134 _1015_/a_193_47# _1015_/a_634_159# 0.11072f
C19135 net224 clknet_0__0460_ 0
C19136 _0179_ _0219_ 0.09814f
C19137 _0983_/a_466_413# VPWR 0.25343f
C19138 _0730_/a_215_47# _1010_/a_634_159# 0
C19139 _0181_ _0345_ 0.14899f
C19140 _0199_ _0208_ 0
C19141 _0329_ _0738_/a_68_297# 0
C19142 _0814_/a_27_47# _0181_ 0.00411f
C19143 _0982_/a_1059_315# acc0.A\[1\] 0.00492f
C19144 net104 _0266_ 0
C19145 hold59/a_49_47# net165 0
C19146 clknet_1_1__leaf__0462_ _1027_/a_193_47# 0.01168f
C19147 pp[27] _0358_ 0
C19148 clkbuf_1_0__f__0458_/a_110_47# net58 0.01922f
C19149 _0339_ _0778_/a_68_297# 0
C19150 _0792_/a_80_21# _0405_ 0.15896f
C19151 _0987_/a_1017_47# _0085_ 0.00125f
C19152 acc0.A\[30\] hold92/a_285_47# 0.01388f
C19153 _1038_/a_27_47# _1038_/a_1059_315# 0.04861f
C19154 _1038_/a_193_47# _1038_/a_466_413# 0.0802f
C19155 _0556_/a_68_297# _1037_/a_634_159# 0
C19156 _0086_ acc0.A\[8\] 0.0413f
C19157 _0655_/a_109_93# _0303_ 0
C19158 _0283_ _0671_/a_199_47# 0
C19159 _0411_ _0797_/a_207_413# 0.07385f
C19160 _0319_ _1008_/a_27_47# 0
C19161 output48/a_27_47# VPWR 0.29849f
C19162 _0247_ clknet_1_0__leaf__0461_ 0.00796f
C19163 control0.state\[2\] _1064_/a_891_413# 0.00279f
C19164 _0856_/a_215_47# net47 0
C19165 control0.state\[0\] _1065_/a_193_47# 0
C19166 control0.state\[1\] _1065_/a_27_47# 0
C19167 hold2/a_49_47# _0181_ 0
C19168 _0340_ _0218_ 0
C19169 pp[29] hold80/a_391_47# 0.01124f
C19170 clknet_1_0__leaf__0458_ _0848_/a_27_47# 0.00396f
C19171 acc0.A\[31\] _0344_ 0
C19172 _1059_/a_561_413# _0158_ 0
C19173 pp[17] pp[18] 0.18126f
C19174 net17 _0468_ 0.04031f
C19175 _0983_/a_466_413# _0983_/a_381_47# 0.03733f
C19176 _0983_/a_193_47# _0983_/a_975_413# 0
C19177 _0983_/a_1059_315# _0983_/a_891_413# 0.31086f
C19178 comp0.B\[4\] clknet_0__0463_ 0
C19179 clknet_1_0__leaf__0465_ _1051_/a_891_413# 0.00452f
C19180 _0217_ hold60/a_49_47# 0.01409f
C19181 clknet_1_0__leaf__0458_ _0218_ 0.4019f
C19182 hold88/a_391_47# _0350_ 0
C19183 clknet_1_0__leaf__0465_ _1045_/a_561_413# 0
C19184 _0352_ _0757_/a_68_297# 0
C19185 _0758_/a_510_47# _0350_ 0.00165f
C19186 _0758_/a_215_47# _0380_ 0.0058f
C19187 net125 _0492_/a_27_47# 0.0027f
C19188 net40 _0995_/a_193_47# 0.00855f
C19189 hold29/a_285_47# VPWR 0.30391f
C19190 clknet_0__0461_ _0245_ 0.02848f
C19191 _0985_/a_634_159# net71 0
C19192 _0200_ net32 0
C19193 _0244_ _0391_ 0
C19194 acc0.A\[31\] _0709_/a_113_47# 0
C19195 _0343_ _0413_ 0
C19196 _0352_ _1025_/a_193_47# 0
C19197 _1026_/a_466_413# _0320_ 0
C19198 net8 comp0.B\[8\] 0
C19199 _0177_ _0176_ 0
C19200 net216 _0350_ 0.02746f
C19201 _0606_/a_392_297# _0237_ 0
C19202 comp0.B\[8\] net32 0
C19203 _1056_/a_193_47# hold35/a_391_47# 0.00107f
C19204 _1056_/a_466_413# hold35/a_49_47# 0.01453f
C19205 _1056_/a_634_159# hold35/a_285_47# 0
C19206 _0206_ net152 0
C19207 _0459_ _0505_/a_27_297# 0
C19208 _0466_ _1068_/a_27_47# 0.02151f
C19209 net2 net143 0
C19210 _0399_ _0114_ 0
C19211 net90 _1007_/a_193_47# 0
C19212 _0118_ net150 0
C19213 hold97/a_391_47# _0320_ 0
C19214 _0831_/a_117_297# _0369_ 0.00113f
C19215 hold33/a_285_47# _1039_/a_193_47# 0
C19216 hold33/a_391_47# _1039_/a_27_47# 0
C19217 _1003_/a_891_413# _0217_ 0.01466f
C19218 _0956_/a_32_297# comp0.B\[15\] 0.11234f
C19219 _0648_/a_277_297# _0276_ 0
C19220 net64 hold88/a_285_47# 0.00658f
C19221 _0280_ _0644_/a_377_297# 0
C19222 _1004_/a_27_47# net50 0
C19223 _0281_ _0418_ 0.11042f
C19224 _0343_ _0827_/a_109_297# 0
C19225 _0330_ _0697_/a_217_297# 0
C19226 _0317_ _0697_/a_300_47# 0.00135f
C19227 _0785_/a_81_21# _0785_/a_384_47# 0.00138f
C19228 _0244_ _0581_/a_27_297# 0.06123f
C19229 _0455_ clknet_1_0__leaf__0461_ 0
C19230 _0467_ net26 0
C19231 _1016_/a_27_47# net166 0.09523f
C19232 _1016_/a_1059_315# _1016_/a_1017_47# 0
C19233 output48/a_27_47# net48 0.22489f
C19234 clkload2/Y _1050_/a_634_159# 0
C19235 net211 acc0.A\[19\] 0.01115f
C19236 VPWR _0354_ 0.23217f
C19237 _0195_ clknet_1_0__leaf__0464_ 0.16787f
C19238 clknet_0__0459_ _0996_/a_634_159# 0
C19239 _0254_ _0369_ 0.01296f
C19240 acc0.A\[16\] _0218_ 0.05601f
C19241 control0.state\[0\] net33 0.00268f
C19242 _0439_ clknet_1_1__leaf__0465_ 0
C19243 _0361_ _0743_/a_51_297# 0
C19244 clknet_1_1__leaf__0462_ _1026_/a_1059_315# 0.01103f
C19245 net113 _1026_/a_634_159# 0
C19246 _0216_ _0705_/a_59_75# 0
C19247 _0478_ _0488_ 0.76572f
C19248 _1028_/a_381_47# acc0.A\[28\] 0
C19249 VPWR clknet_1_1__leaf__0465_ 4.65646f
C19250 _0230_ _0350_ 0
C19251 net49 _0237_ 0
C19252 _0297_ net5 0.04905f
C19253 _0277_ acc0.A\[13\] 0.10413f
C19254 net178 _0252_ 0
C19255 _0476_ hold56/a_391_47# 0
C19256 clknet_1_1__leaf__0459_ _0095_ 0.00313f
C19257 _1057_/a_592_47# _0187_ 0.00262f
C19258 _0780_/a_35_297# _0776_/a_27_47# 0
C19259 _0331_ _0333_ 0
C19260 net217 _0422_ 0.3524f
C19261 _0313_ _0687_/a_59_75# 0.03255f
C19262 _0203_ hold51/a_391_47# 0.02305f
C19263 net85 _0398_ 0
C19264 _0327_ _0701_/a_303_47# 0
C19265 pp[28] _0357_ 0
C19266 control0.state\[1\] hold12/a_285_47# 0
C19267 B[12] clknet_1_1__leaf__0464_ 0.01067f
C19268 acc0.A\[21\] _0468_ 0
C19269 clknet_0__0462_ _0321_ 0.01926f
C19270 VPWR _0215_ 0.74082f
C19271 _0514_/a_27_297# _0189_ 0.12725f
C19272 _0454_ _0265_ 0
C19273 _0179_ _0511_/a_299_297# 0.05209f
C19274 _0534_/a_299_297# _0534_/a_384_47# 0
C19275 net64 _0086_ 0.17916f
C19276 net39 _0994_/a_381_47# 0.02065f
C19277 _0283_ clkbuf_1_1__f__0459_/a_110_47# 0
C19278 _0849_/a_297_297# _0347_ 0
C19279 _0134_ _1037_/a_634_159# 0
C19280 _1032_/a_466_413# _0352_ 0
C19281 hold62/a_285_47# hold62/a_391_47# 0.41909f
C19282 _0984_/a_27_47# _0450_ 0
C19283 _1059_/a_561_413# acc0.A\[14\] 0.00167f
C19284 _0538_/a_51_297# _0142_ 0
C19285 _0538_/a_149_47# net20 0.00472f
C19286 net236 _1068_/a_27_47# 0
C19287 hold42/a_49_47# acc0.A\[11\] 0.03227f
C19288 _1041_/a_561_413# net7 0.00214f
C19289 _0554_/a_68_297# _1035_/a_891_413# 0
C19290 control0.state\[2\] hold84/a_49_47# 0
C19291 clknet_1_1__leaf__0459_ _1057_/a_634_159# 0
C19292 _0780_/a_35_297# _0219_ 0
C19293 _0216_ _0460_ 0.03528f
C19294 _1057_/a_466_413# acc0.A\[11\] 0
C19295 _0593_/a_113_47# net50 0
C19296 _0412_ net5 0.02344f
C19297 hold54/a_285_47# _0130_ 0.00433f
C19298 _0499_/a_59_75# _0495_/a_150_297# 0
C19299 VPWR _0693_/a_68_297# 0.17036f
C19300 _1048_/a_27_47# _0509_/a_27_47# 0
C19301 net193 net32 0
C19302 hold76/a_49_47# _0183_ 0
C19303 _0233_ _0754_/a_51_297# 0.00224f
C19304 _0753_/a_79_21# _0377_ 0.14262f
C19305 _1056_/a_891_413# _1056_/a_1017_47# 0.00617f
C19306 _1056_/a_193_47# net182 0.24369f
C19307 _0323_ _0691_/a_150_297# 0
C19308 hold74/a_49_47# _0306_ 0
C19309 _1004_/a_891_413# hold68/a_285_47# 0.00178f
C19310 _0734_/a_47_47# _1009_/a_193_47# 0
C19311 _1054_/a_561_413# VPWR 0.0031f
C19312 _0643_/a_103_199# _0258_ 0.00298f
C19313 _0315_ _0320_ 0.00194f
C19314 clknet_0_clk _0564_/a_68_297# 0
C19315 _0517_/a_81_21# _0190_ 0.19198f
C19316 _0517_/a_384_47# net16 0
C19317 _0305_ _0394_ 0.00176f
C19318 _0108_ _0195_ 0
C19319 clknet_1_1__leaf__0465_ output62/a_27_47# 0
C19320 acc0.A\[5\] _0987_/a_1059_315# 0.03377f
C19321 _1051_/a_975_413# net73 0
C19322 _0200_ net10 0.6659f
C19323 net59 _0588_/a_113_47# 0
C19324 clknet_1_0__leaf__0459_ _1015_/a_27_47# 0.00138f
C19325 _0802_/a_59_75# _0286_ 0
C19326 _0163_ _1065_/a_634_159# 0.03812f
C19327 _0389_ _0243_ 0.58995f
C19328 _1038_/a_381_47# VPWR 0.07664f
C19329 _0457_ _0216_ 0.01695f
C19330 _0707_/a_544_297# _0336_ 0
C19331 _1041_/a_381_47# A[15] 0
C19332 _0573_/a_27_47# net23 0
C19333 hold39/a_285_47# _0133_ 0.02964f
C19334 _0368_ clknet_1_0__leaf__0460_ 0.00277f
C19335 net104 _0612_/a_59_75# 0
C19336 _0695_/a_80_21# clknet_0__0460_ 0.00106f
C19337 clknet_0_clk clknet_1_1__leaf_clk 0.04126f
C19338 _1067_/a_27_47# _0460_ 0.00114f
C19339 _1067_/a_634_159# clknet_1_0__leaf__0457_ 0.01085f
C19340 comp0.B\[8\] net10 0
C19341 input4/a_75_212# clknet_1_1__leaf__0465_ 0.00712f
C19342 hold36/a_49_47# VPWR 0.31574f
C19343 net203 _0956_/a_32_297# 0.00127f
C19344 _0446_ clkbuf_0__0458_/a_110_47# 0.00325f
C19345 _0983_/a_466_413# clknet_1_0__leaf__0459_ 0
C19346 acc0.A\[7\] net12 0
C19347 clknet_1_0__leaf__0460_ _0618_/a_215_47# 0.00269f
C19348 _0695_/a_300_47# _0250_ 0.00117f
C19349 _0118_ control0.add 0
C19350 _0225_ _0617_/a_68_297# 0
C19351 _0374_ net241 0.10445f
C19352 _0181_ net52 0
C19353 clkbuf_1_1__f__0463_/a_110_47# _0563_/a_240_47# 0.00227f
C19354 clknet_0__0463_ _0563_/a_245_297# 0
C19355 _0241_ _0616_/a_493_297# 0
C19356 _0760_/a_47_47# _0760_/a_377_297# 0.00899f
C19357 hold31/a_285_47# _0988_/a_27_47# 0.00104f
C19358 _0819_/a_81_21# _0181_ 0.00251f
C19359 VPWR _0452_ 0.22797f
C19360 pp[17] _0567_/a_109_47# 0
C19361 net56 _1030_/a_193_47# 0
C19362 _0146_ _0186_ 0
C19363 _0627_/a_109_93# _0252_ 0
C19364 _1031_/a_193_47# _1030_/a_634_159# 0
C19365 _1031_/a_466_413# _1030_/a_27_47# 0
C19366 _1031_/a_27_47# _1030_/a_466_413# 0
C19367 _0714_/a_149_47# _0111_ 0.0013f
C19368 VPWR _0567_/a_27_297# 0.17167f
C19369 net35 _1071_/a_975_413# 0
C19370 _1008_/a_466_413# net244 0
C19371 _0457_ _1067_/a_27_47# 0
C19372 control0.count\[3\] _0483_ 0.01451f
C19373 _0467_ hold84/a_285_47# 0.00115f
C19374 _0180_ _0270_ 0.00591f
C19375 net245 _0277_ 0
C19376 _0298_ acc0.A\[13\] 0.02523f
C19377 _1032_/a_193_47# comp0.B\[15\] 0
C19378 comp0.B\[7\] net147 0
C19379 _0180_ _0987_/a_466_413# 0
C19380 _0782_/a_27_47# _1014_/a_381_47# 0
C19381 clknet_1_0__leaf__0458_ _0112_ 0.00107f
C19382 _1038_/a_193_47# _0550_/a_240_47# 0
C19383 _0382_ hold3/a_285_47# 0
C19384 _0260_ net72 0
C19385 _0712_/a_297_297# _0708_/a_68_297# 0.00389f
C19386 _0138_ net174 0.05835f
C19387 _0343_ _0995_/a_975_413# 0
C19388 _1014_/a_592_47# clknet_1_0__leaf__0461_ 0
C19389 net76 clkbuf_1_1__f__0458_/a_110_47# 0
C19390 _1025_/a_27_47# _1025_/a_1059_315# 0.04875f
C19391 _1025_/a_193_47# _1025_/a_466_413# 0.07855f
C19392 _0359_ _1006_/a_27_47# 0
C19393 net49 _1005_/a_27_47# 0.02096f
C19394 _0355_ net227 0.20312f
C19395 clknet_1_1__leaf__0463_ net25 0.0087f
C19396 _0770_/a_79_21# _0462_ 0.00227f
C19397 clkbuf_1_0__f__0461_/a_110_47# net206 0.01018f
C19398 _1012_/a_193_47# _0345_ 0
C19399 _0858_/a_27_47# net218 0.00244f
C19400 _0269_ _0431_ 0.1075f
C19401 hold82/a_391_47# _0345_ 0.00126f
C19402 _0116_ _0350_ 0
C19403 comp0.B\[1\] _1032_/a_381_47# 0
C19404 _0296_ acc0.A\[13\] 0
C19405 _0179_ _1055_/a_1059_315# 0.00521f
C19406 _0087_ net75 0.00269f
C19407 net45 _0398_ 0.03726f
C19408 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0465_/a_110_47# 0.00208f
C19409 _0274_ _0434_ 0.36271f
C19410 hold55/a_391_47# net202 0.12947f
C19411 input19/a_75_212# _0541_/a_68_297# 0.00119f
C19412 _1055_/a_27_47# _0181_ 0
C19413 hold28/a_49_47# _0195_ 0.00824f
C19414 VPWR _0522_/a_109_297# 0.19764f
C19415 _1070_/a_193_47# _0488_ 0.00243f
C19416 _1070_/a_27_47# _0466_ 0.0016f
C19417 VPWR _0976_/a_76_199# 0.11942f
C19418 hold31/a_391_47# clknet_1_1__leaf__0458_ 0.00376f
C19419 net193 net10 0.02633f
C19420 _0800_/a_51_297# VPWR 0.52835f
C19421 net82 _0369_ 0
C19422 comp0.B\[0\] hold84/a_285_47# 0.00337f
C19423 _0347_ hold72/a_391_47# 0
C19424 net40 _0093_ 0.00162f
C19425 _1059_/a_891_413# net228 0
C19426 _0432_ _0270_ 0
C19427 _0443_ _0256_ 0
C19428 _0999_/a_193_47# _0306_ 0
C19429 _1046_/a_466_413# net10 0.03319f
C19430 _0467_ _1065_/a_561_413# 0.00214f
C19431 _0396_ _0778_/a_150_297# 0
C19432 hold86/a_391_47# clknet_1_0__leaf__0458_ 0
C19433 input31/a_75_212# net153 0
C19434 clknet_1_1__leaf__0463_ _0477_ 0
C19435 _1003_/a_27_47# _0486_ 0
C19436 _1003_/a_193_47# control0.state\[2\] 0.00264f
C19437 _0465_ net134 0.00172f
C19438 _1021_/a_1059_315# _0369_ 0
C19439 control0.count\[3\] control0.count\[1\] 0
C19440 _0996_/a_634_159# _0996_/a_1059_315# 0
C19441 _0996_/a_27_47# _0996_/a_381_47# 0.06222f
C19442 _0996_/a_193_47# _0996_/a_891_413# 0.19489f
C19443 _0174_ _0498_/a_149_47# 0.02736f
C19444 VPWR _0829_/a_27_47# 0.00489f
C19445 _0999_/a_1017_47# _0345_ 0
C19446 clknet_1_0__leaf__0464_ _1048_/a_193_47# 0.00249f
C19447 acc0.A\[2\] net134 0
C19448 hold10/a_391_47# clknet_1_1__leaf__0457_ 0
C19449 _0793_/a_512_297# _0095_ 0
C19450 _0646_/a_377_297# net5 0.00379f
C19451 acc0.A\[16\] _1017_/a_975_413# 0.0014f
C19452 hold56/a_285_47# net203 0.01298f
C19453 _0494_/a_27_47# _0171_ 0
C19454 hold57/a_49_47# _0473_ 0.01244f
C19455 _0559_/a_149_47# _0175_ 0
C19456 hold76/a_391_47# _0248_ 0
C19457 hold8/a_49_47# _1027_/a_27_47# 0.00166f
C19458 clknet_1_0__leaf__0459_ clknet_1_1__leaf__0465_ 0
C19459 VPWR _0996_/a_561_413# 0.00309f
C19460 _0344_ _0999_/a_27_47# 0
C19461 _0317_ _1008_/a_193_47# 0
C19462 _0275_ _0346_ 0.12625f
C19463 _0465_ _0084_ 0
C19464 comp0.B\[7\] net125 0
C19465 _0726_/a_512_297# acc0.A\[29\] 0
C19466 _1059_/a_1059_315# _0347_ 0
C19467 _0454_ _0267_ 0
C19468 hold33/a_285_47# _1041_/a_1059_315# 0.00197f
C19469 _0243_ _0266_ 0
C19470 _1051_/a_193_47# acc0.A\[5\] 0
C19471 _1051_/a_1059_315# _0149_ 0
C19472 _1051_/a_891_413# net137 0
C19473 hold22/a_391_47# _1054_/a_193_47# 0
C19474 _1045_/a_891_413# _1044_/a_891_413# 0.0022f
C19475 _0220_ acc0.A\[30\] 0.60024f
C19476 _0115_ _0240_ 0
C19477 _0762_/a_215_47# net51 0.00387f
C19478 _0992_/a_1059_315# acc0.A\[10\] 0.07857f
C19479 _1051_/a_561_413# net131 0
C19480 _0292_ clkbuf_1_1__f__0465_/a_110_47# 0.02483f
C19481 _0288_ _0218_ 0
C19482 net62 _0986_/a_561_413# 0
C19483 _0369_ _0115_ 0.00812f
C19484 clknet_1_1__leaf__0461_ _0345_ 0.01205f
C19485 _0730_/a_79_21# clkbuf_1_1__f__0460_/a_110_47# 0.01161f
C19486 net78 _0090_ 0.26237f
C19487 net203 _1032_/a_193_47# 0
C19488 _0283_ clknet_1_1__leaf__0465_ 0
C19489 net23 _1067_/a_592_47# 0.00261f
C19490 clknet_0__0465_ _0090_ 0
C19491 _0311_ _0346_ 0
C19492 _0101_ hold66/a_285_47# 0.08922f
C19493 _0787_/a_80_21# _0993_/a_193_47# 0.00344f
C19494 _0787_/a_209_297# _0993_/a_27_47# 0
C19495 _0399_ _0990_/a_466_413# 0.03247f
C19496 _0299_ input6/a_75_212# 0
C19497 hold47/a_49_47# clknet_1_1__leaf__0464_ 0
C19498 _0249_ net241 0
C19499 net245 _0298_ 0
C19500 net191 _0106_ 0
C19501 _0227_ _0232_ 0
C19502 _1002_/a_1059_315# net240 0
C19503 _1002_/a_193_47# _0165_ 0
C19504 _0984_/a_381_47# _0158_ 0
C19505 net104 _0399_ 0.18305f
C19506 _0369_ _0796_/a_297_297# 0.00326f
C19507 control0.sh net29 0.00776f
C19508 _0714_/a_51_297# _1013_/a_27_47# 0.00151f
C19509 _1060_/a_27_47# net229 0
C19510 _1060_/a_381_47# _0506_/a_81_21# 0
C19511 clknet_1_1__leaf__0459_ _0672_/a_510_47# 0
C19512 hold58/a_49_47# _0135_ 0
C19513 clknet_1_1__leaf__0460_ _0776_/a_27_47# 0.00118f
C19514 _1003_/a_634_159# _0467_ 0
C19515 _0181_ _0394_ 0
C19516 net211 net1 0
C19517 _0458_ _0529_/a_373_47# 0
C19518 clkbuf_0__0464_/a_110_47# net20 0.0051f
C19519 _1016_/a_381_47# hold72/a_285_47# 0
C19520 _1030_/a_193_47# _0345_ 0.01459f
C19521 _0662_/a_81_21# _0817_/a_81_21# 0
C19522 clknet_1_0__leaf__0463_ _1040_/a_466_413# 0
C19523 hold3/a_285_47# _1005_/a_634_159# 0
C19524 clknet_0__0464_ _0138_ 0
C19525 _1021_/a_592_47# net88 0.00152f
C19526 _0218_ _0247_ 0.04883f
C19527 _1032_/a_634_159# _1032_/a_381_47# 0
C19528 net9 acc0.A\[6\] 0.46383f
C19529 _1054_/a_1059_315# net140 0
C19530 _1054_/a_466_413# net169 0.04709f
C19531 _1015_/a_27_47# _0113_ 0.09113f
C19532 _1015_/a_1059_315# _1015_/a_1017_47# 0
C19533 _0251_ output63/a_27_47# 0.01261f
C19534 output42/a_27_47# hold98/a_285_47# 0
C19535 _1038_/a_466_413# net29 0
C19536 net113 _0689_/a_68_297# 0
C19537 _0604_/a_113_47# _0346_ 0
C19538 clkbuf_1_0__f__0457_/a_110_47# _0218_ 0.002f
C19539 _0569_/a_27_297# _0569_/a_109_297# 0.17136f
C19540 _0497_/a_68_297# _0492_/a_27_47# 0.00928f
C19541 _0557_/a_240_47# _0208_ 0.06108f
C19542 _0108_ _1010_/a_891_413# 0
C19543 clknet_1_1__leaf__0460_ _0219_ 0.1421f
C19544 control0.state\[2\] _0471_ 0.15604f
C19545 _0753_/a_465_47# clknet_1_0__leaf__0460_ 0
C19546 _1051_/a_27_47# _0180_ 0.03589f
C19547 hold33/a_49_47# net147 0
C19548 acc0.A\[7\] pp[5] 0.0065f
C19549 _0343_ _1031_/a_975_413# 0
C19550 _0400_ _0408_ 0.00114f
C19551 _1014_/a_466_413# net149 0.02842f
C19552 _1038_/a_891_413# _1038_/a_1017_47# 0.00617f
C19553 _1038_/a_193_47# net172 0.22882f
C19554 _1038_/a_634_159# net124 0
C19555 _0211_ _1037_/a_381_47# 0
C19556 _0472_ net7 0
C19557 net33 _1066_/a_193_47# 0.16692f
C19558 clknet_1_1__leaf__0460_ _0728_/a_59_75# 0
C19559 _0729_/a_68_297# _0701_/a_80_21# 0
C19560 hold35/a_391_47# clknet_1_1__leaf__0465_ 0
C19561 hold46/a_391_47# _0548_/a_51_297# 0
C19562 _0731_/a_81_21# _0371_ 0
C19563 _0731_/a_299_297# net216 0
C19564 _0172_ _1043_/a_466_413# 0
C19565 _1067_/a_891_413# net107 0
C19566 _1067_/a_561_413# clknet_1_0__leaf__0461_ 0
C19567 _0464_ _0171_ 0.00543f
C19568 _0476_ _0496_/a_27_47# 0
C19569 _0183_ net58 0
C19570 _0442_ _0087_ 0
C19571 _0661_/a_109_297# _0345_ 0
C19572 _0603_/a_68_297# _0346_ 0.00125f
C19573 _0346_ hold73/a_391_47# 0
C19574 clknet_1_0__leaf__0465_ _1044_/a_381_47# 0.0014f
C19575 pp[1] net141 0.00246f
C19576 comp0.B\[7\] _0473_ 0.08099f
C19577 net167 _0486_ 0
C19578 hold16/a_285_47# _1030_/a_27_47# 0.00287f
C19579 hold36/a_285_47# hold36/a_391_47# 0.41909f
C19580 net11 _0142_ 0
C19581 net58 output63/a_27_47# 0
C19582 _0289_ _0673_/a_337_297# 0.00684f
C19583 _0625_/a_59_75# _0369_ 0.00103f
C19584 _0287_ _0673_/a_253_297# 0
C19585 acc0.A\[21\] _0762_/a_79_21# 0
C19586 net61 clkbuf_0__0458_/a_110_47# 0.00427f
C19587 _0997_/a_27_47# net43 0.04572f
C19588 net9 _0523_/a_384_47# 0
C19589 _0263_ _0448_ 0
C19590 _0216_ _0614_/a_29_53# 0.00198f
C19591 net245 _0995_/a_1017_47# 0
C19592 _0983_/a_27_47# acc0.A\[18\] 0
C19593 _0457_ net100 0
C19594 net66 acc0.A\[8\] 0.5117f
C19595 _0455_ _0218_ 0.01432f
C19596 _0461_ hold40/a_391_47# 0.0022f
C19597 clknet_1_1__leaf__0460_ _1008_/a_634_159# 0.00147f
C19598 clknet_1_0__leaf__0465_ _0528_/a_81_21# 0.00109f
C19599 _0457_ net186 0
C19600 hold45/a_391_47# net4 0.01453f
C19601 _0997_/a_381_47# net42 0.01434f
C19602 hold37/a_391_47# _0148_ 0
C19603 _0371_ _1006_/a_193_47# 0.01087f
C19604 net216 _1006_/a_634_159# 0
C19605 _0726_/a_51_297# _0353_ 0
C19606 net106 _1032_/a_466_413# 0
C19607 _0264_ _0347_ 0
C19608 acc0.A\[12\] _1058_/a_1059_315# 0.11658f
C19609 _0459_ _0184_ 0
C19610 hold32/a_391_47# _1055_/a_193_47# 0
C19611 hold32/a_285_47# _1055_/a_634_159# 0
C19612 _1048_/a_891_413# _1047_/a_891_413# 0
C19613 _0452_ _0453_ 0.05645f
C19614 _0767_/a_145_75# _0387_ 0
C19615 _0101_ _0183_ 0.0216f
C19616 _1054_/a_891_413# acc0.A\[6\] 0
C19617 _1000_/a_27_47# _0461_ 0.02025f
C19618 VPWR _0955_/a_304_297# 0.00579f
C19619 _0520_/a_109_297# net12 0
C19620 _0643_/a_103_199# net72 0.00682f
C19621 _0954_/a_114_297# comp0.B\[10\] 0
C19622 _0294_ _0505_/a_109_47# 0
C19623 _0244_ _0116_ 0.09641f
C19624 _0578_/a_109_297# _0352_ 0.0069f
C19625 _0421_ acc0.A\[10\] 0
C19626 net182 clknet_1_1__leaf__0465_ 0.00289f
C19627 hold32/a_49_47# net181 0
C19628 _0616_/a_292_297# _0246_ 0
C19629 _1036_/a_634_159# _0175_ 0.00549f
C19630 _0240_ _0614_/a_111_297# 0.00108f
C19631 _0181_ hold93/a_49_47# 0.04898f
C19632 _0534_/a_81_21# acc0.A\[1\] 0
C19633 net113 net112 0.00358f
C19634 _0991_/a_27_47# _0991_/a_193_47# 0.97064f
C19635 net58 acc0.A\[15\] 0.05929f
C19636 _0998_/a_592_47# _0399_ 0
C19637 _0998_/a_975_413# _0096_ 0
C19638 _0567_/a_27_297# _0567_/a_373_47# 0.01338f
C19639 _0313_ _0352_ 0.00142f
C19640 _0263_ _0444_ 0
C19641 _0241_ _0771_/a_27_413# 0.00213f
C19642 _0370_ _0350_ 0.04836f
C19643 hold23/a_49_47# _0180_ 0.0406f
C19644 _0243_ _0612_/a_59_75# 0
C19645 hold54/a_391_47# comp0.B\[15\] 0.04654f
C19646 _0502_/a_27_47# net135 0
C19647 acc0.A\[22\] hold4/a_391_47# 0.03089f
C19648 _0183_ hold4/a_285_47# 0.0856f
C19649 net160 _0957_/a_32_297# 0.05516f
C19650 _1008_/a_381_47# hold50/a_285_47# 0
C19651 _1052_/a_891_413# net11 0.01996f
C19652 acc0.A\[8\] _0350_ 0.24874f
C19653 net202 _0352_ 0
C19654 _0982_/a_193_47# _1014_/a_891_413# 0
C19655 _0982_/a_634_159# _1014_/a_1059_315# 0
C19656 net178 pp[8] 0
C19657 _0684_/a_59_75# _0360_ 0
C19658 net55 _0737_/a_35_297# 0
C19659 hold27/a_285_47# _0176_ 0
C19660 _0195_ _1017_/a_381_47# 0.01241f
C19661 net160 _1035_/a_1017_47# 0
C19662 clknet_1_1__leaf__0463_ _0352_ 0
C19663 net189 acc0.A\[11\] 0.02195f
C19664 _0618_/a_215_47# hold94/a_285_47# 0
C19665 _0251_ _0179_ 0.00125f
C19666 _0983_/a_27_47# hold59/a_49_47# 0
C19667 control0.count\[2\] clkbuf_1_0__f_clk/a_110_47# 0.03202f
C19668 _0677_/a_285_47# _0306_ 0.00105f
C19669 _0234_ clknet_1_0__leaf__0460_ 0.26222f
C19670 _1057_/a_381_47# VPWR 0.07542f
C19671 comp0.B\[4\] _1034_/a_1017_47# 0
C19672 clknet_1_1__leaf__0460_ _0746_/a_81_21# 0
C19673 clkbuf_1_1__f__0462_/a_110_47# _1008_/a_466_413# 0
C19674 _0233_ _0219_ 0.01415f
C19675 _0579_/a_27_297# VPWR 0.18581f
C19676 hold35/a_49_47# hold35/a_285_47# 0.22264f
C19677 _0991_/a_193_47# _0350_ 0
C19678 _0548_/a_51_297# net153 0
C19679 hold13/a_285_47# hold57/a_49_47# 0.03151f
C19680 _0174_ _0540_/a_51_297# 0.2145f
C19681 acc0.A\[27\] hold9/a_49_47# 0
C19682 _0362_ _1009_/a_466_413# 0.00478f
C19683 _0222_ _0606_/a_392_297# 0
C19684 _0687_/a_59_75# _0321_ 0.00105f
C19685 _0343_ hold78/a_285_47# 0.03758f
C19686 _0315_ _1007_/a_1059_315# 0
C19687 _0366_ _1007_/a_891_413# 0.06281f
C19688 clknet_0__0464_ net134 0
C19689 comp0.B\[10\] _0540_/a_512_297# 0
C19690 _0621_/a_35_297# acc0.A\[8\] 0
C19691 VPWR _0398_ 0.31859f
C19692 hold11/a_285_47# _0174_ 0
C19693 _0722_/a_79_21# _0347_ 0.12974f
C19694 _0671_/a_199_47# _0345_ 0
C19695 _0976_/a_76_199# _0976_/a_535_374# 0
C19696 _1050_/a_891_413# clknet_1_1__leaf__0464_ 0.00155f
C19697 _1001_/a_466_413# _0580_/a_27_297# 0
C19698 _1001_/a_634_159# _0580_/a_109_297# 0
C19699 _0800_/a_51_297# _0800_/a_149_47# 0.02487f
C19700 clknet_1_0__leaf__0460_ clknet_0__0460_ 0.00539f
C19701 hold57/a_391_47# _0174_ 0.04412f
C19702 net35 _1072_/a_1017_47# 0
C19703 acc0.A\[29\] _0568_/a_27_297# 0.06634f
C19704 _0855_/a_299_297# _0345_ 0.01078f
C19705 _1017_/a_891_413# _0369_ 0
C19706 clkbuf_0__0463_/a_110_47# _0496_/a_27_47# 0
C19707 _0225_ _1023_/a_466_413# 0
C19708 _1052_/a_891_413# hold7/a_391_47# 0
C19709 _1002_/a_27_47# _0352_ 0
C19710 pp[17] _1031_/a_193_47# 0
C19711 _0183_ _0262_ 0
C19712 net49 _0222_ 0
C19713 _0179_ net58 0.01947f
C19714 hold33/a_49_47# _0473_ 0.00846f
C19715 _0607_/a_109_47# _0352_ 0.00163f
C19716 _0369_ net146 0
C19717 _0965_/a_285_47# _0466_ 0.0441f
C19718 _0179_ hold7/a_49_47# 0.00682f
C19719 hold14/a_391_47# _0134_ 0
C19720 _0760_/a_285_47# _0382_ 0.04387f
C19721 _0350_ _0380_ 0.01743f
C19722 net178 _0988_/a_891_413# 0.04568f
C19723 _0458_ _0845_/a_109_47# 0.0178f
C19724 _0183_ _0582_/a_109_297# 0.01661f
C19725 _0180_ A[4] 0
C19726 _0983_/a_891_413# _0399_ 0.04365f
C19727 net51 _1022_/a_1059_315# 0.01703f
C19728 _0183_ net23 0
C19729 net205 _0213_ 0
C19730 VPWR _0277_ 2.9282f
C19731 clknet_1_0__leaf__0463_ _1061_/a_381_47# 0.01913f
C19732 hold68/a_391_47# net176 0.00593f
C19733 net215 hold29/a_391_47# 0
C19734 hold42/a_49_47# A[12] 0
C19735 _0430_ clknet_0__0465_ 0.00328f
C19736 _0835_/a_78_199# _0835_/a_292_297# 0.01295f
C19737 _0975_/a_59_75# clknet_1_0__leaf_clk 0
C19738 _0180_ _0085_ 0
C19739 net76 _0290_ 0.00252f
C19740 hold78/a_49_47# net60 0.33161f
C19741 hold65/a_49_47# _0346_ 0
C19742 net123 _0207_ 0
C19743 _0344_ _0708_/a_68_297# 0
C19744 _0218_ pp[13] 0
C19745 _0195_ _0581_/a_27_297# 0
C19746 _1025_/a_891_413# _1025_/a_1017_47# 0.00617f
C19747 net64 _0350_ 0
C19748 _0369_ pp[3] 0
C19749 net78 _0401_ 0
C19750 hold69/a_285_47# _0462_ 0.01111f
C19751 _0973_/a_27_297# _1067_/a_1059_315# 0
C19752 _0973_/a_109_297# _1067_/a_466_413# 0
C19753 clknet_0__0465_ _0401_ 0.08032f
C19754 _0195_ clkbuf_1_0__f__0464_/a_110_47# 0.01983f
C19755 hold65/a_49_47# net65 0.32604f
C19756 _0982_/a_1059_315# _0216_ 0
C19757 pp[15] acc0.A\[13\] 0
C19758 clk _0972_/a_250_297# 0
C19759 VPWR _0488_ 0.70768f
C19760 comp0.B\[7\] _0497_/a_68_297# 0
C19761 _1001_/a_27_47# control0.add 0.01024f
C19762 _0966_/a_109_297# _0483_ 0.01121f
C19763 _0369_ net223 0.10041f
C19764 _0516_/a_109_47# clknet_1_1__leaf__0465_ 0.00311f
C19765 hold49/a_391_47# comp0.B\[11\] 0
C19766 hold49/a_285_47# comp0.B\[12\] 0.02112f
C19767 clknet_0__0457_ net223 0
C19768 clkbuf_1_0__f__0457_/a_110_47# _0099_ 0.00342f
C19769 comp0.B\[5\] _0175_ 0.02118f
C19770 comp0.B\[3\] _0215_ 0
C19771 _0238_ _1006_/a_27_47# 0
C19772 acc0.A\[11\] _0417_ 0
C19773 _0119_ _1067_/a_27_47# 0
C19774 _0183_ net35 0
C19775 _0516_/a_27_297# _0088_ 0
C19776 net16 _0990_/a_891_413# 0
C19777 _0432_ _0085_ 0
C19778 _0182_ comp0.B\[15\] 0.00119f
C19779 _0262_ acc0.A\[15\] 0.0013f
C19780 net205 _0212_ 0.14494f
C19781 VPWR _0808_/a_81_21# 0.54063f
C19782 _1055_/a_193_47# _0153_ 0
C19783 _0315_ clkbuf_1_0__f__0462_/a_110_47# 0.14357f
C19784 _0998_/a_466_413# _0219_ 0
C19785 _0218_ _0779_/a_297_297# 0
C19786 hold57/a_391_47# _0208_ 0.03475f
C19787 _0822_/a_109_297# _0430_ 0.01334f
C19788 hold77/a_49_47# VPWR 0.33902f
C19789 _0801_/a_113_47# _0414_ 0.00937f
C19790 net64 _0621_/a_35_297# 0.24294f
C19791 _0621_/a_35_297# _0621_/a_117_297# 0.00641f
C19792 _0402_ _0993_/a_193_47# 0
C19793 _0243_ _0399_ 0
C19794 _0581_/a_109_47# _0247_ 0
C19795 _0343_ acc0.A\[23\] 0.08913f
C19796 net168 output63/a_27_47# 0
C19797 _0129_ net60 0.01744f
C19798 _0217_ clknet_1_0__leaf__0461_ 0.09926f
C19799 comp0.B\[6\] control0.sh 0.17016f
C19800 _0462_ _0617_/a_68_297# 0.00304f
C19801 hold53/a_285_47# _0124_ 0
C19802 net1 hold84/a_285_47# 0
C19803 hold63/a_285_47# acc0.A\[25\] 0.00659f
C19804 hold68/a_49_47# hold68/a_391_47# 0.00188f
C19805 clkbuf_1_1__f__0459_/a_110_47# _0345_ 0.02737f
C19806 _0137_ net157 0
C19807 _0158_ _0505_/a_373_47# 0
C19808 _1052_/a_891_413# clknet_1_1__leaf__0458_ 0
C19809 hold79/a_285_47# _0978_/a_109_297# 0
C19810 hold79/a_391_47# _0978_/a_27_297# 0
C19811 acc0.A\[16\] _1016_/a_1059_315# 0.14678f
C19812 _0317_ _0318_ 0.15265f
C19813 _0273_ _0369_ 0
C19814 clknet_1_0__leaf__0463_ _1039_/a_381_47# 0
C19815 _1057_/a_592_47# clknet_1_1__leaf__0465_ 0
C19816 VPWR _1036_/a_975_413# 0.00483f
C19817 _1050_/a_27_47# _0524_/a_27_297# 0
C19818 output43/a_27_47# net43 0.17911f
C19819 hold48/a_49_47# clkbuf_1_1__f__0464_/a_110_47# 0.00143f
C19820 hold24/a_391_47# _0136_ 0.02116f
C19821 net98 _0306_ 0
C19822 clknet_1_1__leaf__0461_ _0394_ 0.00655f
C19823 _0536_/a_51_297# _0138_ 0.00198f
C19824 _0536_/a_240_47# net173 0
C19825 clknet_0__0457_ _0982_/a_891_413# 0
C19826 _1044_/a_1059_315# _1044_/a_891_413# 0.31086f
C19827 _1044_/a_193_47# _1044_/a_975_413# 0
C19828 _1044_/a_466_413# _1044_/a_381_47# 0.03733f
C19829 _0654_/a_27_413# _0808_/a_81_21# 0
C19830 _1065_/a_27_47# _0564_/a_68_297# 0.00173f
C19831 _0109_ acc0.A\[29\] 0.07084f
C19832 net101 _0584_/a_109_47# 0
C19833 VPWR _0353_ 0.2244f
C19834 VPWR _0150_ 0.33089f
C19835 _1038_/a_1059_315# comp0.B\[5\] 0
C19836 _1038_/a_466_413# comp0.B\[6\] 0.00182f
C19837 hold41/a_285_47# _1058_/a_193_47# 0.0028f
C19838 hold41/a_391_47# _1058_/a_27_47# 0
C19839 _0172_ _0522_/a_27_297# 0
C19840 _0815_/a_113_297# _0425_ 0.09112f
C19841 _0815_/a_199_47# _0401_ 0
C19842 acc0.A\[14\] _0852_/a_35_297# 0
C19843 hold22/a_49_47# net169 0
C19844 net131 _1044_/a_975_413# 0
C19845 VPWR _0743_/a_51_297# 0.46588f
C19846 net149 _1048_/a_1059_315# 0
C19847 net18 _0541_/a_68_297# 0.00468f
C19848 _0302_ net238 0
C19849 output36/a_27_47# _1038_/a_193_47# 0
C19850 _0410_ _0795_/a_81_21# 0.11556f
C19851 clknet_1_1__leaf_clk _1065_/a_27_47# 0.31118f
C19852 _0999_/a_193_47# _0778_/a_68_297# 0
C19853 clkload3/Y _0306_ 0
C19854 _0819_/a_81_21# _0990_/a_193_47# 0
C19855 clknet_1_1__leaf__0459_ _0219_ 0.66667f
C19856 _0461_ acc0.A\[19\] 0.04646f
C19857 acc0.A\[12\] pp[10] 0
C19858 _0399_ _0088_ 0.03248f
C19859 net46 _1023_/a_561_413# 0
C19860 pp[19] _1023_/a_891_413# 0.00145f
C19861 _0195_ _1028_/a_193_47# 0.04983f
C19862 net56 _0354_ 0.00152f
C19863 hold49/a_391_47# _0202_ 0.02709f
C19864 _1051_/a_891_413# _0148_ 0.00539f
C19865 _0399_ _0407_ 0
C19866 net49 _0762_/a_297_297# 0
C19867 _1057_/a_27_47# _1057_/a_1059_315# 0.04875f
C19868 _1057_/a_193_47# _1057_/a_466_413# 0.07482f
C19869 _0298_ VPWR 0.9324f
C19870 _0414_ _0286_ 0.00168f
C19871 VPWR _0754_/a_240_47# 0.00143f
C19872 _0579_/a_27_297# clknet_1_0__leaf__0459_ 0.03036f
C19873 net21 input19/a_75_212# 0.13399f
C19874 hold81/a_49_47# _0419_ 0
C19875 net225 _1013_/a_27_47# 0
C19876 VPWR _1064_/a_27_47# 0.47884f
C19877 _0966_/a_27_47# clkbuf_1_0__f_clk/a_110_47# 0
C19878 _0443_ clknet_0__0465_ 0.0145f
C19879 _0800_/a_512_297# _0995_/a_27_47# 0
C19880 _0180_ clkbuf_0__0463_/a_110_47# 0.00183f
C19881 net89 _0467_ 0
C19882 _1059_/a_193_47# _1059_/a_466_413# 0.07409f
C19883 _1059_/a_27_47# _1059_/a_1059_315# 0.04875f
C19884 net199 output52/a_27_47# 0
C19885 _0276_ net41 0.01249f
C19886 acc0.A\[14\] _0081_ 0
C19887 _0459_ control0.add 0
C19888 VPWR _0296_ 0.32532f
C19889 _0179_ _0262_ 0
C19890 hold96/a_49_47# _0123_ 0
C19891 _0849_/a_215_47# net222 0.04614f
C19892 clknet_1_0__leaf__0463_ net174 0.02493f
C19893 _1015_/a_27_47# _0345_ 0
C19894 clkbuf_0__0458_/a_110_47# _0431_ 0
C19895 _0517_/a_384_47# net142 0
C19896 clknet_1_0__leaf__0459_ _0398_ 0.06715f
C19897 _1032_/a_891_413# net202 0
C19898 pp[15] net245 0.06915f
C19899 _0288_ net228 0
C19900 net172 net29 0
C19901 _0982_/a_1059_315# net247 0
C19902 _0330_ _0729_/a_68_297# 0.00191f
C19903 _1032_/a_891_413# clknet_1_1__leaf__0463_ 0
C19904 _0569_/a_109_297# _0127_ 0.00169f
C19905 _1065_/a_193_47# clkbuf_1_1__f_clk/a_110_47# 0.00812f
C19906 _0481_ _0978_/a_27_297# 0.1383f
C19907 _0179_ _1058_/a_466_413# 0
C19908 comp0.B\[13\] _0540_/a_51_297# 0.01315f
C19909 hold46/a_285_47# _0540_/a_240_47# 0
C19910 acc0.A\[14\] _0505_/a_373_47# 0.00197f
C19911 _0386_ _0773_/a_285_297# 0.00786f
C19912 _0388_ _0773_/a_117_297# 0.01205f
C19913 _0244_ _0773_/a_285_47# 0.00284f
C19914 _0180_ net131 0
C19915 net45 _0308_ 0
C19916 _0783_/a_79_21# _0398_ 0.07091f
C19917 _0232_ _0352_ 0.04564f
C19918 net44 hold16/a_285_47# 0
C19919 hold46/a_49_47# _0138_ 0
C19920 _0337_ _0705_/a_59_75# 0.16842f
C19921 _0172_ net196 0.06442f
C19922 hold86/a_49_47# _0846_/a_149_47# 0
C19923 _0551_/a_27_47# net8 0
C19924 _0343_ _1055_/a_381_47# 0
C19925 acc0.A\[27\] _1028_/a_891_413# 0
C19926 net189 _0281_ 0
C19927 hold11/a_391_47# _1046_/a_27_47# 0
C19928 _0293_ _0814_/a_109_47# 0
C19929 clknet_0__0461_ hold72/a_49_47# 0.0228f
C19930 hold17/a_285_47# _0488_ 0
C19931 hold17/a_49_47# _0466_ 0.00975f
C19932 net54 _0322_ 0
C19933 acc0.A\[20\] _0603_/a_150_297# 0.00104f
C19934 _1034_/a_891_413# net24 0
C19935 B[7] clkbuf_1_0__f__0463_/a_110_47# 0
C19936 _0949_/a_59_75# _0949_/a_145_75# 0.00658f
C19937 _1052_/a_193_47# _0186_ 0.00351f
C19938 net54 _0327_ 0
C19939 net111 net113 0
C19940 _0376_ acc0.A\[23\] 0
C19941 _0352_ _1006_/a_561_413# 0
C19942 _0570_/a_109_297# net113 0.04463f
C19943 _0570_/a_373_47# clknet_1_1__leaf__0462_ 0
C19944 VPWR _0995_/a_1017_47# 0
C19945 net186 _1033_/a_193_47# 0
C19946 _0284_ _0993_/a_561_413# 0
C19947 clknet_1_0__leaf__0458_ _0268_ 0.00939f
C19948 _0386_ _0350_ 0
C19949 net168 _0179_ 0.47302f
C19950 net61 net248 0.3671f
C19951 net165 _0465_ 0.02112f
C19952 hold101/a_391_47# acc0.A\[4\] 0
C19953 _0225_ net241 0.0655f
C19954 net247 _0451_ 0
C19955 _0731_/a_299_297# _0370_ 0.04564f
C19956 clkbuf_1_0__f__0464_/a_110_47# _1048_/a_193_47# 0
C19957 _0612_/a_59_75# _0612_/a_145_75# 0.00658f
C19958 _0217_ _0585_/a_27_297# 0.0684f
C19959 _0156_ _0187_ 0.06668f
C19960 clknet_1_1__leaf__0460_ net94 0.1426f
C19961 _0663_/a_207_413# _0425_ 0
C19962 net238 net6 0
C19963 _1014_/a_193_47# clkbuf_0__0457_/a_110_47# 0.00277f
C19964 pp[15] net45 0.01805f
C19965 _1056_/a_1059_315# _0515_/a_81_21# 0.00342f
C19966 _0550_/a_240_47# _0137_ 0
C19967 _0259_ _0275_ 0.8578f
C19968 net216 net92 0
C19969 _0533_/a_109_47# _0182_ 0.00355f
C19970 _0533_/a_109_297# _0180_ 0.03117f
C19971 _0533_/a_27_297# net8 0.19803f
C19972 _0951_/a_209_311# _1062_/a_466_413# 0
C19973 hold43/a_391_47# net190 0.13564f
C19974 output55/a_27_47# hold95/a_49_47# 0.00616f
C19975 control0.state\[1\] clknet_1_0__leaf_clk 0.00466f
C19976 _1016_/a_27_47# _0781_/a_68_297# 0
C19977 net106 net202 0.25016f
C19978 _0651_/a_113_47# _0091_ 0
C19979 _0182_ hold71/a_285_47# 0.00378f
C19980 acc0.A\[1\] hold71/a_391_47# 0.03843f
C19981 _0183_ _1060_/a_466_413# 0.0063f
C19982 clknet_0__0464_ net22 0
C19983 hold33/a_391_47# _0174_ 0
C19984 hold71/a_49_47# net218 0.00119f
C19985 hold32/a_49_47# net179 0
C19986 hold32/a_285_47# net141 0
C19987 comp0.B\[7\] comp0.B\[8\] 0.10988f
C19988 net106 clknet_1_1__leaf__0463_ 0
C19989 net140 net13 0
C19990 clknet_1_1__leaf__0459_ _0511_/a_299_297# 0
C19991 pp[9] pp[1] 0
C19992 _0511_/a_384_47# acc0.A\[11\] 0
C19993 hold53/a_49_47# _1024_/a_1059_315# 0
C19994 _0186_ net12 0.31261f
C19995 pp[8] hold34/a_285_47# 0.0637f
C19996 B[13] _0176_ 0
C19997 _0234_ hold94/a_285_47# 0.00856f
C19998 hold88/a_285_47# _0369_ 0
C19999 _0966_/a_27_47# control0.count\[2\] 0
C20000 _0334_ hold62/a_285_47# 0
C20001 _0546_/a_240_47# _0205_ 0
C20002 _1047_/a_193_47# clknet_1_1__leaf__0457_ 0.0049f
C20003 _1047_/a_381_47# clkbuf_1_1__f__0457_/a_110_47# 0.00109f
C20004 VPWR _1023_/a_975_413# 0.00464f
C20005 A[15] _0206_ 0.0017f
C20006 _0984_/a_27_47# _0849_/a_79_21# 0
C20007 _0446_ _0447_ 0.4996f
C20008 _0209_ _1040_/a_193_47# 0
C20009 _0607_/a_27_297# _0387_ 0
C20010 acc0.A\[27\] _0739_/a_79_21# 0.00118f
C20011 clknet_1_0__leaf__0464_ acc0.A\[15\] 0.01743f
C20012 control0.state\[0\] _0880_/a_27_47# 0
C20013 _0991_/a_466_413# _0991_/a_592_47# 0.00553f
C20014 _0991_/a_634_159# _0991_/a_1017_47# 0
C20015 net160 _0213_ 0.00322f
C20016 net36 VPWR 2.22315f
C20017 _0726_/a_240_47# _0219_ 0.07226f
C20018 _0354_ _0345_ 0.18619f
C20019 hold79/a_285_47# _0480_ 0
C20020 _0536_/a_51_297# net134 0
C20021 _0369_ _0487_ 0.07437f
C20022 comp0.B\[14\] _0138_ 0
C20023 _0195_ _0727_/a_277_47# 0
C20024 net39 _0218_ 0.50986f
C20025 net78 hold70/a_49_47# 0
C20026 hold58/a_285_47# net25 0
C20027 _0794_/a_27_47# _0300_ 0.02739f
C20028 _0794_/a_110_297# _0277_ 0
C20029 clknet_1_0__leaf__0463_ clknet_0__0464_ 0
C20030 _0997_/a_193_47# clknet_1_1__leaf__0461_ 0
C20031 net118 control0.reset 0
C20032 clknet_1_1__leaf__0465_ _0345_ 0.0611f
C20033 _0814_/a_27_47# clknet_1_1__leaf__0465_ 0.00274f
C20034 _0216_ _1029_/a_891_413# 0.0042f
C20035 _0328_ acc0.A\[26\] 0.0043f
C20036 _0799_/a_209_47# net5 0.00297f
C20037 clknet_1_0__leaf__0457_ hold73/a_49_47# 0.00995f
C20038 _0982_/a_27_47# acc0.A\[0\] 0.03659f
C20039 _0793_/a_512_297# _0219_ 0.00109f
C20040 _0982_/a_1059_315# net100 0
C20041 _1004_/a_466_413# acc0.A\[23\] 0
C20042 VPWR _1065_/a_193_47# 0.28442f
C20043 _0086_ _0369_ 0.02683f
C20044 _0363_ clkbuf_0__0462_/a_110_47# 0
C20045 hold64/a_49_47# net223 0
C20046 _0159_ _1046_/a_634_159# 0
C20047 clknet_0__0465_ _0089_ 0
C20048 _1001_/a_975_413# _0183_ 0
C20049 _1001_/a_1017_47# _0217_ 0
C20050 comp0.B\[10\] _0542_/a_51_297# 0
C20051 clknet_1_0__leaf__0463_ _1037_/a_381_47# 0.00166f
C20052 net123 _1037_/a_1059_315# 0
C20053 VPWR _0811_/a_81_21# 0.20233f
C20054 comp0.B\[9\] _0540_/a_51_297# 0
C20055 _0399_ _0996_/a_592_47# 0.00151f
C20056 _0725_/a_80_21# acc0.A\[29\] 0.01916f
C20057 _0995_/a_27_47# _0995_/a_193_47# 0.97383f
C20058 _0800_/a_240_47# _0300_ 0
C20059 _0357_ _0701_/a_80_21# 0.06546f
C20060 _0739_/a_215_47# _0321_ 0
C20061 _0229_ _0383_ 0.72436f
C20062 _0739_/a_79_21# _0364_ 0.06893f
C20063 _0417_ _0281_ 0.01923f
C20064 _0226_ _0369_ 0.2043f
C20065 net26 control0.sh 0.20468f
C20066 _1021_/a_891_413# _0183_ 0.0222f
C20067 clkbuf_1_0__f__0458_/a_110_47# acc0.A\[14\] 0
C20068 _0352_ _0321_ 0
C20069 _1060_/a_466_413# acc0.A\[15\] 0.00403f
C20070 _0454_ _0347_ 0.33084f
C20071 hold11/a_285_47# comp0.B\[9\] 0.00201f
C20072 _0315_ net51 0
C20073 _1058_/a_592_47# acc0.A\[10\] 0
C20074 VPWR output52/a_27_47# 0.31007f
C20075 _0828_/a_113_297# _0434_ 0
C20076 _0367_ _0105_ 0.03481f
C20077 comp0.B\[10\] _0142_ 0.00152f
C20078 _0218_ _0444_ 0.03975f
C20079 _0546_/a_51_297# _1042_/a_891_413# 0
C20080 _0546_/a_240_47# _1042_/a_193_47# 0
C20081 net53 _1007_/a_634_159# 0.00282f
C20082 _1070_/a_1059_315# _1069_/a_27_47# 0.00143f
C20083 _1070_/a_27_47# _1069_/a_1059_315# 0.00143f
C20084 _0661_/a_277_297# _0346_ 0
C20085 _0351_ _0352_ 0.24812f
C20086 hold64/a_285_47# _0982_/a_1059_315# 0
C20087 control0.state\[0\] _1062_/a_27_47# 0.00436f
C20088 _0733_/a_222_93# _0328_ 0.01182f
C20089 acc0.A\[29\] _0128_ 0
C20090 hold74/a_49_47# net221 0
C20091 _0343_ clknet_1_1__leaf__0462_ 0
C20092 _0225_ net177 0
C20093 net76 _0986_/a_1059_315# 0
C20094 _0508_/a_299_297# net229 0.07368f
C20095 _0180_ _0529_/a_109_297# 0.03971f
C20096 _1011_/a_27_47# _1011_/a_1059_315# 0.04875f
C20097 _1011_/a_193_47# _1011_/a_466_413# 0.07855f
C20098 _1016_/a_193_47# _0369_ 0.02278f
C20099 _0179_ clknet_1_0__leaf__0464_ 0.23996f
C20100 pp[27] hold62/a_49_47# 0.00512f
C20101 _1034_/a_193_47# net23 0
C20102 VPWR net33 0.50773f
C20103 pp[9] hold34/a_49_47# 0.03158f
C20104 _1004_/a_592_47# net52 0
C20105 VPWR _1031_/a_1017_47# 0
C20106 _0350_ _1006_/a_466_413# 0.02944f
C20107 net150 net51 0
C20108 _0255_ acc0.A\[6\] 0.00276f
C20109 clknet_0__0465_ _0986_/a_891_413# 0.00518f
C20110 _0195_ _1019_/a_975_413# 0
C20111 _0714_/a_149_47# _0195_ 0.00335f
C20112 _0269_ clkbuf_0__0458_/a_110_47# 0.03923f
C20113 VPWR hold51/a_49_47# 0.28329f
C20114 _0296_ _0283_ 0.01009f
C20115 acc0.A\[10\] _0186_ 0.82243f
C20116 hold55/a_49_47# _1067_/a_891_413# 0
C20117 _0752_/a_27_413# hold4/a_285_47# 0
C20118 _1021_/a_27_47# hold73/a_285_47# 0
C20119 _1021_/a_193_47# hold73/a_49_47# 0
C20120 _0461_ net1 0.04233f
C20121 pp[17] _0221_ 0
C20122 _0274_ _0186_ 0.02607f
C20123 net215 net50 0.02783f
C20124 _1020_/a_1059_315# VPWR 0.46103f
C20125 _0350_ _0986_/a_466_413# 0.00151f
C20126 hold33/a_49_47# _0200_ 0.00128f
C20127 hold74/a_391_47# _0459_ 0.00387f
C20128 _0452_ _0345_ 0.04051f
C20129 hold12/a_391_47# VPWR 0.18314f
C20130 hold41/a_285_47# pp[9] 0.00291f
C20131 net189 A[12] 0
C20132 clk _0975_/a_145_75# 0
C20133 _0955_/a_32_297# comp0.B\[6\] 0.13347f
C20134 net162 _0336_ 0.01413f
C20135 _0955_/a_114_297# comp0.B\[5\] 0.00672f
C20136 _0955_/a_304_297# comp0.B\[3\] 0
C20137 VPWR _0515_/a_81_21# 0.21181f
C20138 _0567_/a_27_297# _0345_ 0.00652f
C20139 net172 _0137_ 0
C20140 _0404_ _0794_/a_27_47# 0.09904f
C20141 _0789_/a_75_199# _0277_ 0.06359f
C20142 _0789_/a_201_297# _0300_ 0.00793f
C20143 _0789_/a_208_47# _0297_ 0.00377f
C20144 _1004_/a_1017_47# clknet_1_0__leaf__0460_ 0
C20145 _0305_ _0748_/a_299_297# 0.05782f
C20146 _0680_/a_217_297# _0294_ 0.0248f
C20147 _0523_/a_299_297# _0193_ 0.00863f
C20148 _0524_/a_27_297# _0987_/a_27_47# 0.0238f
C20149 clknet_0__0457_ clkbuf_0__0457_/a_110_47# 1.703f
C20150 clknet_1_1__leaf__0459_ _0799_/a_209_297# 0.00143f
C20151 _0195_ _0116_ 0.04346f
C20152 _1025_/a_592_47# acc0.A\[25\] 0.00256f
C20153 hold33/a_49_47# comp0.B\[8\] 0.3055f
C20154 net65 _0828_/a_199_47# 0
C20155 acc0.A\[7\] _0828_/a_113_297# 0
C20156 net55 _1010_/a_466_413# 0
C20157 _0828_/a_113_297# _0989_/a_1059_315# 0
C20158 _1020_/a_381_47# _1015_/a_193_47# 0
C20159 _1020_/a_193_47# _1015_/a_381_47# 0
C20160 _0181_ clknet_1_0__leaf__0457_ 0.14993f
C20161 _0179_ _1060_/a_466_413# 0
C20162 _0583_/a_27_297# net221 0
C20163 net54 _1008_/a_561_413# 0
C20164 _0486_ _0974_/a_448_47# 0.0581f
C20165 _0217_ _0218_ 0.02463f
C20166 output44/a_27_47# hold61/a_49_47# 0.00616f
C20167 _0271_ _0825_/a_68_297# 0
C20168 control0.add _0772_/a_79_21# 0.01534f
C20169 hold45/a_49_47# clknet_1_1__leaf__0465_ 0
C20170 _0516_/a_27_297# _0516_/a_109_297# 0.17136f
C20171 _1037_/a_27_47# _0552_/a_68_297# 0.00127f
C20172 clknet_0__0457_ _1019_/a_561_413# 0.00129f
C20173 _1010_/a_634_159# _0347_ 0.00831f
C20174 acc0.A\[30\] _0347_ 0
C20175 hold28/a_49_47# acc0.A\[15\] 0
C20176 _0236_ net92 0
C20177 _1051_/a_634_159# clknet_1_1__leaf__0464_ 0
C20178 hold63/a_49_47# _0195_ 0
C20179 hold63/a_285_47# net210 0.01066f
C20180 _0800_/a_149_47# _0298_ 0
C20181 _0190_ _0088_ 0
C20182 net55 _1009_/a_1059_315# 0.08595f
C20183 _0800_/a_51_297# _0345_ 0.11794f
C20184 _0368_ hold90/a_285_47# 0
C20185 _1045_/a_1059_315# clknet_1_1__leaf__0464_ 0.00886f
C20186 _1036_/a_634_159# _1036_/a_381_47# 0
C20187 clknet_1_1__leaf__0459_ _0810_/a_113_47# 0
C20188 _0290_ _0986_/a_193_47# 0
C20189 _0401_ _0986_/a_27_47# 0
C20190 _0346_ _0990_/a_466_413# 0
C20191 _0244_ _0386_ 0.68771f
C20192 hold97/a_285_47# hold9/a_49_47# 0
C20193 control0.sh hold84/a_285_47# 0.00317f
C20194 _0517_/a_299_297# _0988_/a_193_47# 0
C20195 net104 _0346_ 0
C20196 _1072_/a_27_47# _0487_ 0
C20197 _1049_/a_381_47# net154 0
C20198 _1020_/a_1059_315# net48 0
C20199 _0523_/a_81_21# _0150_ 0.11556f
C20200 _0725_/a_209_297# _0725_/a_303_47# 0
C20201 _0111_ _0342_ 0.00332f
C20202 net120 _0457_ 0
C20203 _0433_ _0434_ 0.00126f
C20204 pp[28] _0723_/a_297_47# 0.00121f
C20205 clknet_1_0__leaf__0463_ _0553_/a_149_47# 0
C20206 _0343_ _0429_ 0.21132f
C20207 _1041_/a_27_47# net18 0
C20208 _0458_ _1048_/a_27_47# 0
C20209 _1041_/a_193_47# net198 0
C20210 input14/a_75_212# net13 0
C20211 _0796_/a_215_47# acc0.A\[15\] 0.00176f
C20212 _0238_ _0247_ 0
C20213 _0389_ clknet_1_0__leaf__0460_ 0.00226f
C20214 _1065_/a_1059_315# _0215_ 0
C20215 _0654_/a_207_413# _0419_ 0.01112f
C20216 _0178_ _1048_/a_592_47# 0
C20217 output36/a_27_47# net29 0
C20218 _0467_ clkbuf_0_clk/a_110_47# 0.04162f
C20219 _0529_/a_27_297# net10 0.18568f
C20220 hold33/a_391_47# comp0.B\[13\] 0
C20221 _1041_/a_891_413# hold6/a_49_47# 0
C20222 _1041_/a_466_413# hold6/a_391_47# 0
C20223 net172 comp0.B\[6\] 0
C20224 hold69/a_285_47# _0312_ 0.01652f
C20225 _0965_/a_47_47# net167 0
C20226 control0.count\[3\] _0981_/a_109_297# 0
C20227 _0172_ _0193_ 0
C20228 _0996_/a_466_413# _0219_ 0
C20229 VPWR _0308_ 1.19663f
C20230 _0163_ _1062_/a_193_47# 0.00121f
C20231 _0992_/a_27_47# _0282_ 0
C20232 clknet_1_0__leaf__0462_ _1024_/a_634_159# 0.00275f
C20233 _0467_ _1063_/a_634_159# 0.00857f
C20234 _1058_/a_193_47# net4 0.45349f
C20235 _0742_/a_81_21# net51 0
C20236 B[12] B[11] 0.17109f
C20237 _1021_/a_193_47# _0181_ 0.03451f
C20238 _0399_ _0516_/a_109_297# 0
C20239 net36 _1038_/a_592_47# 0.00276f
C20240 pp[0] _1038_/a_561_413# 0
C20241 _1049_/a_381_47# _0465_ 0
C20242 _0329_ _0355_ 0
C20243 net194 net20 0
C20244 clkload0/a_27_47# clkbuf_1_0__f_clk/a_110_47# 0.00295f
C20245 _0624_/a_59_75# _0255_ 0
C20246 net224 hold77/a_285_47# 0.01139f
C20247 _1012_/a_27_47# net239 0
C20248 _1012_/a_891_413# _0720_/a_68_297# 0.00492f
C20249 _0428_ _0990_/a_1059_315# 0.08224f
C20250 net61 _0447_ 0.21036f
C20251 hold86/a_391_47# _0448_ 0.01657f
C20252 net149 clkbuf_1_1__f__0457_/a_110_47# 0.07473f
C20253 _0585_/a_109_297# clknet_1_1__leaf__0457_ 0
C20254 net111 hold8/a_285_47# 0
C20255 net97 acc0.A\[28\] 0.00151f
C20256 _1054_/a_193_47# _0989_/a_27_47# 0
C20257 _1054_/a_27_47# _0989_/a_193_47# 0
C20258 _0736_/a_56_297# _0107_ 0.00416f
C20259 _0570_/a_27_297# hold8/a_391_47# 0
C20260 _0570_/a_109_297# hold8/a_285_47# 0
C20261 _1057_/a_891_413# _1057_/a_1017_47# 0.00617f
C20262 _1057_/a_193_47# net189 0.51577f
C20263 clkbuf_0__0463_/a_110_47# _0498_/a_51_297# 0
C20264 _0269_ _0986_/a_975_413# 0
C20265 pp[17] _0344_ 0
C20266 _0195_ _0534_/a_384_47# 0
C20267 _0111_ _1013_/a_592_47# 0.00188f
C20268 net1 _0465_ 0
C20269 _0209_ _0207_ 0.42936f
C20270 _0607_/a_373_47# clknet_0__0461_ 0
C20271 _0579_/a_27_297# _0579_/a_373_47# 0.01338f
C20272 _0179_ hold28/a_49_47# 0.05656f
C20273 clknet_0__0463_ comp0.B\[10\] 0.01197f
C20274 _0216_ hold62/a_49_47# 0
C20275 _0195_ hold62/a_391_47# 0.04355f
C20276 _0379_ net93 0
C20277 _0730_/a_79_21# clkbuf_1_1__f__0462_/a_110_47# 0
C20278 _0093_ _0995_/a_27_47# 0.20784f
C20279 _1059_/a_193_47# _0157_ 0.26097f
C20280 _1059_/a_891_413# _1059_/a_1017_47# 0.00617f
C20281 _0789_/a_75_199# _0298_ 0.10389f
C20282 _0789_/a_201_297# _0404_ 0.01098f
C20283 _1059_/a_634_159# net145 0
C20284 _1041_/a_1059_315# _1041_/a_1017_47# 0
C20285 _0693_/a_68_297# net52 0.1232f
C20286 _0369_ net41 0
C20287 net231 _1062_/a_1017_47# 0.00137f
C20288 _0528_/a_81_21# _0148_ 0.115f
C20289 _0528_/a_384_47# net170 0.01004f
C20290 net36 _0453_ 0.09184f
C20291 _0568_/a_109_47# _0219_ 0
C20292 _0500_/a_27_47# _0145_ 0.08603f
C20293 pp[15] VPWR 0.47095f
C20294 _0510_/a_109_297# _0186_ 0.05708f
C20295 clknet_1_0__leaf__0465_ clknet_1_1__leaf__0464_ 0.06039f
C20296 _0433_ _0989_/a_1059_315# 0
C20297 _0811_/a_81_21# _0283_ 0.05219f
C20298 _0221_ _0355_ 0.30671f
C20299 _1055_/a_27_47# clknet_1_1__leaf__0465_ 0.04896f
C20300 net248 _0431_ 0
C20301 _0181_ _1047_/a_891_413# 0
C20302 _0710_/a_109_47# _0341_ 0.00138f
C20303 _0710_/a_109_297# _0340_ 0.00905f
C20304 _0779_/a_79_21# _0347_ 0.12066f
C20305 clknet_1_0__leaf_clk _1068_/a_634_159# 0
C20306 _0443_ _0986_/a_27_47# 0.00858f
C20307 _0592_/a_68_297# _0380_ 0
C20308 clknet_1_0__leaf__0458_ net222 0.00138f
C20309 _0352_ _0771_/a_27_413# 0.02055f
C20310 clknet_1_1__leaf__0463_ net122 0.18497f
C20311 net168 hold83/a_49_47# 0.0466f
C20312 _0310_ _0347_ 0.00927f
C20313 clknet_1_1__leaf__0460_ _1007_/a_193_47# 0.00134f
C20314 pp[16] hold98/a_49_47# 0
C20315 _0107_ net224 0
C20316 _0693_/a_150_297# clknet_1_0__leaf__0460_ 0
C20317 _0399_ _0096_ 0.16288f
C20318 _0369_ net217 0.25631f
C20319 _1030_/a_381_47# clknet_1_1__leaf__0462_ 0
C20320 net120 _0475_ 0
C20321 hold32/a_391_47# pp[8] 0.04703f
C20322 _0536_/a_51_297# net22 0.17441f
C20323 VPWR _0686_/a_301_297# 0
C20324 _0850_/a_68_297# _0181_ 0
C20325 _0248_ _0218_ 0
C20326 _0372_ _0294_ 0.11824f
C20327 _0125_ net114 0.04192f
C20328 _0974_/a_79_199# _1068_/a_27_47# 0.00155f
C20329 _1054_/a_1059_315# _0087_ 0.00102f
C20330 VPWR _1008_/a_381_47# 0.07829f
C20331 _0981_/a_27_297# clkbuf_1_0__f_clk/a_110_47# 0
C20332 _0331_ acc0.A\[29\] 0
C20333 net158 _1046_/a_381_47# 0.12138f
C20334 _0180_ net170 0.1181f
C20335 hold11/a_49_47# net132 0
C20336 _0338_ _0723_/a_27_413# 0
C20337 _0335_ _0723_/a_207_413# 0.00721f
C20338 _0891_/a_27_47# _1015_/a_634_159# 0
C20339 _1028_/a_27_47# _1027_/a_1059_315# 0
C20340 _1020_/a_1059_315# clknet_1_0__leaf__0459_ 0.01089f
C20341 output55/a_27_47# _1011_/a_27_47# 0
C20342 _0467_ _1062_/a_381_47# 0
C20343 net21 net18 0.02213f
C20344 net89 net1 0
C20345 _0180_ _0845_/a_109_297# 0
C20346 net5 _0668_/a_79_21# 0
C20347 clknet_1_0__leaf__0458_ _0182_ 0.58024f
C20348 _0798_/a_113_297# _0409_ 0.00101f
C20349 _0341_ _1013_/a_193_47# 0
C20350 _0340_ _1013_/a_27_47# 0
C20351 _0179_ hold47/a_391_47# 0.00232f
C20352 net144 _0513_/a_299_297# 0.00997f
C20353 net168 input13/a_75_212# 0
C20354 clknet_1_0__leaf__0463_ _0536_/a_51_297# 0.00349f
C20355 _0369_ _0744_/a_27_47# 0.35949f
C20356 _0545_/a_68_297# _0545_/a_150_297# 0.00477f
C20357 _0408_ hold91/a_391_47# 0
C20358 _0368_ clknet_0__0462_ 0
C20359 _0369_ _0760_/a_47_47# 0.01046f
C20360 _0217_ _0112_ 0.36038f
C20361 clknet_1_1__leaf__0460_ _0328_ 0.02382f
C20362 _0699_/a_68_297# _0331_ 0.10723f
C20363 _0299_ _0995_/a_193_47# 0.00408f
C20364 _0221_ _0569_/a_27_297# 0
C20365 hold33/a_391_47# comp0.B\[9\] 0.03245f
C20366 _1010_/a_193_47# hold95/a_285_47# 0
C20367 _1010_/a_27_47# hold95/a_391_47# 0
C20368 pp[28] _0356_ 0
C20369 VPWR _0652_/a_109_297# 0.00778f
C20370 _1030_/a_27_47# net239 0
C20371 clknet_1_0__leaf__0462_ _0577_/a_109_297# 0.01333f
C20372 _1031_/a_27_47# _1031_/a_193_47# 0.97099f
C20373 net8 _0199_ 0.13907f
C20374 clkload0/a_27_47# control0.count\[2\] 0.00137f
C20375 net34 clk 0.0577f
C20376 _0951_/a_209_311# _0160_ 0.0255f
C20377 hold69/a_391_47# _0219_ 0
C20378 _0183_ _0158_ 0.12105f
C20379 hold19/a_285_47# _0181_ 0
C20380 _1014_/a_193_47# _0350_ 0
C20381 _0343_ clknet_1_1__leaf__0458_ 0.15287f
C20382 VPWR _0563_/a_149_47# 0
C20383 B[8] _0546_/a_240_47# 0
C20384 _0457_ _1034_/a_466_413# 0
C20385 control0.state\[1\] _1063_/a_381_47# 0.0165f
C20386 hold26/a_285_47# _0545_/a_68_297# 0
C20387 net207 _1014_/a_891_413# 0
C20388 hold44/a_49_47# hold44/a_391_47# 0.00188f
C20389 clknet_1_0__leaf__0462_ _1022_/a_1017_47# 0
C20390 _1005_/a_466_413# _1005_/a_381_47# 0.03733f
C20391 _1005_/a_193_47# _1005_/a_975_413# 0
C20392 _1005_/a_1059_315# _1005_/a_891_413# 0.31086f
C20393 _0731_/a_299_297# _0731_/a_384_47# 0
C20394 _0705_/a_59_75# _0333_ 0
C20395 _0534_/a_81_21# net247 0.03581f
C20396 _0769_/a_81_21# _0616_/a_215_47# 0
C20397 net152 _0139_ 0.04056f
C20398 _0955_/a_32_297# net26 0
C20399 _0984_/a_193_47# _0082_ 0.54237f
C20400 _0984_/a_1059_315# net222 0.00581f
C20401 _1066_/a_193_47# _1062_/a_27_47# 0
C20402 _1066_/a_27_47# _1062_/a_193_47# 0
C20403 _0188_ _0186_ 0.05163f
C20404 clkbuf_1_1__f__0463_/a_110_47# net17 0
C20405 _1060_/a_193_47# _0507_/a_109_297# 0
C20406 _1013_/a_634_159# _1013_/a_1059_315# 0
C20407 _1013_/a_27_47# _1013_/a_381_47# 0.06222f
C20408 _1013_/a_193_47# _1013_/a_891_413# 0.19683f
C20409 clknet_1_0__leaf__0465_ net247 0
C20410 _0125_ _0365_ 0
C20411 _0991_/a_381_47# net67 0
C20412 _0991_/a_592_47# _0089_ 0.00288f
C20413 VPWR _0527_/a_27_297# 0.19128f
C20414 _1002_/a_27_47# _1002_/a_634_159# 0.14145f
C20415 hold46/a_49_47# net22 0
C20416 _1017_/a_27_47# _0583_/a_27_297# 0
C20417 hold26/a_49_47# hold26/a_285_47# 0.22264f
C20418 _0309_ _0775_/a_510_47# 0
C20419 _1027_/a_27_47# _0347_ 0
C20420 _0424_ _0218_ 0
C20421 _0617_/a_150_297# _0219_ 0
C20422 _0367_ _0359_ 0.14577f
C20423 _0315_ _0324_ 0.20238f
C20424 _0766_/a_109_297# _0393_ 0
C20425 _0985_/a_561_413# _0261_ 0
C20426 _0985_/a_975_413# _0262_ 0
C20427 _1017_/a_193_47# net43 0
C20428 _0607_/a_27_297# acc0.A\[16\] 0.09177f
C20429 _0286_ _0419_ 0.02959f
C20430 net165 _1060_/a_634_159# 0
C20431 clknet_1_1__leaf__0459_ _0997_/a_891_413# 0.02439f
C20432 _0467_ net185 0
C20433 output59/a_27_47# _0350_ 0
C20434 clknet_1_1__leaf__0459_ _0992_/a_592_47# 0.00163f
C20435 VPWR _0989_/a_634_159# 0.18372f
C20436 hold32/a_285_47# pp[9] 0.00219f
C20437 _0217_ net240 0
C20438 _0357_ _0330_ 0.19161f
C20439 VPWR hold1/a_391_47# 0.18384f
C20440 _0095_ _0219_ 0.00659f
C20441 hold64/a_391_47# _1019_/a_891_413# 0.00406f
C20442 _0174_ net195 0.14974f
C20443 _0180_ _0525_/a_81_21# 0.01436f
C20444 _1038_/a_891_413# _1040_/a_193_47# 0
C20445 _1038_/a_1059_315# _1040_/a_634_159# 0
C20446 _1012_/a_1059_315# hold92/a_391_47# 0.0103f
C20447 VPWR _0992_/a_634_159# 0.18025f
C20448 _0343_ _0263_ 0
C20449 _0343_ clkload4/Y 0.01605f
C20450 _0217_ _0099_ 0.04494f
C20451 _0768_/a_27_47# _0347_ 0.00301f
C20452 net103 _0790_/a_35_297# 0
C20453 _0995_/a_466_413# _0995_/a_592_47# 0.00553f
C20454 _0995_/a_634_159# _0995_/a_1017_47# 0
C20455 _0765_/a_79_21# _0765_/a_297_297# 0.01735f
C20456 _0680_/a_80_21# _0359_ 0.0107f
C20457 net10 _0196_ 0
C20458 hold46/a_49_47# clknet_1_0__leaf__0463_ 0
C20459 VPWR _1061_/a_27_47# 0.68215f
C20460 _0437_ _0829_/a_109_297# 0
C20461 _0565_/a_512_297# clknet_1_0__leaf__0461_ 0
C20462 _0343_ _0582_/a_373_47# 0
C20463 hold59/a_391_47# acc0.A\[18\] 0
C20464 _0983_/a_891_413# _0346_ 0
C20465 _0158_ acc0.A\[15\] 0.04033f
C20466 _0732_/a_80_21# _0460_ 0
C20467 net82 _0507_/a_27_297# 0.0054f
C20468 _0501_/a_27_47# _0180_ 0.19093f
C20469 _1070_/a_1059_315# _0489_ 0
C20470 _0244_ _0854_/a_79_21# 0
C20471 _1034_/a_27_47# _0173_ 0.0469f
C20472 _1034_/a_193_47# _0213_ 0.01888f
C20473 _1034_/a_891_413# _0561_/a_149_47# 0
C20474 _1034_/a_1059_315# _0561_/a_240_47# 0
C20475 net185 comp0.B\[0\] 0
C20476 _0579_/a_27_297# _0345_ 0
C20477 hold64/a_391_47# net206 0
C20478 _0217_ _0581_/a_109_47# 0.00231f
C20479 _0183_ _0581_/a_27_297# 0.18198f
C20480 net36 net30 0
C20481 net145 _0082_ 0
C20482 VPWR _0428_ 0.82473f
C20483 _0183_ acc0.A\[14\] 0.16541f
C20484 net32 _1042_/a_381_47# 0.01657f
C20485 _0139_ _1042_/a_466_413# 0
C20486 _1018_/a_1059_315# _0459_ 0
C20487 net53 net93 0
C20488 _0369_ net66 0.61168f
C20489 hold86/a_49_47# acc0.A\[15\] 0.00454f
C20490 net56 _0353_ 0.00789f
C20491 acc0.A\[21\] net213 0
C20492 _0168_ _1069_/a_193_47# 0
C20493 _1070_/a_634_159# clknet_1_0__leaf_clk 0
C20494 _0975_/a_59_75# _0970_/a_27_297# 0.00484f
C20495 VPWR _1069_/a_466_413# 0.25726f
C20496 control0.state\[1\] _1062_/a_1017_47# 0
C20497 VPWR hold60/a_391_47# 0.16799f
C20498 hold27/a_391_47# net173 0
C20499 _1034_/a_466_413# _0475_ 0
C20500 _0398_ _0345_ 0
C20501 _1056_/a_27_47# _1058_/a_27_47# 0
C20502 clkbuf_1_0__f__0460_/a_110_47# _0460_ 0.02624f
C20503 _1011_/a_634_159# net97 0
C20504 _1011_/a_891_413# _1011_/a_1017_47# 0.00617f
C20505 _0274_ net62 0.09761f
C20506 _0985_/a_634_159# _0186_ 0.00549f
C20507 _0239_ _0347_ 0.03762f
C20508 _1000_/a_193_47# _0614_/a_29_53# 0
C20509 _0399_ _0304_ 0
C20510 _0644_/a_47_47# hold91/a_285_47# 0
C20511 clkbuf_0__0462_/a_110_47# _0686_/a_219_297# 0.01043f
C20512 input34/a_27_47# _0162_ 0
C20513 _0182_ _0532_/a_299_297# 0.06414f
C20514 _0180_ _0532_/a_81_21# 0
C20515 _1006_/a_27_47# _1006_/a_891_413# 0.03206f
C20516 _1006_/a_193_47# _1006_/a_1059_315# 0.03405f
C20517 _1006_/a_634_159# _1006_/a_466_413# 0.23992f
C20518 output37/a_27_47# _0187_ 0
C20519 _0538_/a_512_297# VPWR 0.00729f
C20520 clkload2/Y _0196_ 0.00103f
C20521 _0532_/a_81_21# net218 0.06277f
C20522 _0993_/a_27_47# _0807_/a_68_297# 0
C20523 net45 _0997_/a_592_47# 0
C20524 _0250_ _0460_ 0.07072f
C20525 _0972_/a_584_47# _0487_ 0.00205f
C20526 comp0.B\[14\] net22 0
C20527 pp[8] _0153_ 0.006f
C20528 _0316_ hold97/a_391_47# 0.00577f
C20529 _0984_/a_27_47# _0984_/a_634_159# 0.14145f
C20530 _0347_ _1026_/a_466_413# 0
C20531 clknet_1_0__leaf__0462_ _0756_/a_129_47# 0
C20532 _0212_ _1034_/a_193_47# 0
C20533 _0808_/a_81_21# _0808_/a_266_47# 0.04342f
C20534 _1055_/a_975_413# VPWR 0.00733f
C20535 net182 _0515_/a_81_21# 0
C20536 _0243_ _0346_ 0
C20537 _0102_ _1024_/a_466_413# 0
C20538 _0352_ _1024_/a_1059_315# 0
C20539 _1003_/a_561_413# VPWR 0.00309f
C20540 _0251_ _0435_ 0.00993f
C20541 hold65/a_49_47# _0253_ 0.00514f
C20542 _0982_/a_193_47# _0117_ 0
C20543 _0457_ net118 0.01086f
C20544 hold77/a_285_47# hold77/a_391_47# 0.41909f
C20545 clknet_0__0464_ _1049_/a_381_47# 0
C20546 _0955_/a_32_297# hold84/a_285_47# 0
C20547 net35 _1068_/a_891_413# 0.00681f
C20548 _1039_/a_27_47# VPWR 0.42411f
C20549 _0343_ clknet_1_0__leaf__0461_ 0
C20550 comp0.B\[6\] _0474_ 0.30826f
C20551 pp[9] net4 0
C20552 _0712_/a_79_21# _1031_/a_193_47# 0
C20553 _0986_/a_27_47# _0986_/a_891_413# 0.03224f
C20554 _0986_/a_193_47# _0986_/a_1059_315# 0.03405f
C20555 _0986_/a_634_159# _0986_/a_466_413# 0.23992f
C20556 net148 _0987_/a_891_413# 0
C20557 _0194_ _0987_/a_27_47# 0
C20558 _0277_ _0345_ 0.19244f
C20559 net49 net151 0
C20560 _0715_/a_27_47# VPWR 0.38483f
C20561 _1017_/a_634_159# _0181_ 0.01776f
C20562 _1023_/a_634_159# _1023_/a_381_47# 0
C20563 _0616_/a_78_199# _1006_/a_27_47# 0
C20564 clkbuf_1_0__f__0461_/a_110_47# _0247_ 0.0344f
C20565 _0240_ _0350_ 0
C20566 net224 _0322_ 0
C20567 _0179_ _0158_ 0.07112f
C20568 _0344_ _0567_/a_109_297# 0.03138f
C20569 _0627_/a_215_53# _0271_ 0
C20570 _0297_ _0669_/a_29_53# 0
C20571 output36/a_27_47# comp0.B\[6\] 0
C20572 _0747_/a_79_21# acc0.A\[24\] 0
C20573 _1042_/a_466_413# _1042_/a_561_413# 0.00772f
C20574 _1042_/a_634_159# _1042_/a_975_413# 0
C20575 _0369_ _0350_ 0.39878f
C20576 hold59/a_49_47# hold59/a_391_47# 0.00188f
C20577 _0156_ clknet_1_1__leaf__0465_ 0.02636f
C20578 acc0.A\[14\] acc0.A\[15\] 0.59561f
C20579 _1019_/a_27_47# control0.add 0
C20580 clknet_1_0__leaf__0458_ _0089_ 0
C20581 _0181_ _1060_/a_1017_47# 0.00114f
C20582 _0114_ net221 0
C20583 net165 _0115_ 0
C20584 clknet_0__0457_ _0350_ 0
C20585 net224 _0327_ 0
C20586 input12/a_75_212# net12 0.10944f
C20587 net22 _0543_/a_68_297# 0
C20588 _1003_/a_27_47# clknet_0_clk 0
C20589 _0516_/a_109_297# _0190_ 0.00176f
C20590 _0516_/a_373_47# net16 0.00188f
C20591 _1037_/a_1059_315# _0209_ 0.00178f
C20592 _1010_/a_1017_47# _0352_ 0
C20593 net96 _0347_ 0.00455f
C20594 _0401_ _0288_ 0.06735f
C20595 output42/a_27_47# _0297_ 0
C20596 output50/a_27_47# pp[24] 0
C20597 clknet_1_1__leaf__0464_ _1044_/a_466_413# 0.01332f
C20598 _1045_/a_27_47# net20 0.00571f
C20599 hold86/a_49_47# _0179_ 0
C20600 clknet_1_1__leaf__0460_ _0108_ 0.23754f
C20601 net137 clknet_1_1__leaf__0464_ 0.2185f
C20602 _0179_ _1050_/a_561_413# 0
C20603 _0093_ _0299_ 0
C20604 _0699_/a_68_297# _1008_/a_27_47# 0
C20605 comp0.B\[3\] _1065_/a_193_47# 0.00133f
C20606 net58 _0435_ 0
C20607 net243 _0757_/a_68_297# 0.10105f
C20608 _0625_/a_59_75# _0442_ 0
C20609 _1036_/a_634_159# comp0.B\[4\] 0
C20610 _1036_/a_891_413# net161 0
C20611 _0447_ _0431_ 0
C20612 clknet_0__0460_ hold90/a_285_47# 0
C20613 _0346_ _0088_ 0
C20614 _0466_ _1064_/a_634_159# 0
C20615 pp[30] net209 0.0301f
C20616 net10 _1042_/a_381_47# 0.01201f
C20617 _0346_ _0407_ 0
C20618 net120 _1033_/a_193_47# 0
C20619 _0305_ _0508_/a_81_21# 0
C20620 hold18/a_285_47# acc0.A\[1\] 0
C20621 hold18/a_49_47# _0182_ 0
C20622 _0598_/a_297_47# net213 0
C20623 _0230_ hold66/a_285_47# 0
C20624 _0742_/a_299_297# _0359_ 0
C20625 _0742_/a_81_21# _0324_ 0
C20626 _0226_ hold66/a_391_47# 0
C20627 _0153_ _0988_/a_891_413# 0
C20628 _0984_/a_193_47# net145 0
C20629 _0107_ hold77/a_391_47# 0
C20630 net31 _0176_ 0.02466f
C20631 _0404_ net79 0
C20632 _1059_/a_27_47# _0506_/a_81_21# 0
C20633 _0808_/a_81_21# _0345_ 0.14179f
C20634 _0316_ _0315_ 0
C20635 _0621_/a_35_297# _0369_ 0.00145f
C20636 pp[29] _1011_/a_193_47# 0
C20637 _0387_ _0679_/a_68_297# 0
C20638 VPWR _1040_/a_975_413# 0.00468f
C20639 _0992_/a_891_413# clknet_1_1__leaf__0465_ 0
C20640 clknet_1_0__leaf__0460_ net50 0.00427f
C20641 clknet_0__0463_ _0177_ 0
C20642 net240 _0971_/a_81_21# 0
C20643 _0315_ _0347_ 0
C20644 control0.reset _0175_ 0.02997f
C20645 _1036_/a_891_413# net26 0.00309f
C20646 _0743_/a_51_297# _0743_/a_149_47# 0.02487f
C20647 _0998_/a_27_47# _0459_ 0
C20648 clknet_1_0__leaf__0458_ _0986_/a_891_413# 0
C20649 _1002_/a_27_47# net220 0
C20650 _1054_/a_193_47# net11 0.03128f
C20651 clknet_1_0__leaf__0462_ net110 0.11724f
C20652 _0391_ hold40/a_285_47# 0
C20653 net223 hold40/a_391_47# 0
C20654 _0313_ acc0.A\[27\] 0
C20655 hold34/a_285_47# A[10] 0.03571f
C20656 _0178_ clknet_1_1__leaf__0457_ 0.08938f
C20657 _0571_/a_27_297# _0571_/a_373_47# 0.01338f
C20658 _0662_/a_299_297# _0292_ 0
C20659 _0353_ _0345_ 0
C20660 acc0.A\[3\] _0465_ 0
C20661 _0743_/a_51_297# _0345_ 0.11536f
C20662 _0999_/a_1059_315# _0218_ 0.08636f
C20663 net125 net201 0
C20664 _0856_/a_215_47# acc0.A\[1\] 0.0487f
C20665 net33 comp0.B\[3\] 0
C20666 _0409_ net41 0.00502f
C20667 _0606_/a_215_297# _0372_ 0
C20668 _0179_ acc0.A\[14\] 0
C20669 _0305_ _0246_ 0.00345f
C20670 _0311_ _0245_ 0
C20671 control0.sh _0465_ 0.0016f
C20672 clknet_1_0__leaf__0464_ _1049_/a_891_413# 0
C20673 acc0.A\[2\] acc0.A\[3\] 0.02455f
C20674 net133 _1049_/a_466_413# 0
C20675 _0258_ VPWR 0.80638f
C20676 hold41/a_391_47# A[10] 0
C20677 _0179_ clkbuf_1_0__f__0464_/a_110_47# 0.04362f
C20678 _1058_/a_1059_315# acc0.A\[11\] 0
C20679 _0217_ hold3/a_285_47# 0
C20680 net150 hold3/a_391_47# 0.13645f
C20681 _0279_ _0403_ 0.56696f
C20682 _1000_/a_27_47# net223 0
C20683 VPWR _1035_/a_466_413# 0.25821f
C20684 _1053_/a_1059_315# _1052_/a_891_413# 0
C20685 _1001_/a_193_47# net45 0
C20686 _0298_ _0345_ 0
C20687 _0225_ hold4/a_49_47# 0.00251f
C20688 _0754_/a_512_297# _0377_ 0
C20689 _0754_/a_51_297# _0219_ 0.13909f
C20690 _0754_/a_240_47# _0345_ 0.00634f
C20691 _0272_ _0270_ 0
C20692 _0982_/a_634_159# _0181_ 0.04108f
C20693 _0179_ _1053_/a_634_159# 0
C20694 _0549_/a_68_297# net29 0.00733f
C20695 _0992_/a_634_159# _0283_ 0
C20696 _0992_/a_193_47# _0286_ 0
C20697 _0844_/a_79_21# _0350_ 0
C20698 _1056_/a_891_413# output66/a_27_47# 0
C20699 _1056_/a_27_47# pp[8] 0
C20700 acc0.A\[21\] hold73/a_391_47# 0.00106f
C20701 _0313_ _0364_ 0.15713f
C20702 _0458_ _0643_/a_253_47# 0
C20703 _1064_/a_27_47# _1064_/a_466_413# 0.26005f
C20704 _1064_/a_193_47# _1064_/a_634_159# 0.12729f
C20705 _0296_ _0345_ 0.04868f
C20706 net158 clknet_1_0__leaf__0465_ 0.01076f
C20707 _0837_/a_81_21# _0271_ 0
C20708 net224 _0306_ 0
C20709 _0396_ _0352_ 0.31943f
C20710 clknet_1_1__leaf__0459_ _0786_/a_217_297# 0.00151f
C20711 clk _1068_/a_466_413# 0
C20712 _1054_/a_634_159# hold7/a_285_47# 0
C20713 _1018_/a_193_47# _1017_/a_193_47# 0.00131f
C20714 pp[16] clknet_1_1__leaf__0459_ 0
C20715 clkbuf_0_clk/a_110_47# net1 0
C20716 VPWR net113 0.84429f
C20717 _0295_ _0304_ 0.07867f
C20718 _0255_ _0826_/a_219_297# 0.1286f
C20719 hold65/a_49_47# output61/a_27_47# 0
C20720 _1038_/a_891_413# _0207_ 0.00764f
C20721 _0769_/a_299_297# _0771_/a_27_413# 0
C20722 _0769_/a_81_21# _0771_/a_215_297# 0.01092f
C20723 net58 _0456_ 0
C20724 _0712_/a_79_21# _0712_/a_297_297# 0.05317f
C20725 _0587_/a_27_47# hold92/a_391_47# 0
C20726 _1051_/a_634_159# net148 0
C20727 _0455_ net222 0
C20728 _1033_/a_634_159# comp0.B\[0\] 0.01202f
C20729 net132 net20 0
C20730 _0163_ net17 0
C20731 _0348_ _0723_/a_27_413# 0.00126f
C20732 _0568_/a_27_297# clknet_1_1__leaf__0462_ 0.00187f
C20733 VPWR _0994_/a_975_413# 0.00464f
C20734 _0343_ _1060_/a_891_413# 0.002f
C20735 net159 _1068_/a_1059_315# 0
C20736 control0.state\[0\] _0970_/a_114_47# 0.00179f
C20737 control0.state\[1\] _0970_/a_27_297# 0
C20738 _0170_ clkbuf_1_0__f_clk/a_110_47# 0.00203f
C20739 net167 clknet_0_clk 0.03983f
C20740 hold19/a_285_47# clknet_1_1__leaf__0461_ 0
C20741 clknet_1_0__leaf__0458_ _0854_/a_215_47# 0.00121f
C20742 clknet_0__0465_ _0841_/a_297_297# 0
C20743 _1010_/a_381_47# _0350_ 0.01189f
C20744 _0576_/a_109_297# net50 0
C20745 _0477_ _0951_/a_296_53# 0
C20746 net145 net67 0
C20747 hold13/a_391_47# _1034_/a_891_413# 0
C20748 _0259_ _0990_/a_466_413# 0
C20749 _0339_ net209 0.00521f
C20750 net44 net239 0.15171f
C20751 _0565_/a_149_47# _0173_ 0.02555f
C20752 _0565_/a_51_297# _0208_ 0.15218f
C20753 _0305_ net103 0.0346f
C20754 net88 net202 0.00239f
C20755 net157 _0465_ 0.08021f
C20756 net61 _0275_ 0
C20757 hold65/a_285_47# _0518_/a_27_297# 0
C20758 _0479_ clknet_1_0__leaf_clk 0.00178f
C20759 _0989_/a_27_47# acc0.A\[6\] 0
C20760 _0846_/a_240_47# _0350_ 0.00277f
C20761 hold70/a_285_47# net37 0.00333f
C20762 VPWR _0720_/a_150_297# 0.00246f
C20763 hold36/a_285_47# _0538_/a_240_47# 0
C20764 _0383_ _0382_ 0.05257f
C20765 _1056_/a_193_47# _0988_/a_1059_315# 0
C20766 _1056_/a_27_47# _0988_/a_891_413# 0
C20767 _0995_/a_381_47# _0219_ 0
C20768 comp0.B\[4\] comp0.B\[5\] 0.25142f
C20769 clknet_0__0462_ clknet_0__0460_ 0
C20770 _0174_ _0204_ 0.16477f
C20771 _0695_/a_472_297# _0323_ 0.00127f
C20772 _0695_/a_80_21# _0327_ 0.11839f
C20773 net214 _0399_ 0.00436f
C20774 net175 _0261_ 0
C20775 _0180_ _0498_/a_240_47# 0
C20776 _0222_ _0232_ 0.06064f
C20777 input31/a_75_212# B[8] 0.19861f
C20778 _1037_/a_27_47# VPWR 0.71572f
C20779 net247 hold71/a_391_47# 0.04768f
C20780 clkbuf_1_1__f_clk/a_110_47# _0880_/a_27_47# 0.01306f
C20781 comp0.B\[10\] net198 0.21846f
C20782 _0183_ _1016_/a_634_159# 0
C20783 _1031_/a_466_413# _1031_/a_592_47# 0.00553f
C20784 _1031_/a_634_159# _1031_/a_1017_47# 0
C20785 _0289_ _0786_/a_80_21# 0.17233f
C20786 _0080_ clkbuf_1_1__f__0457_/a_110_47# 0
C20787 _1041_/a_466_413# VPWR 0.24364f
C20788 _0416_ _0403_ 0.08928f
C20789 net105 acc0.A\[0\] 0.0032f
C20790 _1022_/a_193_47# _1005_/a_27_47# 0
C20791 pp[15] _0995_/a_634_159# 0.00431f
C20792 _1005_/a_381_47# _0103_ 0.13417f
C20793 _0244_ _0240_ 0.19273f
C20794 _0325_ _0367_ 0
C20795 _0474_ net26 0
C20796 clknet_0__0458_ clknet_0__0465_ 0.17533f
C20797 _0244_ _0369_ 0
C20798 _1060_/a_1059_315# net5 0
C20799 _1060_/a_634_159# _0185_ 0.00167f
C20800 _0366_ _1025_/a_193_47# 0
C20801 _1054_/a_193_47# clknet_1_1__leaf__0458_ 0
C20802 _0857_/a_27_47# clkbuf_1_1__f_clk/a_110_47# 0
C20803 _1002_/a_381_47# _1002_/a_561_413# 0.00123f
C20804 _1002_/a_27_47# net88 0.29632f
C20805 _1002_/a_891_413# _1002_/a_975_413# 0.00851f
C20806 _1014_/a_1059_315# _0264_ 0
C20807 _1027_/a_634_159# _0365_ 0
C20808 _1027_/a_27_47# _0106_ 0
C20809 _1021_/a_1059_315# net1 0.01547f
C20810 clknet_1_0__leaf__0465_ net148 0.07467f
C20811 acc0.A\[20\] VPWR 1.12421f
C20812 net29 _1040_/a_891_413# 0
C20813 _0268_ _0448_ 0
C20814 _0269_ _0447_ 0.00167f
C20815 _0984_/a_592_47# clknet_1_0__leaf__0458_ 0
C20816 _0820_/a_79_21# _0820_/a_215_47# 0.04584f
C20817 net36 _0345_ 0.0238f
C20818 net165 net146 0
C20819 _0466_ clknet_1_0__leaf__0460_ 0
C20820 hold28/a_285_47# _1049_/a_1059_315# 0.0054f
C20821 _0710_/a_109_47# acc0.A\[30\] 0
C20822 _0343_ _0642_/a_27_413# 0.00332f
C20823 clkbuf_1_0__f__0459_/a_110_47# clkload4/Y 0.00214f
C20824 hold64/a_49_47# _0350_ 0.02136f
C20825 _0154_ _1055_/a_891_413# 0
C20826 VPWR _0997_/a_592_47# 0
C20827 _0309_ _0347_ 0.02048f
C20828 _1038_/a_466_413# net174 0
C20829 _0183_ _1019_/a_975_413# 0
C20830 _0799_/a_80_21# _0297_ 0
C20831 net175 _0509_/a_27_47# 0
C20832 _1001_/a_27_47# net46 0.00182f
C20833 net104 net221 0
C20834 pp[26] hold8/a_49_47# 0
C20835 net54 hold8/a_391_47# 0.00529f
C20836 _1041_/a_634_159# _0550_/a_51_297# 0
C20837 _0437_ _0827_/a_27_47# 0
C20838 hold77/a_391_47# _0327_ 0
C20839 _0109_ clknet_1_1__leaf__0462_ 0.00242f
C20840 _0285_ net38 0.05693f
C20841 _0822_/a_109_297# clknet_0__0458_ 0.0017f
C20842 _0170_ control0.count\[2\] 0
C20843 pp[28] _1011_/a_891_413# 0.00103f
C20844 net69 _0853_/a_68_297# 0.02065f
C20845 _0089_ _0288_ 0
C20846 net36 hold2/a_49_47# 0
C20847 net230 net138 0.00199f
C20848 _0146_ _0196_ 0
C20849 clknet_1_0__leaf__0463_ _1046_/a_561_413# 0
C20850 _0811_/a_81_21# _0345_ 0.00869f
C20851 net82 _0185_ 0
C20852 _0398_ _0394_ 0
C20853 _0096_ _0306_ 0
C20854 net10 _0449_ 0
C20855 _0183_ _0116_ 0.02313f
C20856 _0176_ _0548_/a_240_47# 0.00163f
C20857 _1000_/a_634_159# _0393_ 0
C20858 _0412_ _0799_/a_80_21# 0
C20859 _0800_/a_51_297# _0411_ 0.00152f
C20860 comp0.B\[12\] _1044_/a_193_47# 0
C20861 _0680_/a_80_21# _0238_ 0.07921f
C20862 _0924_/a_27_47# _0935_/a_27_47# 0.01126f
C20863 _0268_ _0444_ 0
C20864 _1066_/a_27_47# net17 0
C20865 net207 _0580_/a_27_297# 0
C20866 _0254_ _0622_/a_109_47# 0.01114f
C20867 clknet_1_0__leaf__0458_ _1014_/a_466_413# 0
C20868 _0486_ _0484_ 0
C20869 control0.state\[2\] _0485_ 0.31319f
C20870 _0592_/a_68_297# _0592_/a_150_297# 0.00477f
C20871 control0.count\[1\] _1069_/a_592_47# 0
C20872 VPWR _0167_ 0.53472f
C20873 hold39/a_285_47# clknet_1_1__leaf__0463_ 0.01117f
C20874 _0619_/a_68_297# _0619_/a_150_297# 0.00477f
C20875 comp0.B\[2\] _0473_ 0
C20876 A[0] input17/a_75_212# 0.00319f
C20877 input1/a_27_47# B[0] 0.00125f
C20878 acc0.A\[20\] net48 0.58445f
C20879 comp0.B\[12\] net131 0.00124f
C20880 _1018_/a_891_413# _0218_ 0.00192f
C20881 _0397_ _0218_ 0
C20882 _1030_/a_891_413# _0220_ 0.00605f
C20883 _1030_/a_1059_315# _0336_ 0.02346f
C20884 _0414_ _0994_/a_193_47# 0
C20885 net235 _0181_ 0
C20886 hold30/a_391_47# net110 0
C20887 _0323_ _0743_/a_240_47# 0
C20888 _0172_ hold1/a_285_47# 0
C20889 _0369_ _1005_/a_1059_315# 0
C20890 _1017_/a_634_159# clknet_1_1__leaf__0461_ 0
C20891 _0216_ _1011_/a_381_47# 0.0039f
C20892 _1000_/a_891_413# _0245_ 0
C20893 _0216_ _1006_/a_193_47# 0.02058f
C20894 _0343_ _0218_ 0.74295f
C20895 _0462_ _0318_ 0
C20896 _0199_ _0146_ 0
C20897 _1006_/a_466_413# net92 0
C20898 _0656_/a_145_75# _0288_ 0
C20899 _0143_ VPWR 0.30845f
C20900 _0993_/a_381_47# net246 0
C20901 VPWR _0880_/a_27_47# 0.23988f
C20902 _0570_/a_27_297# hold9/a_285_47# 0.00104f
C20903 net59 _0341_ 0
C20904 _0984_/a_381_47# _0984_/a_561_413# 0.00123f
C20905 _0984_/a_27_47# net70 0.22753f
C20906 _0984_/a_891_413# _0984_/a_975_413# 0.00851f
C20907 _0201_ net129 0
C20908 _0200_ hold6/a_49_47# 0
C20909 _1031_/a_381_47# _0219_ 0
C20910 _0216_ acc0.A\[25\] 0.28243f
C20911 net79 _0419_ 0
C20912 _0808_/a_368_297# _0091_ 0
C20913 clkload3/Y _1017_/a_27_47# 0
C20914 _0439_ _0988_/a_193_47# 0.00144f
C20915 acc0.A\[19\] net223 0.01038f
C20916 net43 net219 0
C20917 _0765_/a_79_21# _0369_ 0.13639f
C20918 net122 input28/a_75_212# 0.00149f
C20919 net234 _0459_ 0
C20920 VPWR _0988_/a_193_47# 0.29903f
C20921 _0514_/a_109_297# acc0.A\[10\] 0.0015f
C20922 _0390_ acc0.A\[20\] 0
C20923 hold97/a_391_47# _0106_ 0
C20924 pp[10] acc0.A\[11\] 0
C20925 _0474_ hold84/a_285_47# 0
C20926 _1015_/a_27_47# clknet_1_0__leaf__0457_ 0
C20927 _1059_/a_27_47# _0184_ 0.00246f
C20928 _0285_ hold81/a_285_47# 0
C20929 _0344_ _1031_/a_27_47# 0
C20930 _0730_/a_510_47# VPWR 0
C20931 hold78/a_285_47# _1031_/a_1059_315# 0
C20932 _1058_/a_1059_315# _0281_ 0
C20933 net168 _1054_/a_466_413# 0.01442f
C20934 _0463_ _0138_ 0
C20935 VPWR _0953_/a_32_297# 0.35491f
C20936 net12 net73 0
C20937 _1056_/a_634_159# _0186_ 0.00599f
C20938 VPWR hold92/a_391_47# 0.20383f
C20939 _0857_/a_27_47# VPWR 0.27212f
C20940 net46 _0459_ 0
C20941 net103 _0181_ 0.03729f
C20942 _1023_/a_381_47# net109 0
C20943 _1023_/a_891_413# net177 0.00204f
C20944 _1023_/a_634_159# acc0.A\[23\] 0
C20945 _1037_/a_891_413# _0175_ 0.00121f
C20946 _0300_ _0301_ 0
C20947 _0369_ _1006_/a_634_159# 0
C20948 hold32/a_391_47# A[10] 0
C20949 net59 _0722_/a_79_21# 0
C20950 _0697_/a_217_297# _0686_/a_27_53# 0
C20951 _0195_ _0571_/a_109_47# 0.00346f
C20952 _0216_ _0571_/a_27_297# 0.20886f
C20953 net155 _0571_/a_109_297# 0.00291f
C20954 _0467_ _0487_ 0.45978f
C20955 clknet_1_0__leaf__0465_ _0837_/a_81_21# 0.00129f
C20956 _1011_/a_1059_315# _0335_ 0
C20957 output67/a_27_47# VPWR 0.33464f
C20958 _0433_ _0186_ 0.38495f
C20959 clkbuf_1_1__f__0462_/a_110_47# _0690_/a_68_297# 0.00131f
C20960 _1037_/a_381_47# control0.sh 0
C20961 _0217_ _0721_/a_27_47# 0
C20962 _0337_ hold62/a_49_47# 0.01077f
C20963 _0257_ acc0.A\[6\] 0
C20964 _0757_/a_68_297# _0378_ 0
C20965 _0350_ _0756_/a_47_47# 0
C20966 _1016_/a_27_47# _0307_ 0
C20967 _0263_ _0842_/a_59_75# 0.13141f
C20968 _0119_ net118 0
C20969 VPWR net72 0.3159f
C20970 _0399_ _0434_ 0.0841f
C20971 _1001_/a_193_47# VPWR 0.3003f
C20972 hold36/a_391_47# clkbuf_0__0464_/a_110_47# 0.0049f
C20973 _0129_ _1031_/a_891_413# 0.01053f
C20974 net163 _1031_/a_466_413# 0.00296f
C20975 net7 _0176_ 0.02405f
C20976 acc0.A\[16\] _0781_/a_150_297# 0
C20977 _0988_/a_193_47# output62/a_27_47# 0
C20978 VPWR _1062_/a_27_47# 0.6398f
C20979 _0342_ _0195_ 0.01595f
C20980 _0616_/a_78_199# _0247_ 0.20562f
C20981 _1059_/a_891_413# net229 0
C20982 _0128_ hold61/a_391_47# 0.01879f
C20983 _0148_ clknet_1_1__leaf__0464_ 0
C20984 clkbuf_1_1__f_clk/a_110_47# net107 0.00191f
C20985 output57/a_27_47# net57 0.2163f
C20986 _1038_/a_1059_315# _1037_/a_891_413# 0
C20987 _1038_/a_891_413# _1037_/a_1059_315# 0.00119f
C20988 clkbuf_1_0__f__0457_/a_110_47# _0616_/a_78_199# 0
C20989 VPWR hold8/a_285_47# 0.2878f
C20990 _0490_ _0488_ 0.0747f
C20991 clkbuf_0__0457_/a_110_47# hold40/a_391_47# 0
C20992 _0487_ comp0.B\[0\] 0
C20993 _0997_/a_891_413# _0095_ 0
C20994 comp0.B\[6\] _0549_/a_68_297# 0.0017f
C20995 comp0.B\[5\] _0549_/a_150_297# 0
C20996 _0677_/a_47_47# _0393_ 0
C20997 net234 _0265_ 0.15738f
C20998 _0165_ _0163_ 0
C20999 net193 hold6/a_49_47# 0
C21000 _0111_ pp[31] 0
C21001 acc0.A\[20\] clknet_1_0__leaf__0459_ 0.00115f
C21002 _0743_/a_240_47# net237 0.05932f
C21003 _1053_/a_634_159# hold83/a_49_47# 0.00127f
C21004 _1053_/a_27_47# hold83/a_391_47# 0.00249f
C21005 _1053_/a_193_47# hold83/a_285_47# 0.00356f
C21006 _0195_ _0334_ 0.06447f
C21007 net42 pp[14] 0
C21008 _1065_/a_634_159# _1065_/a_466_413# 0.23992f
C21009 _1065_/a_193_47# _1065_/a_1059_315# 0.03405f
C21010 _1065_/a_27_47# _1065_/a_891_413# 0.03089f
C21011 _0395_ _0306_ 0
C21012 VPWR _0561_/a_51_297# 0.47233f
C21013 _0217_ _0760_/a_285_47# 0.0016f
C21014 _0183_ _0760_/a_377_297# 0.00152f
C21015 net232 _1066_/a_1059_315# 0
C21016 _0121_ _0183_ 0.19945f
C21017 _0787_/a_209_297# _0418_ 0
C21018 _0787_/a_303_47# _0281_ 0.00169f
C21019 _0251_ net169 0
C21020 _0998_/a_193_47# _0218_ 0.0065f
C21021 _1036_/a_466_413# _1035_/a_27_47# 0.00205f
C21022 _0571_/a_373_47# _0125_ 0
C21023 clknet_0__0464_ net157 0
C21024 net202 _1067_/a_891_413# 0
C21025 _0601_/a_150_297# acc0.A\[23\] 0
C21026 _1003_/a_27_47# _0228_ 0
C21027 _0985_/a_193_47# _0270_ 0
C21028 _0776_/a_27_47# _0219_ 0.00407f
C21029 _0707_/a_75_199# _0707_/a_544_297# 0.01759f
C21030 _1033_/a_1059_315# _0565_/a_149_47# 0
C21031 hold79/a_285_47# _1070_/a_27_47# 0
C21032 hold79/a_49_47# _1070_/a_193_47# 0
C21033 _0954_/a_220_297# _1042_/a_193_47# 0
C21034 _1014_/a_27_47# _1014_/a_193_47# 0.96236f
C21035 clknet_1_1__leaf__0463_ _1067_/a_891_413# 0.00104f
C21036 _0508_/a_299_297# hold82/a_285_47# 0.00142f
C21037 VPWR _1047_/a_634_159# 0.18719f
C21038 _0811_/a_299_297# _0811_/a_384_47# 0
C21039 hold17/a_391_47# clknet_1_0__leaf_clk 0.00435f
C21040 _0285_ _0282_ 0
C21041 _0627_/a_109_93# clknet_0__0465_ 0.00592f
C21042 _0195_ _1013_/a_592_47# 0.00112f
C21043 _0238_ _0248_ 0.17427f
C21044 _0457_ _0526_/a_27_47# 0
C21045 output67/a_27_47# input4/a_75_212# 0
C21046 input5/a_75_212# net5 0.1085f
C21047 A[13] acc0.A\[13\] 0.00506f
C21048 output55/a_27_47# net59 0
C21049 net133 _0147_ 0
C21050 hold101/a_285_47# hold101/a_391_47# 0.41909f
C21051 net173 net152 0
C21052 _0399_ acc0.A\[7\] 0
C21053 hold57/a_391_47# net8 0
C21054 VPWR _1007_/a_891_413# 0.18755f
C21055 _0996_/a_27_47# _0459_ 0.00137f
C21056 VPWR _0133_ 0.82663f
C21057 _0172_ _1040_/a_561_413# 0
C21058 _0550_/a_240_47# net174 0
C21059 _1058_/a_561_413# VPWR 0.00292f
C21060 _0179_ _1051_/a_1059_315# 0
C21061 _0467_ net119 0.00141f
C21062 net68 _0181_ 0.14017f
C21063 _0534_/a_384_47# acc0.A\[15\] 0.00147f
C21064 net61 hold65/a_49_47# 0.00676f
C21065 _0179_ net139 0
C21066 _0493_/a_27_47# _0208_ 0
C21067 _0171_ _0213_ 0
C21068 _0404_ _0301_ 0
C21069 _0279_ acc0.A\[13\] 0
C21070 _1055_/a_193_47# net16 0.0119f
C21071 _0316_ _0698_/a_199_47# 0
C21072 _1064_/a_1059_315# _1064_/a_1017_47# 0
C21073 _0558_/a_68_297# VPWR 0.19528f
C21074 acc0.A\[27\] _0321_ 0
C21075 _0275_ _0431_ 0.04916f
C21076 clknet_1_0__leaf__0458_ _0852_/a_285_47# 0
C21077 _0728_/a_59_75# _0219_ 0.05103f
C21078 acc0.A\[27\] clkbuf_0__0460_/a_110_47# 0
C21079 output52/a_27_47# net52 0.20296f
C21080 clk _0166_ 0
C21081 _0669_/a_29_53# _0669_/a_183_297# 0.00868f
C21082 _1018_/a_27_47# net103 0
C21083 hold41/a_49_47# A[11] 0
C21084 pp[15] _0345_ 0
C21085 clknet_1_1__leaf_clk _1063_/a_381_47# 0
C21086 _0218_ net38 0.00188f
C21087 net112 _1025_/a_193_47# 0.00979f
C21088 VPWR hold80/a_391_47# 0.19214f
C21089 _0712_/a_79_21# _0344_ 0.13832f
C21090 _1002_/a_27_47# _1067_/a_891_413# 0.00153f
C21091 A[14] _0218_ 0
C21092 output37/a_27_47# clknet_1_1__leaf__0465_ 0.00111f
C21093 clkbuf_1_0__f__0459_/a_110_47# _1060_/a_891_413# 0.00735f
C21094 net137 net148 0
C21095 _0983_/a_891_413# net221 0
C21096 _0343_ _1017_/a_975_413# 0
C21097 _1002_/a_1059_315# _0383_ 0
C21098 _1002_/a_381_47# _0369_ 0
C21099 _0234_ _0227_ 0.1653f
C21100 _1025_/a_193_47# acc0.A\[24\] 0.00294f
C21101 net230 hold83/a_285_47# 0.01016f
C21102 _0192_ hold83/a_391_47# 0
C21103 net119 comp0.B\[0\] 0.03081f
C21104 _1056_/a_891_413# _1056_/a_975_413# 0.00851f
C21105 _0257_ _0624_/a_59_75# 0.02222f
C21106 control0.state\[1\] _0967_/a_487_297# 0
C21107 _0226_ _0374_ 0.02168f
C21108 hold65/a_391_47# net63 0
C21109 net43 _0352_ 0.35593f
C21110 _0181_ net143 0.03373f
C21111 _0985_/a_466_413# net61 0
C21112 _1013_/a_466_413# _0339_ 0
C21113 _0636_/a_145_75# _0186_ 0
C21114 hold24/a_285_47# clkbuf_1_0__f__0463_/a_110_47# 0.02321f
C21115 net11 acc0.A\[6\] 0.03975f
C21116 _0457_ _0175_ 0
C21117 _0352_ hold73/a_285_47# 0.00251f
C21118 _0429_ acc0.A\[6\] 0
C21119 pp[27] net57 0.16944f
C21120 _0393_ _0242_ 0.06127f
C21121 _0321_ _0364_ 0.43f
C21122 hold13/a_285_47# comp0.B\[2\] 0
C21123 _0222_ _1022_/a_193_47# 0.05709f
C21124 _0855_/a_81_21# net149 0.09825f
C21125 _0259_ _0088_ 0
C21126 _0854_/a_215_47# _0455_ 0.00837f
C21127 _0854_/a_79_21# _0081_ 0.05088f
C21128 _1037_/a_27_47# _1036_/a_27_47# 0
C21129 VPWR net107 0.4114f
C21130 _0322_ _0329_ 0.05704f
C21131 _0350_ _0084_ 0
C21132 hold21/a_49_47# net12 0
C21133 _0648_/a_27_297# clkbuf_1_1__f__0459_/a_110_47# 0.01056f
C21134 _1058_/a_1059_315# A[12] 0
C21135 _0999_/a_27_47# _0352_ 0.22041f
C21136 _0329_ _0327_ 0.36532f
C21137 _0413_ _0997_/a_466_413# 0.00127f
C21138 hold28/a_285_47# net175 0.04257f
C21139 _0498_/a_51_297# _0498_/a_240_47# 0.03076f
C21140 _0830_/a_510_47# _0437_ 0.003f
C21141 comp0.B\[4\] hold84/a_49_47# 0
C21142 _0841_/a_79_21# _0986_/a_193_47# 0.00378f
C21143 clknet_1_1__leaf__0460_ _1028_/a_193_47# 0
C21144 A[10] _0153_ 0.0047f
C21145 net35 clkbuf_1_0__f_clk/a_110_47# 0.0038f
C21146 _0179_ _0422_ 0.03055f
C21147 net10 _0540_/a_51_297# 0
C21148 _0313_ hold97/a_285_47# 0
C21149 _1015_/a_891_413# clknet_1_0__leaf__0461_ 0.00276f
C21150 net82 clknet_0__0459_ 0.04607f
C21151 _1034_/a_193_47# _0131_ 0
C21152 clknet_1_0__leaf__0465_ _1052_/a_592_47# 0
C21153 net36 _1040_/a_27_47# 0
C21154 _0442_ acc0.A\[4\] 0.00105f
C21155 net197 _1028_/a_27_47# 0
C21156 _0287_ _0402_ 0
C21157 _0195_ _1014_/a_193_47# 0
C21158 hold11/a_285_47# net10 0
C21159 _0180_ _0524_/a_109_297# 0.01796f
C21160 comp0.B\[11\] _0176_ 0.26401f
C21161 _0516_/a_373_47# net142 0
C21162 clknet_1_0__leaf__0458_ _0844_/a_297_47# 0
C21163 hold51/a_285_47# hold51/a_391_47# 0.41909f
C21164 _0351_ _0110_ 0
C21165 _0856_/a_79_21# _1014_/a_1059_315# 0
C21166 net11 _0523_/a_384_47# 0
C21167 _0260_ net10 0
C21168 clkbuf_1_0__f__0460_/a_110_47# _0373_ 0
C21169 _0368_ _0352_ 0.03863f
C21170 _1001_/a_193_47# clknet_1_0__leaf__0459_ 0
C21171 _0327_ _0221_ 0.12708f
C21172 clkbuf_1_0__f__0457_/a_110_47# _0384_ 0
C21173 _0512_/a_373_47# _0181_ 0.00165f
C21174 control0.sh _1062_/a_381_47# 0
C21175 _1018_/a_193_47# net219 0.00111f
C21176 net146 _0185_ 0.0045f
C21177 _0727_/a_109_47# _0333_ 0
C21178 _0356_ _0701_/a_80_21# 0
C21179 _1008_/a_27_47# _1008_/a_1059_315# 0.04875f
C21180 _1008_/a_193_47# _1008_/a_466_413# 0.07482f
C21181 _0416_ acc0.A\[13\] 0
C21182 _0488_ _1069_/a_381_47# 0
C21183 _0466_ _1069_/a_891_413# 0
C21184 _0976_/a_76_199# control0.count\[0\] 0.36904f
C21185 hold16/a_285_47# net163 0.01002f
C21186 output56/a_27_47# pp[28] 0.15844f
C21187 _1020_/a_634_159# _1020_/a_592_47# 0
C21188 output43/a_27_47# _0995_/a_27_47# 0
C21189 hold76/a_285_47# net211 0
C21190 _1002_/a_1017_47# _0100_ 0.00109f
C21191 acc0.A\[23\] _0377_ 0
C21192 _0400_ _0406_ 0.27046f
C21193 _0408_ net42 0.18329f
C21194 _0182_ _0448_ 0
C21195 _1035_/a_27_47# comp0.B\[6\] 0
C21196 _1035_/a_193_47# comp0.B\[5\] 0
C21197 _1035_/a_466_413# comp0.B\[3\] 0
C21198 clkbuf_1_0__f__0464_/a_110_47# _1049_/a_891_413# 0.00846f
C21199 _0239_ _0607_/a_109_297# 0.0038f
C21200 _1055_/a_27_47# _0515_/a_81_21# 0
C21201 output59/a_27_47# _0195_ 0.01119f
C21202 _0311_ _0326_ 0
C21203 _0483_ clkbuf_0_clk/a_110_47# 0
C21204 hold28/a_391_47# _0147_ 0.04376f
C21205 _0746_/a_81_21# _0219_ 0
C21206 clknet_0__0458_ _0986_/a_27_47# 0.00797f
C21207 acc0.A\[27\] _1009_/a_27_47# 0
C21208 _0217_ clkbuf_1_0__f__0461_/a_110_47# 0
C21209 _1028_/a_381_47# hold50/a_49_47# 0.00167f
C21210 clknet_0__0457_ _1014_/a_27_47# 0.01698f
C21211 _0183_ _0380_ 0
C21212 _0515_/a_299_297# _0515_/a_384_47# 0
C21213 _0475_ _0175_ 0.23306f
C21214 _0188_ _0512_/a_109_47# 0
C21215 _0346_ _0304_ 0.50082f
C21216 _1031_/a_891_413# hold61/a_285_47# 0
C21217 _0411_ _0277_ 0
C21218 _1013_/a_1059_315# net99 0
C21219 net46 _0772_/a_79_21# 0.01379f
C21220 hold14/a_49_47# VPWR 0.27727f
C21221 _0313_ _0366_ 0.10857f
C21222 _0314_ _0315_ 0.39903f
C21223 _1041_/a_634_159# _0172_ 0.01843f
C21224 _1041_/a_1059_315# net180 0
C21225 _1041_/a_466_413# net30 0
C21226 _0452_ _0635_/a_27_47# 0
C21227 _0559_/a_245_297# _0133_ 0
C21228 control0.count\[3\] net159 0
C21229 _0109_ hold80/a_49_47# 0
C21230 _0992_/a_634_159# _0345_ 0
C21231 _0645_/a_285_47# net41 0.06705f
C21232 clkbuf_1_1__f__0457_/a_110_47# hold71/a_285_47# 0
C21233 _0195_ _0724_/a_113_297# 0.01358f
C21234 hold94/a_391_47# _0754_/a_240_47# 0
C21235 hold21/a_391_47# input15/a_75_212# 0.01627f
C21236 _0991_/a_193_47# acc0.A\[15\] 0
C21237 _0838_/a_109_297# _0271_ 0
C21238 _0441_ _1051_/a_1059_315# 0
C21239 clknet_0__0459_ _0796_/a_297_297# 0
C21240 _0176_ _0202_ 0.80774f
C21241 hold63/a_285_47# net53 0
C21242 _1072_/a_891_413# _0468_ 0
C21243 _0226_ _0249_ 0
C21244 hold42/a_391_47# _1058_/a_27_47# 0.00609f
C21245 hold42/a_285_47# _1058_/a_193_47# 0.00661f
C21246 net26 _0549_/a_68_297# 0
C21247 VPWR _0535_/a_68_297# 0.15735f
C21248 net86 _0393_ 0.11854f
C21249 _0578_/a_27_297# net150 0.09077f
C21250 _1058_/a_27_47# _1057_/a_891_413# 0.00868f
C21251 _1058_/a_193_47# _1057_/a_1059_315# 0
C21252 _1058_/a_634_159# _1057_/a_466_413# 0.012f
C21253 _1058_/a_891_413# _1057_/a_27_47# 0.00868f
C21254 _1058_/a_466_413# _1057_/a_634_159# 0.012f
C21255 _1058_/a_1059_315# _1057_/a_193_47# 0
C21256 VPWR _0336_ 0.3834f
C21257 _0083_ _0446_ 0
C21258 clknet_1_1__leaf__0460_ net216 0.0512f
C21259 _0403_ net246 0
C21260 _0458_ _0530_/a_299_297# 0
C21261 net207 _0117_ 0
C21262 clk _0168_ 0
C21263 B[9] hold5/a_391_47# 0.00247f
C21264 pp[16] _0095_ 0
C21265 _0218_ _0793_/a_51_297# 0
C21266 _0428_ _0345_ 0
C21267 net168 hold22/a_49_47# 0.03441f
C21268 _0946_/a_30_53# net1 0
C21269 net35 control0.count\[2\] 0.0103f
C21270 _0576_/a_27_297# clknet_1_0__leaf__0460_ 0.00125f
C21271 _1000_/a_561_413# _0347_ 0.00156f
C21272 _1000_/a_1059_315# _0352_ 0.00629f
C21273 net185 control0.sh 0.03603f
C21274 VPWR _1063_/a_561_413# 0.00213f
C21275 _0284_ _0654_/a_207_413# 0.06788f
C21276 net103 clknet_1_1__leaf__0461_ 0.13781f
C21277 _0216_ net57 0.00226f
C21278 _0195_ net155 0.38088f
C21279 net210 _0216_ 0.00871f
C21280 clkbuf_0__0457_/a_110_47# acc0.A\[19\] 0.00111f
C21281 VPWR _0959_/a_300_47# 0
C21282 hold36/a_285_47# _0473_ 0
C21283 VPWR _0585_/a_109_47# 0
C21284 clknet_1_1__leaf__0458_ acc0.A\[6\] 0.84088f
C21285 net46 net51 0.11212f
C21286 _0739_/a_79_21# hold50/a_285_47# 0
C21287 _0126_ hold9/a_285_47# 0.04981f
C21288 _0443_ _0444_ 0.16884f
C21289 clknet_0__0458_ clknet_1_0__leaf__0458_ 0.02413f
C21290 _0286_ _0420_ 0
C21291 _0275_ _0269_ 0.13072f
C21292 _0347_ hold50/a_391_47# 0.05815f
C21293 _0130_ net118 0
C21294 _0548_/a_51_297# _0548_/a_149_47# 0.02487f
C21295 VPWR _1060_/a_561_413# 0.00358f
C21296 net114 net244 0
C21297 pp[28] _0707_/a_315_47# 0
C21298 clkload1/a_110_47# _0346_ 0
C21299 _1056_/a_27_47# A[10] 0
C21300 _0584_/a_109_297# _0208_ 0
C21301 hold65/a_285_47# clkbuf_1_0__f__0465_/a_110_47# 0.00359f
C21302 _0179_ acc0.A\[8\] 0.02769f
C21303 hold36/a_285_47# clkbuf_1_1__f__0464_/a_110_47# 0
C21304 clknet_0_clk _1063_/a_27_47# 0.01181f
C21305 _0985_/a_193_47# hold23/a_49_47# 0.00243f
C21306 _0985_/a_27_47# hold23/a_285_47# 0.0016f
C21307 VPWR _0174_ 2.93239f
C21308 hold2/a_49_47# hold60/a_391_47# 0
C21309 net168 net169 0.28344f
C21310 _0174_ _1043_/a_561_413# 0
C21311 VPWR _1050_/a_27_47# 0.69445f
C21312 clkbuf_0__0458_/a_110_47# _0447_ 0.00463f
C21313 _0195_ _0240_ 0
C21314 clknet_0_clk _0974_/a_448_47# 0.00259f
C21315 _0511_/a_81_21# _0511_/a_384_47# 0.00138f
C21316 _0452_ _0850_/a_68_297# 0.10698f
C21317 hold89/a_391_47# _0486_ 0.00136f
C21318 hold21/a_49_47# pp[5] 0.00315f
C21319 net109 acc0.A\[23\] 0
C21320 acc0.A\[7\] _0619_/a_68_297# 0.17492f
C21321 pp[9] input16/a_75_212# 0.01585f
C21322 _0195_ _0369_ 0.01992f
C21323 _0331_ clknet_1_1__leaf__0462_ 0.22661f
C21324 _0179_ _0991_/a_193_47# 0
C21325 net206 _0242_ 0
C21326 clknet_0__0457_ _0195_ 0.01205f
C21327 _0369_ net92 0
C21328 _0715_/a_27_47# _0345_ 0
C21329 _1044_/a_1017_47# net20 0.00184f
C21330 _0557_/a_51_297# net28 0
C21331 pp[27] _1010_/a_1059_315# 0
C21332 _0217_ _0182_ 0.01667f
C21333 _0298_ _0411_ 0.27035f
C21334 hold36/a_285_47# _0186_ 0
C21335 pp[15] _0791_/a_113_297# 0
C21336 _0216_ _0125_ 0.04483f
C21337 net69 _1060_/a_27_47# 0
C21338 _0457_ _1015_/a_592_47# 0.00113f
C21339 _0532_/a_81_21# _1048_/a_891_413# 0.00357f
C21340 _0198_ _1048_/a_27_47# 0
C21341 _0536_/a_51_297# net157 0.12984f
C21342 _0195_ _0852_/a_117_297# 0
C21343 _1037_/a_592_47# B[6] 0
C21344 hold18/a_285_47# net247 0.06076f
C21345 VPWR _0772_/a_297_297# 0.00781f
C21346 clkbuf_1_0__f__0463_/a_110_47# _0138_ 0
C21347 _0248_ clkbuf_1_0__f__0461_/a_110_47# 0
C21348 _0376_ _0606_/a_109_53# 0
C21349 net45 _1017_/a_1017_47# 0
C21350 _1020_/a_193_47# _0461_ 0.00176f
C21351 _1020_/a_381_47# _0891_/a_27_47# 0
C21352 _1018_/a_1059_315# _0347_ 0.01285f
C21353 _0578_/a_27_297# control0.add 0.04919f
C21354 _1039_/a_1017_47# _0172_ 0
C21355 _1021_/a_592_47# VPWR 0
C21356 net172 _1037_/a_381_47# 0
C21357 net55 net95 0
C21358 _0305_ _0663_/a_207_413# 0
C21359 _0762_/a_510_47# _0383_ 0.00898f
C21360 net180 _0953_/a_114_297# 0.00179f
C21361 net84 _0796_/a_510_47# 0
C21362 _0365_ net244 0
C21363 hold65/a_49_47# _0431_ 0
C21364 _1000_/a_634_159# _0773_/a_35_297# 0.00318f
C21365 clknet_1_1__leaf__0459_ acc0.A\[14\] 0
C21366 net56 _0720_/a_150_297# 0
C21367 net149 _0566_/a_27_47# 0
C21368 _0346_ _0811_/a_384_47# 0
C21369 _1009_/a_27_47# _1009_/a_634_159# 0.14145f
C21370 _0308_ _0394_ 0.45819f
C21371 VPWR _0518_/a_27_297# 0.21056f
C21372 net36 _1061_/a_466_413# 0
C21373 _0576_/a_27_297# _0576_/a_109_297# 0.17136f
C21374 _0295_ _0421_ 0
C21375 pp[10] A[12] 0.03889f
C21376 hold35/a_49_47# _0186_ 0
C21377 _0642_/a_298_297# VPWR 0.19957f
C21378 VPWR _0208_ 3.02905f
C21379 hold5/a_285_47# _0204_ 0
C21380 net27 _0175_ 0.12122f
C21381 _0677_/a_129_47# _0352_ 0
C21382 _0313_ _0689_/a_68_297# 0.00557f
C21383 net36 net171 0.03886f
C21384 clknet_0_clk _1062_/a_1059_315# 0.03972f
C21385 hold66/a_49_47# _1005_/a_381_47# 0
C21386 _1036_/a_193_47# net121 0.03572f
C21387 _1036_/a_27_47# _0133_ 0.00123f
C21388 _0186_ _0522_/a_109_47# 0.0033f
C21389 net111 _1025_/a_193_47# 0.00677f
C21390 _1036_/a_891_413# B[15] 0
C21391 _1068_/a_381_47# _0487_ 0
C21392 _0967_/a_109_93# net1 0.03793f
C21393 net1 _0487_ 0.04604f
C21394 _0992_/a_1059_315# _0811_/a_299_297# 0
C21395 _0992_/a_891_413# _0811_/a_81_21# 0
C21396 _0707_/a_544_297# _0338_ 0.00226f
C21397 _0707_/a_201_297# _0339_ 0.02047f
C21398 _0218_ _0842_/a_59_75# 0.01847f
C21399 hold79/a_49_47# VPWR 0.32246f
C21400 net64 _0179_ 0
C21401 comp0.B\[11\] _1042_/a_975_413# 0
C21402 _0389_ _0241_ 0.22112f
C21403 _1014_/a_466_413# _1014_/a_592_47# 0.00553f
C21404 _1014_/a_634_159# _1014_/a_1017_47# 0
C21405 _1071_/a_634_159# _1071_/a_1059_315# 0
C21406 _1071_/a_27_47# _1071_/a_381_47# 0.06222f
C21407 _1071_/a_193_47# _1071_/a_891_413# 0.19497f
C21408 _0187_ net143 0.0034f
C21409 net59 acc0.A\[30\] 0.21561f
C21410 _1015_/a_466_413# _0208_ 0.04248f
C21411 _0331_ net242 0
C21412 hold96/a_49_47# hold96/a_285_47# 0.22264f
C21413 _0985_/a_561_413# _0458_ 0
C21414 net61 _0828_/a_199_47# 0
C21415 _0852_/a_35_297# _0852_/a_117_297# 0.00641f
C21416 _0476_ _1034_/a_891_413# 0
C21417 _0179_ _0423_ 0.01162f
C21418 _0233_ _0230_ 0.21304f
C21419 _0343_ _0792_/a_80_21# 0.14629f
C21420 _0458_ _1049_/a_1059_315# 0
C21421 _0183_ _0386_ 0
C21422 _0251_ _0830_/a_79_21# 0
C21423 _1035_/a_27_47# net26 0.02393f
C21424 _0346_ clknet_1_0__leaf__0460_ 0.02031f
C21425 VPWR B[0] 0.26075f
C21426 net139 input13/a_75_212# 0
C21427 _0815_/a_113_297# _0181_ 0.00867f
C21428 clknet_1_0__leaf__0463_ _0463_ 0.00591f
C21429 _0226_ net1 0
C21430 _0436_ pp[3] 0
C21431 _0437_ _0989_/a_193_47# 0.03869f
C21432 net212 _0989_/a_634_159# 0
C21433 hold25/a_285_47# hold25/a_391_47# 0.41909f
C21434 net188 net2 0
C21435 hold98/a_285_47# net41 0.00103f
C21436 _0857_/a_27_47# comp0.B\[3\] 0
C21437 _0381_ hold73/a_391_47# 0
C21438 _1015_/a_634_159# net17 0
C21439 _0284_ _0286_ 0.06599f
C21440 _1026_/a_975_413# acc0.A\[25\] 0
C21441 _0455_ _0852_/a_285_47# 0
C21442 net36 _1039_/a_466_413# 0.03335f
C21443 _0295_ _0809_/a_81_21# 0.06036f
C21444 _0778_/a_68_297# _0395_ 0
C21445 acc0.A\[29\] _0705_/a_59_75# 0
C21446 net88 _1067_/a_466_413# 0
C21447 _0195_ _1048_/a_634_159# 0
C21448 hold18/a_391_47# _0846_/a_240_47# 0
C21449 _0343_ output64/a_27_47# 0
C21450 _1012_/a_634_159# _0352_ 0.01825f
C21451 net54 hold9/a_285_47# 0.02943f
C21452 _0819_/a_81_21# _0428_ 0.13985f
C21453 _0819_/a_299_297# _0427_ 0.04683f
C21454 clknet_0__0459_ net146 0.00147f
C21455 clknet_1_0__leaf__0460_ hold94/a_49_47# 0
C21456 _0183_ _1059_/a_975_413# 0
C21457 _0343_ _1016_/a_1059_315# 0.0084f
C21458 _0288_ net229 0
C21459 _0083_ net61 0.25462f
C21460 clknet_1_0__leaf__0465_ hold83/a_391_47# 0
C21461 clkbuf_0__0461_/a_110_47# _0218_ 0.09773f
C21462 _0579_/a_27_297# clknet_1_0__leaf__0457_ 0
C21463 _0216_ _1010_/a_1059_315# 0
C21464 _0981_/a_373_47# net167 0.003f
C21465 _0981_/a_27_297# _0170_ 0.11027f
C21466 _1052_/a_1059_315# _0180_ 0
C21467 _0521_/a_81_21# VPWR 0.23151f
C21468 _0148_ net148 0
C21469 net102 _1060_/a_27_47# 0
C21470 hold49/a_391_47# net196 0.13054f
C21471 _1016_/a_466_413# acc0.A\[17\] 0
C21472 hold20/a_49_47# control0.count\[3\] 0.30118f
C21473 _0963_/a_285_297# control0.count\[1\] 0.0129f
C21474 _0998_/a_27_47# _0347_ 0
C21475 _0273_ _0436_ 0.00389f
C21476 _0255_ _0831_/a_35_297# 0
C21477 net36 _0634_/a_113_47# 0
C21478 _0533_/a_109_297# _0181_ 0.01019f
C21479 _0232_ _0366_ 0
C21480 _0424_ _0401_ 0.0334f
C21481 _0280_ clkbuf_1_1__f__0459_/a_110_47# 0.09472f
C21482 hold23/a_285_47# _0197_ 0.03492f
C21483 comp0.B\[2\] net25 0
C21484 _0313_ acc0.A\[24\] 0
C21485 acc0.A\[16\] _0678_/a_68_297# 0
C21486 _0498_/a_512_297# _0159_ 0
C21487 _0234_ _0352_ 0.18466f
C21488 _0084_ _0986_/a_634_159# 0.00894f
C21489 _0445_ _0986_/a_1059_315# 0
C21490 hold96/a_285_47# net90 0
C21491 _0358_ acc0.A\[29\] 0.00204f
C21492 _0592_/a_68_297# _0756_/a_47_47# 0.0279f
C21493 _0399_ _0988_/a_466_413# 0.00167f
C21494 hold96/a_49_47# _1024_/a_27_47# 0
C21495 _1053_/a_27_47# net9 0
C21496 _1038_/a_1059_315# _0136_ 0.03643f
C21497 net172 _0553_/a_149_47# 0
C21498 comp0.B\[2\] _1033_/a_592_47# 0.00112f
C21499 _0557_/a_240_47# _0134_ 0
C21500 _0577_/a_27_297# _0103_ 0
C21501 net190 _1028_/a_592_47# 0.00164f
C21502 _0126_ _1028_/a_381_47# 0.11511f
C21503 clknet_1_1__leaf__0459_ _0798_/a_199_47# 0
C21504 net1 clkbuf_0__0457_/a_110_47# 0.00785f
C21505 comp0.B\[13\] VPWR 0.7472f
C21506 _0715_/a_27_47# _0819_/a_81_21# 0
C21507 clknet_1_1__leaf__0462_ _1008_/a_27_47# 0.00896f
C21508 hold42/a_285_47# pp[9] 0.00131f
C21509 comp0.B\[3\] _0561_/a_51_297# 0.00194f
C21510 VPWR A[13] 0.42496f
C21511 _1032_/a_466_413# _0565_/a_51_297# 0.00117f
C21512 _0330_ _0356_ 0.01344f
C21513 VPWR _1046_/a_193_47# 0.27357f
C21514 _1022_/a_193_47# _1022_/a_466_413# 0.08301f
C21515 _1022_/a_27_47# _1022_/a_1059_315# 0.04875f
C21516 acc0.A\[31\] _1013_/a_1059_315# 0.02739f
C21517 net44 _0393_ 0.00461f
C21518 _0645_/a_47_47# _0644_/a_47_47# 0.00181f
C21519 _1003_/a_975_413# clknet_1_0__leaf__0460_ 0
C21520 _1021_/a_1059_315# _0462_ 0
C21521 _1052_/a_27_47# _0525_/a_81_21# 0
C21522 _1059_/a_975_413# acc0.A\[15\] 0
C21523 clknet_0__0460_ _0352_ 0.02438f
C21524 _0811_/a_299_297# _0421_ 0.06051f
C21525 _0957_/a_114_297# comp0.B\[6\] 0.00319f
C21526 hold38/a_49_47# clknet_1_1__leaf__0463_ 0.02845f
C21527 _0335_ acc0.A\[30\] 0
C21528 _1008_/a_634_159# net94 0
C21529 _1008_/a_891_413# _1008_/a_1017_47# 0.00617f
C21530 _1055_/a_634_159# _1055_/a_381_47# 0
C21531 _0488_ control0.count\[0\] 0.11328f
C21532 _0279_ VPWR 0.49029f
C21533 hold24/a_49_47# hold24/a_285_47# 0.22264f
C21534 _1020_/a_975_413# _0118_ 0
C21535 _0559_/a_240_47# _0173_ 0.01701f
C21536 clkbuf_0__0461_/a_110_47# _0775_/a_215_47# 0
C21537 _0559_/a_245_297# _0208_ 0
C21538 _0133_ comp0.B\[3\] 0.02851f
C21539 _0771_/a_27_413# _0771_/a_298_297# 0.00498f
C21540 _1054_/a_27_47# net63 0
C21541 hold14/a_49_47# _1036_/a_27_47# 0.01435f
C21542 _1003_/a_193_47# _1003_/a_891_413# 0.19489f
C21543 _1003_/a_27_47# _1003_/a_381_47# 0.06222f
C21544 _1003_/a_634_159# _1003_/a_1059_315# 0
C21545 hold97/a_285_47# _0321_ 0.00251f
C21546 _1055_/a_891_413# net181 0
C21547 _0679_/a_150_297# _0310_ 0
C21548 hold64/a_49_47# _0195_ 0
C21549 _0388_ _0372_ 0
C21550 _0466_ _0974_/a_222_93# 0.00938f
C21551 VPWR _0970_/a_114_47# 0.00198f
C21552 acc0.A\[20\] _0345_ 0
C21553 _0949_/a_59_75# _0467_ 0
C21554 net247 _1048_/a_27_47# 0
C21555 net185 _0955_/a_32_297# 0.09488f
C21556 _0558_/a_68_297# comp0.B\[3\] 0
C21557 hold81/a_285_47# net228 0.00832f
C21558 hold55/a_285_47# _0584_/a_27_297# 0
C21559 net47 acc0.A\[18\] 0.00403f
C21560 clknet_1_0__leaf__0459_ _0208_ 0.04322f
C21561 _0343_ _0238_ 0.54427f
C21562 VPWR _0747_/a_79_21# 0.44507f
C21563 _1054_/a_193_47# net15 0.02796f
C21564 hold67/a_391_47# _0401_ 0
C21565 net29 _0173_ 0
C21566 _1032_/a_592_47# comp0.B\[0\] 0
C21567 _0997_/a_891_413# _0219_ 0
C21568 _0997_/a_592_47# _0345_ 0.00128f
C21569 net235 _0438_ 0
C21570 _0216_ _0779_/a_215_47# 0
C21571 _0855_/a_81_21# net206 0
C21572 _1004_/a_634_159# _0347_ 0
C21573 _0180_ clknet_1_1__leaf__0457_ 0.30799f
C21574 clknet_1_1__leaf__0457_ net218 0.07988f
C21575 hold87/a_391_47# _0181_ 0.05964f
C21576 VPWR _0639_/a_109_297# 0.00652f
C21577 _1054_/a_27_47# _1053_/a_891_413# 0.01154f
C21578 _1054_/a_193_47# _1053_/a_1059_315# 0.00103f
C21579 VPWR hold9/a_49_47# 0.27456f
C21580 _0799_/a_80_21# _0799_/a_209_47# 0.01013f
C21581 _0317_ _0350_ 0
C21582 _0598_/a_382_297# VPWR 0.00453f
C21583 _0773_/a_35_297# _0242_ 0
C21584 VPWR _0987_/a_27_47# 0.61555f
C21585 hold42/a_49_47# net144 0.0056f
C21586 _0270_ _0636_/a_59_75# 0
C21587 _1058_/a_634_159# net189 0.00536f
C21588 net165 _0350_ 0.18582f
C21589 _0557_/a_240_47# _0554_/a_68_297# 0
C21590 _0516_/a_27_297# _0186_ 0.1385f
C21591 net58 _0219_ 0.47268f
C21592 _0951_/a_368_53# _0468_ 0
C21593 _0347_ hold81/a_49_47# 0
C21594 _0464_ clknet_1_0__leaf__0464_ 0.2005f
C21595 _1000_/a_27_47# _0244_ 0.00177f
C21596 _1000_/a_1059_315# _0769_/a_299_297# 0
C21597 pp[30] _0339_ 0.08028f
C21598 VPWR _1029_/a_27_47# 0.77451f
C21599 _0315_ _0360_ 0.02623f
C21600 _0982_/a_634_159# _0452_ 0
C21601 _0982_/a_193_47# _0266_ 0
C21602 _1016_/a_592_47# clknet_1_1__leaf__0461_ 0.00164f
C21603 clknet_1_0__leaf_clk _1064_/a_1059_315# 0
C21604 _1048_/a_27_47# _1048_/a_466_413# 0.27314f
C21605 _1048_/a_193_47# _1048_/a_634_159# 0.11072f
C21606 _1015_/a_1059_315# _0178_ 0
C21607 _0717_/a_303_47# pp[28] 0
C21608 net87 _0218_ 0
C21609 _0106_ hold50/a_391_47# 0
C21610 _0350_ acc0.A\[19\] 0.3589f
C21611 VPWR comp0.B\[9\] 0.59855f
C21612 clknet_1_1__leaf__0460_ _0370_ 0.02988f
C21613 clknet_1_1__leaf__0465_ _0508_/a_81_21# 0.02922f
C21614 _0622_/a_109_47# _0086_ 0
C21615 _0346_ _0434_ 0
C21616 _0555_/a_245_297# VPWR 0.00955f
C21617 _0506_/a_299_297# net229 0.05874f
C21618 _0416_ VPWR 0.51208f
C21619 VPWR _1033_/a_561_413# 0.00213f
C21620 _0387_ _0677_/a_47_47# 0
C21621 net124 _0547_/a_68_297# 0
C21622 net36 _1037_/a_466_413# 0
C21623 _1044_/a_891_413# _0141_ 0
C21624 _0243_ _0245_ 0.05414f
C21625 clknet_1_0__leaf__0465_ _1049_/a_561_413# 0
C21626 hold59/a_49_47# net47 0
C21627 clkbuf_1_1__f__0462_/a_110_47# _0365_ 0
C21628 hold55/a_49_47# VPWR 0.32013f
C21629 hold26/a_49_47# _0473_ 0
C21630 net65 _0434_ 0.01243f
C21631 _0783_/a_215_47# _0218_ 0
C21632 _0101_ _0219_ 0
C21633 _0183_ _0854_/a_79_21# 0
C21634 _0494_/a_27_47# _0213_ 0.00292f
C21635 _0642_/a_27_413# acc0.A\[6\] 0
C21636 _0151_ _1054_/a_634_159# 0
C21637 _0399_ _0186_ 0.55916f
C21638 clkbuf_1_1__f__0463_/a_110_47# _0560_/a_68_297# 0.00128f
C21639 _0349_ _0722_/a_79_21# 0.06784f
C21640 hold57/a_49_47# hold57/a_391_47# 0.00188f
C21641 _1020_/a_27_47# net23 0
C21642 _1010_/a_634_159# _1010_/a_592_47# 0
C21643 clknet_1_0__leaf__0462_ _1004_/a_975_413# 0
C21644 _0276_ acc0.A\[15\] 0.00202f
C21645 _1056_/a_466_413# _0514_/a_27_297# 0
C21646 hold55/a_391_47# _1015_/a_193_47# 0
C21647 hold92/a_391_47# _0345_ 0
C21648 hold6/a_285_47# _0546_/a_51_297# 0.01385f
C21649 _0978_/a_27_297# _0978_/a_109_47# 0.00393f
C21650 _1040_/a_634_159# _1040_/a_381_47# 0
C21651 hold36/a_391_47# net194 0
C21652 _0795_/a_81_21# _0795_/a_384_47# 0.00138f
C21653 _0266_ _0450_ 0.00238f
C21654 _0979_/a_27_297# _0979_/a_373_47# 0.01338f
C21655 _0226_ _0225_ 0
C21656 _0146_ _1048_/a_975_413# 0.00165f
C21657 hold19/a_49_47# _0399_ 0
C21658 _0233_ _0121_ 0
C21659 _0527_/a_27_297# _0527_/a_373_47# 0.01338f
C21660 _0249_ _0350_ 0
C21661 _0216_ _1027_/a_634_159# 0.04504f
C21662 _0195_ _1027_/a_1059_315# 0
C21663 _0751_/a_29_53# _0618_/a_79_21# 0
C21664 _0131_ _0171_ 0
C21665 _1002_/a_592_47# _0217_ 0.00105f
C21666 _1002_/a_1017_47# net150 0
C21667 VPWR _1019_/a_193_47# 0.27883f
C21668 _0532_/a_299_297# clkbuf_1_1__f__0457_/a_110_47# 0
C21669 _0372_ _1006_/a_1059_315# 0
C21670 _0319_ acc0.A\[25\] 0
C21671 net1 _0760_/a_47_47# 0
C21672 _0241_ _0612_/a_59_75# 0
C21673 _0743_/a_51_297# hold90/a_391_47# 0
C21674 clknet_0__0463_ _0562_/a_150_297# 0
C21675 acc0.A\[14\] _0996_/a_466_413# 0.00211f
C21676 _0846_/a_149_47# _0846_/a_240_47# 0.06872f
C21677 _0537_/a_68_297# _1045_/a_27_47# 0
C21678 pp[15] _0411_ 0.00195f
C21679 net45 _1016_/a_381_47# 0
C21680 _1067_/a_634_159# _1067_/a_381_47# 0
C21681 net72 _0345_ 0
C21682 _0174_ net30 0.0024f
C21683 clknet_1_0__leaf__0465_ _0834_/a_109_297# 0
C21684 _1001_/a_193_47# _0345_ 0.0238f
C21685 _1036_/a_27_47# _0208_ 0
C21686 _0458_ net175 0
C21687 _0195_ pp[31] 0.00234f
C21688 _0346_ _0992_/a_1059_315# 0
C21689 _0462_ _0614_/a_111_297# 0
C21690 net123 _0176_ 0
C21691 _0985_/a_193_47# _0529_/a_109_297# 0
C21692 _0985_/a_634_159# _0529_/a_27_297# 0
C21693 _1072_/a_466_413# _1071_/a_891_413# 0.00156f
C21694 _1004_/a_193_47# _0757_/a_68_297# 0
C21695 net65 acc0.A\[7\] 0.35895f
C21696 net9 A[5] 0
C21697 _1009_/a_891_413# _1009_/a_975_413# 0.00851f
C21698 _1009_/a_381_47# _1009_/a_561_413# 0.00123f
C21699 pp[8] net16 0.01664f
C21700 net65 _0989_/a_1059_315# 0.1116f
C21701 acc0.A\[7\] _0989_/a_466_413# 0.00179f
C21702 _0252_ _0989_/a_193_47# 0.47005f
C21703 net235 clknet_1_1__leaf__0465_ 0.00262f
C21704 _0989_/a_193_47# _0989_/a_381_47# 0.09503f
C21705 _0989_/a_634_159# _0989_/a_891_413# 0.03684f
C21706 _0989_/a_27_47# _0989_/a_561_413# 0.0027f
C21707 VPWR _0191_ 0.24451f
C21708 clknet_1_0__leaf__0462_ hold29/a_49_47# 0.0082f
C21709 _0218_ acc0.A\[6\] 0
C21710 _0854_/a_79_21# acc0.A\[15\] 0
C21711 _0544_/a_51_297# _1042_/a_27_47# 0
C21712 _1065_/a_1017_47# control0.reset 0
C21713 _0248_ _0616_/a_78_199# 0.10637f
C21714 _0717_/a_209_297# _0338_ 0.00375f
C21715 _0348_ _0707_/a_544_297# 0.0072f
C21716 _0717_/a_209_47# _0335_ 0
C21717 output58/a_27_47# VPWR 0.44203f
C21718 _0982_/a_1017_47# VPWR 0
C21719 _0476_ _1066_/a_592_47# 0
C21720 _0992_/a_193_47# _0992_/a_381_47# 0.10164f
C21721 _0992_/a_634_159# _0992_/a_891_413# 0.03684f
C21722 _0992_/a_27_47# _0992_/a_561_413# 0.0027f
C21723 _0424_ _0089_ 0.00164f
C21724 _0835_/a_78_199# net62 0
C21725 clkbuf_1_0__f__0457_/a_110_47# _0749_/a_81_21# 0
C21726 _0606_/a_392_297# VPWR 0
C21727 VPWR _1053_/a_381_47# 0.07542f
C21728 _0349_ output55/a_27_47# 0
C21729 _0181_ _0264_ 0.02203f
C21730 _0125_ _1027_/a_891_413# 0.02212f
C21731 acc0.A\[27\] _1027_/a_975_413# 0
C21732 net54 _0739_/a_297_297# 0.00244f
C21733 hold10/a_285_47# control0.reset 0.00123f
C21734 _0354_ _1029_/a_466_413# 0
C21735 net234 _0347_ 0
C21736 _0959_/a_80_21# comp0.B\[6\] 0
C21737 _0959_/a_217_297# comp0.B\[5\] 0
C21738 hold94/a_49_47# hold94/a_285_47# 0.22264f
C21739 _0275_ clkbuf_0__0458_/a_110_47# 0
C21740 _0996_/a_381_47# _0094_ 0.11749f
C21741 _0996_/a_975_413# _0410_ 0
C21742 _0996_/a_592_47# net238 0
C21743 _1045_/a_891_413# _1043_/a_193_47# 0
C21744 _0793_/a_51_297# _0792_/a_80_21# 0
C21745 _0113_ _0208_ 0.514f
C21746 hold75/a_391_47# _0267_ 0.00838f
C21747 _1000_/a_891_413# clknet_0__0461_ 0
C21748 _0262_ _0219_ 0
C21749 hold10/a_49_47# _0465_ 0.00911f
C21750 hold76/a_285_47# _0461_ 0.01198f
C21751 hold10/a_391_47# _1061_/a_1059_315# 0
C21752 _0983_/a_1059_315# net219 0
C21753 _1061_/a_27_47# _1061_/a_466_413# 0.27314f
C21754 _1061_/a_193_47# _1061_/a_634_159# 0.12729f
C21755 _0742_/a_81_21# _0360_ 0
C21756 net62 A[9] 0
C21757 _0659_/a_68_297# _0990_/a_466_413# 0
C21758 net49 VPWR 1.48482f
C21759 _0626_/a_150_297# _0257_ 0
C21760 _0683_/a_113_47# clknet_1_1__leaf__0460_ 0
C21761 hold101/a_49_47# _0837_/a_81_21# 0.0023f
C21762 _0124_ _1026_/a_466_413# 0
C21763 _0572_/a_109_297# net112 0
C21764 _0216_ _1026_/a_891_413# 0.06367f
C21765 _1007_/a_193_47# _0219_ 0.00127f
C21766 _0689_/a_150_297# _0360_ 0
C21767 _0689_/a_68_297# _0321_ 0.13209f
C21768 _0302_ net6 0.06664f
C21769 clkbuf_0__0459_/a_110_47# _0507_/a_109_297# 0
C21770 net22 clkbuf_1_0__f__0463_/a_110_47# 0
C21771 net226 clkbuf_1_0__f_clk/a_110_47# 0.00375f
C21772 clkload0/a_27_47# net35 0.01963f
C21773 _0313_ _0570_/a_109_297# 0
C21774 _1065_/a_27_47# _1063_/a_27_47# 0
C21775 acc0.A\[27\] _0332_ 0
C21776 _0216_ _1024_/a_592_47# 0
C21777 acc0.A\[16\] _0675_/a_68_297# 0.18064f
C21778 _0817_/a_585_47# acc0.A\[9\] 0
C21779 _0817_/a_368_297# _0288_ 0
C21780 _0629_/a_59_75# _0629_/a_145_75# 0.00658f
C21781 _0648_/a_27_297# _0277_ 0.18215f
C21782 clknet_1_1__leaf__0458_ _0826_/a_219_297# 0.01729f
C21783 _0190_ _0988_/a_466_413# 0
C21784 net46 _0104_ 0
C21785 _0804_/a_297_297# _0414_ 0
C21786 clkbuf_0__0459_/a_110_47# hold82/a_49_47# 0
C21787 _1020_/a_561_413# acc0.A\[20\] 0
C21788 hold2/a_391_47# _1047_/a_27_47# 0
C21789 hold2/a_285_47# _1047_/a_193_47# 0
C21790 _0217_ _1014_/a_466_413# 0.03422f
C21791 _0183_ _1014_/a_193_47# 0
C21792 acc0.A\[27\] _0685_/a_68_297# 0.21114f
C21793 _0152_ A[8] 0
C21794 _0195_ net134 0
C21795 _1042_/a_1059_315# net195 0
C21796 _1065_/a_193_47# clknet_1_0__leaf__0457_ 0
C21797 _0182_ _0530_/a_81_21# 0
C21798 _0197_ hold71/a_285_47# 0.00105f
C21799 _0805_/a_27_47# _0993_/a_193_47# 0
C21800 _1033_/a_1017_47# _0215_ 0
C21801 _0984_/a_561_413# acc0.A\[15\] 0
C21802 pp[16] _0219_ 0
C21803 clknet_1_1__leaf__0459_ _0422_ 0.05577f
C21804 _0343_ _0991_/a_466_413# 0.00415f
C21805 _0234_ _0237_ 0.01343f
C21806 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# 1.68035f
C21807 VPWR _1028_/a_891_413# 0.17553f
C21808 _1069_/a_1059_315# _1069_/a_891_413# 0.31086f
C21809 _1069_/a_193_47# _1069_/a_975_413# 0
C21810 _1069_/a_466_413# _1069_/a_381_47# 0.03733f
C21811 hold4/a_391_47# net177 0
C21812 clknet_0__0463_ _0495_/a_68_297# 0.0014f
C21813 VPWR _0812_/a_297_297# 0.00777f
C21814 B[13] net198 0
C21815 _0718_/a_47_47# pp[30] 0.00223f
C21816 _1059_/a_193_47# acc0.A\[13\] 0.00977f
C21817 clknet_0__0465_ _0990_/a_27_47# 0.0027f
C21818 net56 _0336_ 0
C21819 hold69/a_49_47# _0359_ 0
C21820 net10 net195 0
C21821 _0328_ _0219_ 0.09839f
C21822 _0954_/a_32_297# comp0.B\[12\] 0.18249f
C21823 acc0.A\[4\] acc0.A\[3\] 0
C21824 _1037_/a_891_413# comp0.B\[4\] 0
C21825 _0536_/a_240_47# _0172_ 0.03321f
C21826 _1041_/a_634_159# _1040_/a_193_47# 0.00161f
C21827 _1041_/a_193_47# _1040_/a_634_159# 0
C21828 _1041_/a_27_47# _1040_/a_466_413# 0
C21829 _1041_/a_466_413# _1040_/a_27_47# 0
C21830 _1031_/a_466_413# _0220_ 0.02325f
C21831 _0681_/a_113_47# acc0.A\[25\] 0
C21832 hold66/a_285_47# _0369_ 0.04258f
C21833 net213 _0762_/a_79_21# 0.08135f
C21834 _0399_ _1017_/a_193_47# 0
C21835 net48 net49 0.06638f
C21836 hold85/a_285_47# _0466_ 0
C21837 _0219_ _0599_/a_113_47# 0
C21838 _0408_ net5 0
C21839 _1030_/a_466_413# net209 0.00296f
C21840 _0244_ acc0.A\[19\] 0
C21841 VPWR _0512_/a_27_297# 0.24817f
C21842 _1039_/a_27_47# net171 0
C21843 _1018_/a_634_159# clknet_0__0461_ 0
C21844 _0718_/a_285_47# pp[28] 0.00317f
C21845 _0176_ _0544_/a_149_47# 0
C21846 _0346_ _0421_ 0.01183f
C21847 _0624_/a_59_75# _0218_ 0.00988f
C21848 _0241_ _0399_ 0
C21849 _1002_/a_466_413# _0181_ 0.00118f
C21850 _0294_ acc0.A\[18\] 0
C21851 _0480_ _0978_/a_109_297# 0.00206f
C21852 _0415_ _0286_ 0
C21853 _0416_ _0283_ 0.00142f
C21854 _0680_/a_80_21# _0679_/a_68_297# 0
C21855 _0743_/a_240_47# clkbuf_1_0__f__0462_/a_110_47# 0
C21856 _1034_/a_1059_315# _0176_ 0
C21857 acc0.A\[9\] acc0.A\[10\] 0.015f
C21858 _0233_ _0380_ 0
C21859 _0126_ acc0.A\[28\] 0
C21860 hold75/a_49_47# _0446_ 0
C21861 _0231_ _0350_ 0.02867f
C21862 _0538_/a_149_47# _0538_/a_240_47# 0.06872f
C21863 _0538_/a_51_297# _0201_ 0.1051f
C21864 _0462_ net223 0
C21865 _1037_/a_975_413# net26 0
C21866 _0799_/a_80_21# _0668_/a_79_21# 0
C21867 comp0.B\[6\] _0173_ 0.2891f
C21868 _1032_/a_891_413# net201 0
C21869 comp0.B\[3\] _0208_ 0.00569f
C21870 _1022_/a_193_47# net151 0.26134f
C21871 _1022_/a_891_413# _1022_/a_1017_47# 0.00617f
C21872 _0107_ clknet_0__0462_ 0
C21873 clknet_1_1__leaf__0463_ _0565_/a_51_297# 0.00452f
C21874 _1065_/a_193_47# _1062_/a_466_413# 0
C21875 _0822_/a_109_297# _0990_/a_27_47# 0
C21876 clknet_1_0__leaf__0459_ _1019_/a_193_47# 0.03083f
C21877 hold2/a_391_47# clknet_1_0__leaf__0461_ 0.00705f
C21878 _1018_/a_27_47# _0264_ 0
C21879 _0677_/a_285_47# clknet_0__0461_ 0
C21880 net87 _0099_ 0
C21881 net199 _1025_/a_193_47# 0
C21882 _0994_/a_634_159# _0994_/a_381_47# 0
C21883 _1020_/a_1059_315# clknet_1_0__leaf__0457_ 0
C21884 hold12/a_49_47# _0460_ 0.00141f
C21885 VPWR clkbuf_1_0__f__0465_/a_110_47# 1.23349f
C21886 _0284_ net79 0.04586f
C21887 _0275_ _0986_/a_975_413# 0
C21888 net211 _1001_/a_592_47# 0.00164f
C21889 VPWR hold5/a_285_47# 0.33236f
C21890 _0292_ _0422_ 0.00714f
C21891 clkbuf_0__0462_/a_110_47# _0359_ 0.00554f
C21892 _1055_/a_891_413# net179 0.00273f
C21893 _1055_/a_381_47# net141 0
C21894 _0313_ _0361_ 0
C21895 VPWR _0739_/a_79_21# 0.50988f
C21896 hold56/a_391_47# _0564_/a_68_297# 0.01001f
C21897 _1023_/a_193_47# net51 0.04476f
C21898 _0337_ net57 0
C21899 hold22/a_391_47# _1053_/a_27_47# 0
C21900 hold22/a_285_47# _1053_/a_193_47# 0
C21901 _0430_ _0343_ 0.03007f
C21902 _0804_/a_79_21# _0277_ 0
C21903 net226 control0.count\[2\] 0
C21904 net23 hold84/a_391_47# 0
C21905 _1003_/a_466_413# _0101_ 0.03877f
C21906 _1003_/a_1059_315# net89 0
C21907 net36 _1047_/a_891_413# 0.0569f
C21908 _0954_/a_114_297# _0202_ 0.00267f
C21909 _0648_/a_27_297# _0298_ 0.00827f
C21910 _0279_ _0789_/a_75_199# 0
C21911 hold26/a_391_47# _0174_ 0.03008f
C21912 _0426_ _0350_ 0
C21913 net83 net42 0.08309f
C21914 _0248_ _0384_ 0.19261f
C21915 _0533_/a_27_297# net201 0
C21916 _1039_/a_27_47# _1039_/a_466_413# 0.26005f
C21917 _1039_/a_193_47# _1039_/a_634_159# 0.11072f
C21918 _0343_ _0784_/a_113_47# 0
C21919 _0557_/a_51_297# clknet_0__0463_ 0
C21920 hold56/a_391_47# clknet_1_1__leaf_clk 0
C21921 _1020_/a_634_159# _0457_ 0
C21922 net185 _0474_ 0.3208f
C21923 _0343_ _0401_ 0.00117f
C21924 _0501_/a_27_47# _0181_ 0
C21925 net163 net239 0
C21926 _0985_/a_193_47# net170 0.0014f
C21927 _1054_/a_1017_47# _0191_ 0
C21928 acc0.A\[27\] _0738_/a_68_297# 0.00235f
C21929 input4/a_75_212# _0512_/a_27_297# 0
C21930 net36 _0850_/a_68_297# 0
C21931 _0346_ _0809_/a_81_21# 0.05926f
C21932 _0498_/a_51_297# clknet_1_1__leaf__0457_ 0.16379f
C21933 _1010_/a_193_47# _0332_ 0.00117f
C21934 _0172_ _1046_/a_27_47# 0.03825f
C21935 net126 VPWR 0.43373f
C21936 net143 clknet_1_1__leaf__0465_ 0.13714f
C21937 _0844_/a_297_47# _0448_ 0.00107f
C21938 _0729_/a_150_297# clknet_1_1__leaf__0462_ 0
C21939 _0657_/a_109_297# net67 0
C21940 _1004_/a_592_47# _0102_ 0.00164f
C21941 _0987_/a_27_47# _0523_/a_81_21# 0
C21942 _0311_ _0616_/a_215_47# 0
C21943 _1026_/a_27_47# _1026_/a_634_159# 0.14145f
C21944 net157 clkbuf_0__0457_/a_110_47# 0
C21945 net33 _1062_/a_466_413# 0
C21946 VPWR input11/a_75_212# 0.19444f
C21947 _0343_ net222 0
C21948 clknet_0__0458_ hold31/a_391_47# 0
C21949 _0985_/a_27_47# clknet_1_0__leaf__0458_ 0.00143f
C21950 _0983_/a_561_413# _0347_ 0
C21951 _0752_/a_27_413# _1005_/a_891_413# 0
C21952 _0327_ hold90/a_285_47# 0
C21953 net64 _0641_/a_113_47# 0
C21954 net169 _1053_/a_634_159# 0
C21955 net140 _1053_/a_466_413# 0.02345f
C21956 net220 hold73/a_285_47# 0.02667f
C21957 _0982_/a_193_47# _0399_ 0
C21958 _0385_ hold73/a_49_47# 0.12858f
C21959 _0222_ _0618_/a_215_47# 0.07693f
C21960 clknet_1_0__leaf__0465_ net9 0.09343f
C21961 clknet_1_0__leaf__0461_ _0611_/a_68_297# 0.01226f
C21962 clknet_0_clk _0484_ 0
C21963 VPWR input8/a_75_212# 0.27091f
C21964 VPWR _0792_/a_209_47# 0
C21965 clknet_0__0459_ net41 0.02759f
C21966 _1024_/a_193_47# _1024_/a_592_47# 0.00135f
C21967 _1024_/a_466_413# _1024_/a_561_413# 0.00772f
C21968 _1024_/a_634_159# _1024_/a_975_413# 0
C21969 net144 net189 0
C21970 _0217_ _1067_/a_193_47# 0.00225f
C21971 _0355_ _0723_/a_27_413# 0
C21972 _0217_ _0383_ 0
C21973 _0183_ _0369_ 0.49299f
C21974 net205 _0211_ 0
C21975 _0190_ _0186_ 0.02128f
C21976 VPWR _0745_/a_193_47# 0
C21977 _0718_/a_47_47# _0339_ 0.01112f
C21978 clknet_0__0457_ _0183_ 0.08672f
C21979 _1021_/a_891_413# _1020_/a_27_47# 0
C21980 _1011_/a_381_47# _0333_ 0
C21981 _0234_ _0600_/a_253_297# 0
C21982 _0985_/a_381_47# _0182_ 0.00143f
C21983 _0336_ _0345_ 0.00302f
C21984 hold36/a_285_47# _1045_/a_193_47# 0.00207f
C21985 hold36/a_391_47# _1045_/a_27_47# 0
C21986 net33 _0561_/a_149_47# 0
C21987 _0514_/a_109_47# clknet_1_1__leaf__0465_ 0.00312f
C21988 _0369_ output63/a_27_47# 0.00113f
C21989 _0644_/a_129_47# acc0.A\[13\] 0.00282f
C21990 comp0.B\[2\] _1032_/a_891_413# 0
C21991 _0601_/a_68_297# net51 0.15527f
C21992 input3/a_75_212# clknet_1_1__leaf__0465_ 0.00724f
C21993 _0982_/a_1017_47# _0453_ 0
C21994 net68 _0452_ 0
C21995 _0953_/a_32_297# _1040_/a_27_47# 0
C21996 clk _1064_/a_891_413# 0.00407f
C21997 _0949_/a_59_75# net1 0.05848f
C21998 _1048_/a_193_47# net134 0.00664f
C21999 _1048_/a_1059_315# _1048_/a_1017_47# 0
C22000 hold42/a_391_47# A[10] 0
C22001 _0712_/a_465_47# _0220_ 0
C22002 _1034_/a_975_413# clknet_1_1__leaf__0463_ 0
C22003 _0552_/a_68_297# net8 0
C22004 _0399_ _0410_ 0.17617f
C22005 VPWR _0956_/a_220_297# 0.00418f
C22006 _0086_ pp[4] 0
C22007 VPWR _1016_/a_381_47# 0.07235f
C22008 _0731_/a_81_21# _0250_ 0.05947f
C22009 _0607_/a_27_297# _0397_ 0
C22010 _1068_/a_27_47# _0468_ 0.07787f
C22011 _0343_ _1013_/a_27_47# 0.00387f
C22012 _0981_/a_109_297# clkbuf_0_clk/a_110_47# 0
C22013 net167 clknet_1_0__leaf_clk 0.01588f
C22014 _0399_ net62 0.07299f
C22015 _0389_ _0352_ 0.03138f
C22016 _0399_ _0450_ 0
C22017 net36 _0135_ 0
C22018 _0200_ _0545_/a_68_297# 0
C22019 net236 _0958_/a_27_47# 0
C22020 _1060_/a_466_413# _0219_ 0
C22021 net15 acc0.A\[6\] 0.05235f
C22022 _0804_/a_79_21# _0298_ 0
C22023 _0804_/a_297_297# _0404_ 0
C22024 acc0.A\[16\] _0677_/a_47_47# 0.00146f
C22025 _0151_ net140 0
C22026 _0310_ _0678_/a_150_297# 0
C22027 comp0.B\[1\] _1015_/a_1059_315# 0
C22028 _1051_/a_193_47# _0522_/a_27_297# 0
C22029 hold16/a_49_47# _0336_ 0.0367f
C22030 hold16/a_285_47# _0220_ 0.00139f
C22031 clkbuf_1_0__f__0460_/a_110_47# _1006_/a_193_47# 0.00208f
C22032 hold69/a_391_47# net216 0.13119f
C22033 _1056_/a_891_413# net2 0.00308f
C22034 _1056_/a_466_413# _0189_ 0.0022f
C22035 hold69/a_285_47# _0371_ 0.02976f
C22036 hold6/a_391_47# net32 0.00629f
C22037 _0369_ acc0.A\[15\] 0.03701f
C22038 hold26/a_49_47# _0200_ 0.005f
C22039 _1040_/a_891_413# net174 0.04302f
C22040 _1053_/a_1059_315# acc0.A\[6\] 0
C22041 _1053_/a_193_47# net13 0
C22042 clknet_0__0457_ acc0.A\[15\] 0
C22043 clknet_1_0__leaf__0465_ _1054_/a_891_413# 0
C22044 hold79/a_391_47# _0466_ 0.00253f
C22045 _0486_ net91 0
C22046 _0832_/a_113_47# _0350_ 0
C22047 _0979_/a_373_47# _0169_ 0
C22048 net63 _0523_/a_299_297# 0
C22049 _0249_ _1006_/a_634_159# 0
C22050 hold33/a_391_47# comp0.B\[7\] 0
C22051 _0250_ _1006_/a_193_47# 0
C22052 _0216_ _0379_ 0
C22053 _1072_/a_193_47# _1072_/a_592_47# 0.00135f
C22054 _1072_/a_466_413# _1072_/a_561_413# 0.00772f
C22055 _1072_/a_634_159# _1072_/a_975_413# 0
C22056 VPWR _0757_/a_68_297# 0.15429f
C22057 _0751_/a_183_297# _0249_ 0
C22058 _0841_/a_79_21# _0445_ 0.07612f
C22059 net55 clkbuf_0__0462_/a_110_47# 0.00293f
C22060 _0137_ net153 0
C22061 _0216_ _0372_ 0.02798f
C22062 clknet_0__0458_ _0448_ 0
C22063 hold39/a_49_47# clkbuf_1_1__f__0463_/a_110_47# 0
C22064 _0698_/a_113_297# _0321_ 0.00262f
C22065 net101 net149 0
C22066 _0801_/a_113_47# _0347_ 0
C22067 hold26/a_49_47# comp0.B\[8\] 0
C22068 _0640_/a_215_297# _0640_/a_297_297# 0.00659f
C22069 comp0.B\[2\] net106 0
C22070 VPWR _1025_/a_193_47# 0.30838f
C22071 _0772_/a_297_297# _0345_ 0
C22072 _0183_ _0844_/a_79_21# 0
C22073 net161 _0173_ 0
C22074 net187 net118 0
C22075 hold31/a_391_47# net178 0.13549f
C22076 net207 _1015_/a_193_47# 0
C22077 _1019_/a_193_47# _0113_ 0
C22078 _1012_/a_193_47# _0722_/a_79_21# 0
C22079 _0538_/a_240_47# clkbuf_0__0464_/a_110_47# 0
C22080 _0592_/a_68_297# _0374_ 0
C22081 _0730_/a_79_21# _0318_ 0
C22082 VPWR hold95/a_285_47# 0.36064f
C22083 _0476_ _0215_ 0
C22084 _0217_ _1024_/a_634_159# 0
C22085 acc0.A\[8\] _0435_ 0
C22086 _0572_/a_109_297# net111 0
C22087 _1004_/a_891_413# _0380_ 0.00231f
C22088 _0717_/a_209_297# _0348_ 0.00192f
C22089 VPWR net246 0.27959f
C22090 hold75/a_49_47# net61 0
C22091 _0997_/a_466_413# _0997_/a_561_413# 0.00772f
C22092 _0997_/a_634_159# _0997_/a_975_413# 0
C22093 _0640_/a_297_297# _0465_ 0
C22094 _0856_/a_79_21# _0181_ 0
C22095 _1037_/a_27_47# net24 0.00118f
C22096 net71 _0446_ 0
C22097 _0322_ clknet_0__0462_ 0.05856f
C22098 _0880_/a_27_47# hold93/a_49_47# 0
C22099 _0181_ _0986_/a_1017_47# 0
C22100 _0204_ _1042_/a_1059_315# 0.00222f
C22101 net198 _1042_/a_634_159# 0.01811f
C22102 net18 _1042_/a_193_47# 0.03485f
C22103 hold36/a_391_47# net132 0
C22104 _0293_ clknet_0__0465_ 0
C22105 VPWR _1051_/a_975_413# 0.0049f
C22106 _0349_ _1010_/a_634_159# 0.02738f
C22107 _0251_ net58 0
C22108 _0327_ clknet_0__0462_ 0.33984f
C22109 net26 _0173_ 0.30884f
C22110 _0349_ acc0.A\[30\] 0
C22111 hold7/a_285_47# net154 0.01044f
C22112 acc0.A\[12\] _0993_/a_193_47# 0
C22113 net39 _0993_/a_634_159# 0
C22114 VPWR _1045_/a_1017_47# 0
C22115 _0959_/a_80_21# hold84/a_285_47# 0
C22116 _0208_ _0345_ 0.0212f
C22117 _0783_/a_297_297# _0347_ 0.00564f
C22118 clkbuf_1_0__f__0458_/a_110_47# _0084_ 0
C22119 clknet_0__0458_ _0444_ 0.01897f
C22120 net36 _0497_/a_150_297# 0.00123f
C22121 _0268_ _0842_/a_59_75# 0.00159f
C22122 net230 net13 0.02824f
C22123 _0793_/a_245_297# _0408_ 0.0019f
C22124 _1045_/a_1059_315# net129 0
C22125 _0793_/a_240_47# _0400_ 0
C22126 clkbuf_0__0460_/a_110_47# _0691_/a_68_297# 0.01244f
C22127 _0286_ _0347_ 0
C22128 _1027_/a_193_47# _1027_/a_381_47# 0.09799f
C22129 _1027_/a_634_159# _1027_/a_891_413# 0.03684f
C22130 _1027_/a_27_47# _1027_/a_561_413# 0.0027f
C22131 net63 _0172_ 0
C22132 _0179_ _0369_ 0.49351f
C22133 _0741_/a_109_297# _0315_ 0.00178f
C22134 clknet_1_0__leaf__0463_ _0548_/a_245_297# 0
C22135 pp[7] hold65/a_391_47# 0
C22136 _0481_ _0466_ 0.09185f
C22137 _0996_/a_1059_315# net41 0.09303f
C22138 net10 _0204_ 0
C22139 _0465_ _1061_/a_975_413# 0
C22140 _0226_ _0462_ 0.00172f
C22141 _1061_/a_1059_315# _1061_/a_1017_47# 0
C22142 _1061_/a_193_47# net147 0.01358f
C22143 VPWR _1032_/a_466_413# 0.2493f
C22144 net69 net206 0
C22145 comp0.B\[5\] input25/a_75_212# 0
C22146 _0305_ _1009_/a_466_413# 0
C22147 _0460_ acc0.A\[23\] 0
C22148 VPWR _0824_/a_145_75# 0
C22149 _0798_/a_113_297# _0297_ 0
C22150 net66 _0990_/a_592_47# 0
C22151 _0659_/a_68_297# _0088_ 0
C22152 net219 _0612_/a_59_75# 0
C22153 _0581_/a_109_297# acc0.A\[18\] 0.00262f
C22154 _0225_ _0350_ 0.00306f
C22155 _0143_ _0527_/a_373_47# 0
C22156 hold6/a_391_47# net10 0.05252f
C22157 clknet_0__0457_ hold40/a_285_47# 0.02073f
C22158 hold101/a_285_47# _0442_ 0.00828f
C22159 _0197_ _0845_/a_193_297# 0
C22160 net155 acc0.A\[26\] 0.00751f
C22161 _1054_/a_561_413# A[4] 0
C22162 net119 _0955_/a_32_297# 0
C22163 clknet_1_0__leaf__0458_ _0197_ 0
C22164 _0340_ _1030_/a_27_47# 0
C22165 _0844_/a_79_21# acc0.A\[15\] 0.00419f
C22166 _1032_/a_193_47# _1015_/a_891_413# 0
C22167 _0960_/a_27_47# _1071_/a_27_47# 0.00114f
C22168 _1035_/a_1059_315# _1035_/a_891_413# 0.31086f
C22169 _1035_/a_193_47# _1035_/a_975_413# 0
C22170 _1035_/a_466_413# _1035_/a_381_47# 0.03733f
C22171 hold85/a_391_47# net33 0.00113f
C22172 output45/a_27_47# _0111_ 0
C22173 _0280_ _0277_ 0.00308f
C22174 pp[10] _0511_/a_81_21# 0
C22175 _0770_/a_297_47# _0350_ 0.01167f
C22176 _1035_/a_27_47# B[15] 0
C22177 _1053_/a_27_47# A[7] 0.00861f
C22178 _1000_/a_634_159# _0247_ 0.0288f
C22179 net44 _0387_ 0.00711f
C22180 net162 _0338_ 0
C22181 _0412_ _0798_/a_113_297# 0.12969f
C22182 _0559_/a_240_47# net204 0
C22183 _0292_ _0423_ 0.02617f
C22184 init B[4] 0.03078f
C22185 _1013_/a_891_413# clknet_1_1__leaf__0461_ 0
C22186 _1062_/a_27_47# hold93/a_49_47# 0
C22187 _0753_/a_79_21# _0103_ 0
C22188 _0727_/a_109_47# acc0.A\[29\] 0
C22189 net205 _0210_ 0
C22190 _0764_/a_299_297# _0764_/a_384_47# 0
C22191 _0252_ _0988_/a_27_47# 0
C22192 _0343_ _0089_ 0.03213f
C22193 _0569_/a_27_297# net115 0
C22194 acc0.A\[29\] _1029_/a_891_413# 0.01054f
C22195 _1011_/a_193_47# _0726_/a_51_297# 0
C22196 clknet_1_0__leaf__0459_ _1016_/a_381_47# 0
C22197 _1069_/a_561_413# clknet_1_0__leaf_clk 0
C22198 _1069_/a_466_413# control0.count\[0\] 0
C22199 net236 _0481_ 0
C22200 _1069_/a_381_47# _0167_ 0.12224f
C22201 _1033_/a_27_47# _1065_/a_27_47# 0
C22202 _0278_ _0093_ 0
C22203 _0993_/a_27_47# _0650_/a_150_297# 0
C22204 _0993_/a_193_47# _0650_/a_68_297# 0
C22205 _0454_ _0181_ 0.06041f
C22206 _0209_ _0176_ 0.09454f
C22207 net64 _0435_ 0.00103f
C22208 _1052_/a_193_47# _0524_/a_27_297# 0
C22209 _1052_/a_27_47# _0524_/a_109_297# 0
C22210 clknet_1_1__leaf__0460_ _0334_ 0
C22211 input19/a_75_212# clknet_1_1__leaf__0464_ 0
C22212 acc0.A\[31\] output60/a_27_47# 0
C22213 net204 net29 0.00222f
C22214 hold33/a_49_47# hold33/a_391_47# 0.00188f
C22215 _1041_/a_27_47# net174 0
C22216 hold25/a_285_47# clknet_1_0__leaf__0463_ 0.00789f
C22217 net125 _0935_/a_27_47# 0.00313f
C22218 net125 _1061_/a_193_47# 0.03693f
C22219 hold64/a_391_47# _0217_ 0
C22220 hold64/a_49_47# _0183_ 0.01126f
C22221 _0577_/a_109_297# _0217_ 0.0865f
C22222 _0577_/a_109_47# net150 0.00137f
C22223 _0577_/a_27_297# acc0.A\[22\] 0.12312f
C22224 _0953_/a_304_297# _1061_/a_27_47# 0
C22225 _0846_/a_240_47# acc0.A\[15\] 0
C22226 _0211_ net160 0.06041f
C22227 net137 net9 0
C22228 _0750_/a_27_47# _0219_ 0.00144f
C22229 _0778_/a_68_297# _0778_/a_150_297# 0.00477f
C22230 hold69/a_49_47# _0238_ 0.00128f
C22231 _0181_ _0505_/a_27_297# 0.1167f
C22232 _0100_ _0181_ 0.00102f
C22233 _0170_ net35 0
C22234 hold15/a_49_47# hold15/a_285_47# 0.22264f
C22235 _0305_ _0310_ 0.02691f
C22236 _0577_/a_373_47# net151 0
C22237 _0785_/a_81_21# _0291_ 0
C22238 _0173_ hold84/a_285_47# 0
C22239 net106 _1015_/a_193_47# 0
C22240 _0524_/a_27_297# net12 0.18833f
C22241 _0151_ input14/a_75_212# 0.01018f
C22242 _0673_/a_253_297# net228 0
C22243 pp[11] _0993_/a_193_47# 0
C22244 pp[25] _0195_ 0
C22245 net53 _0216_ 0.02692f
C22246 _1065_/a_193_47# _0160_ 0
C22247 _0343_ _0986_/a_891_413# 0
C22248 comp0.B\[11\] _0542_/a_51_297# 0
C22249 input34/a_27_47# rst 0.19704f
C22250 _0575_/a_373_47# acc0.A\[25\] 0
C22251 _0520_/a_27_297# _0520_/a_109_297# 0.17136f
C22252 _0982_/a_634_159# net36 0.03564f
C22253 _0396_ _0097_ 0.0013f
C22254 net45 _1013_/a_634_159# 0.00911f
C22255 hold24/a_49_47# clknet_1_0__leaf__0463_ 0.00888f
C22256 hold26/a_391_47# comp0.B\[9\] 0.05021f
C22257 _0780_/a_35_297# _0240_ 0
C22258 _0236_ _0617_/a_150_297# 0
C22259 _0179_ _1048_/a_634_159# 0.0023f
C22260 _0260_ _0274_ 0.03196f
C22261 _0705_/a_59_75# hold61/a_391_47# 0
C22262 _0463_ control0.sh 0
C22263 _0780_/a_35_297# _0369_ 0
C22264 _1043_/a_27_47# _1042_/a_27_47# 0
C22265 _0255_ _0271_ 0.22691f
C22266 net45 _0607_/a_109_47# 0
C22267 net86 acc0.A\[16\] 0
C22268 _0777_/a_47_47# _0347_ 0.00401f
C22269 _0234_ _0222_ 0.07675f
C22270 _0343_ _0616_/a_78_199# 0
C22271 comp0.B\[4\] net27 0.35939f
C22272 _0280_ _0298_ 0
C22273 _0993_/a_193_47# _0993_/a_592_47# 0.00135f
C22274 _0993_/a_466_413# _0993_/a_561_413# 0.00772f
C22275 _0993_/a_634_159# _0993_/a_975_413# 0
C22276 _0255_ _0987_/a_891_413# 0.00185f
C22277 _0279_ _0345_ 0
C22278 _0816_/a_68_297# acc0.A\[9\] 0.07578f
C22279 _0181_ _0506_/a_81_21# 0.00839f
C22280 net102 net206 0
C22281 clknet_0__0463_ net7 0.00296f
C22282 net49 _1023_/a_27_47# 0
C22283 hold18/a_391_47# net165 0.13584f
C22284 _1039_/a_193_47# net125 0.01327f
C22285 _1039_/a_1059_315# _1039_/a_1017_47# 0
C22286 output64/a_27_47# acc0.A\[6\] 0.02475f
C22287 hold31/a_49_47# _0274_ 0.02912f
C22288 acc0.A\[1\] net175 0
C22289 _0218_ _0611_/a_68_297# 0.01323f
C22290 _1039_/a_466_413# _0953_/a_32_297# 0
C22291 _0973_/a_27_297# clknet_1_0__leaf__0460_ 0.01652f
C22292 _0713_/a_27_47# _0352_ 0
C22293 _0280_ _0296_ 0.55154f
C22294 _0580_/a_27_297# _0580_/a_109_47# 0.00393f
C22295 _0663_/a_297_47# _0293_ 0
C22296 _0673_/a_103_199# _0347_ 0.06448f
C22297 _0672_/a_79_21# _0347_ 0
C22298 _0399_ net219 0
C22299 _0179_ _0846_/a_240_47# 0.03313f
C22300 clknet_1_0__leaf__0463_ _1048_/a_193_47# 0
C22301 _0465_ _0261_ 0.01476f
C22302 net135 _0528_/a_384_47# 0
C22303 _0190_ net62 0
C22304 _1059_/a_193_47# VPWR 0.3058f
C22305 _1026_/a_891_413# _1026_/a_975_413# 0.00851f
C22306 _1026_/a_27_47# net112 0.23672f
C22307 _1026_/a_381_47# _1026_/a_561_413# 0.00123f
C22308 net33 _0160_ 0.07162f
C22309 _0361_ _0321_ 0
C22310 _0985_/a_634_159# _0449_ 0
C22311 clknet_1_0__leaf__0461_ hold93/a_391_47# 0.00507f
C22312 A[10] net16 0.00122f
C22313 _0361_ clkbuf_0__0460_/a_110_47# 0.00132f
C22314 _0187_ net37 0.02821f
C22315 net36 _0206_ 0
C22316 _0697_/a_217_297# _0324_ 0.04994f
C22317 net141 clknet_1_1__leaf__0458_ 0.00206f
C22318 _0172_ hold5/a_49_47# 0
C22319 net169 net139 0
C22320 net58 _0262_ 0.1301f
C22321 acc0.A\[2\] _0261_ 0.18442f
C22322 _0720_/a_68_297# net239 0.10522f
C22323 _0718_/a_377_297# _0348_ 0.00284f
C22324 _0181_ _1009_/a_466_413# 0.00363f
C22325 net192 _0186_ 0
C22326 _0195_ net165 0
C22327 _0466_ _0477_ 0
C22328 _0695_/a_472_297# _0324_ 0.00412f
C22329 _1024_/a_1059_315# acc0.A\[24\] 0.0855f
C22330 _0542_/a_51_297# _0202_ 0
C22331 net61 net71 0
C22332 _0454_ _1018_/a_27_47# 0
C22333 net227 acc0.A\[28\] 0
C22334 _0639_/a_109_297# _0345_ 0
C22335 hold30/a_49_47# net50 0
C22336 hold36/a_285_47# _1044_/a_27_47# 0.00127f
C22337 hold9/a_49_47# _0345_ 0
C22338 clk _0471_ 0.02394f
C22339 hold66/a_285_47# hold66/a_391_47# 0.41909f
C22340 _0284_ _0301_ 0
C22341 _0527_/a_109_297# _0186_ 0.02774f
C22342 _0230_ _0754_/a_51_297# 0.04496f
C22343 net57 _0333_ 0.0318f
C22344 net24 _0561_/a_51_297# 0
C22345 _0375_ _0232_ 0
C22346 _0662_/a_81_21# _0662_/a_384_47# 0.00138f
C22347 _0346_ _0186_ 0
C22348 _0343_ _0854_/a_215_47# 0
C22349 _0251_ net168 0
C22350 _1057_/a_381_47# net143 0
C22351 hold36/a_49_47# net131 0
C22352 _0174_ _1040_/a_27_47# 0.02898f
C22353 _1037_/a_27_47# _1037_/a_466_413# 0.27314f
C22354 _1037_/a_193_47# _1037_/a_634_159# 0.11072f
C22355 control0.state\[0\] _0978_/a_27_297# 0
C22356 pp[16] _0997_/a_891_413# 0
C22357 _0463_ net157 0
C22358 _0182_ _0147_ 0
C22359 _0180_ net135 0
C22360 _0402_ _0992_/a_27_47# 0
C22361 hold4/a_49_47# hold4/a_391_47# 0.00188f
C22362 _0627_/a_215_53# _0445_ 0
C22363 _0202_ _0142_ 0
C22364 comp0.B\[10\] _1040_/a_634_159# 0
C22365 _0972_/a_250_297# _0951_/a_109_93# 0
C22366 net65 _0186_ 0.18325f
C22367 hold48/a_285_47# net20 0
C22368 _1029_/a_27_47# _0345_ 0
C22369 _0785_/a_81_21# _0290_ 0
C22370 _0785_/a_299_297# _0423_ 0
C22371 _0253_ _0434_ 0.44938f
C22372 hold48/a_49_47# hold48/a_391_47# 0.00188f
C22373 _0195_ acc0.A\[19\] 0.04177f
C22374 net126 net30 0
C22375 _0305_ _0768_/a_27_47# 0
C22376 _0352_ net50 0.00249f
C22377 _1041_/a_1059_315# _1041_/a_891_413# 0.31086f
C22378 _1041_/a_193_47# _1041_/a_975_413# 0
C22379 _1041_/a_466_413# _1041_/a_381_47# 0.03733f
C22380 _1048_/a_891_413# clknet_1_1__leaf__0457_ 0
C22381 _0133_ net24 0
C22382 VPWR _0991_/a_891_413# 0.23341f
C22383 net87 _0721_/a_27_47# 0.00125f
C22384 _0157_ _0661_/a_205_297# 0
C22385 _0465_ _0509_/a_27_47# 0
C22386 _1054_/a_27_47# _0180_ 0.03442f
C22387 clknet_1_1__leaf__0463_ clkbuf_1_1__f_clk/a_110_47# 0
C22388 _0243_ _0769_/a_81_21# 0.0735f
C22389 control0.reset clknet_1_0__leaf__0461_ 0
C22390 clknet_1_0__leaf__0460_ net17 0
C22391 _1015_/a_1017_47# comp0.B\[15\] 0
C22392 _0158_ _0219_ 0.01757f
C22393 output56/a_27_47# _1030_/a_27_47# 0
C22394 _0416_ _0345_ 0.00225f
C22395 hold42/a_49_47# A[11] 0
C22396 _0176_ _1043_/a_466_413# 0
C22397 _0409_ acc0.A\[15\] 0
C22398 acc0.A\[2\] _0509_/a_27_47# 0.04508f
C22399 A[5] A[7] 0.1786f
C22400 _0399_ _0637_/a_56_297# 0
C22401 _1039_/a_193_47# _0473_ 0.02402f
C22402 _0569_/a_109_297# acc0.A\[28\] 0.00776f
C22403 _0275_ _0447_ 0
C22404 clkbuf_0__0464_/a_110_47# net147 0
C22405 _0852_/a_35_297# net165 0
C22406 _1051_/a_193_47# _0193_ 0
C22407 hold86/a_49_47# _0219_ 0.05115f
C22408 _0247_ _0242_ 0.09035f
C22409 _0305_ _0184_ 0
C22410 _0399_ _0812_/a_510_47# 0
C22411 _0532_/a_81_21# _0531_/a_27_297# 0
C22412 _0305_ _0239_ 0
C22413 _1057_/a_27_47# net3 0
C22414 clkbuf_1_0__f__0457_/a_110_47# _0242_ 0
C22415 _0310_ _0181_ 0.02285f
C22416 hold97/a_285_47# _0738_/a_68_297# 0
C22417 net232 hold84/a_285_47# 0.00325f
C22418 VPWR _1011_/a_193_47# 0.30717f
C22419 _0752_/a_27_413# _0369_ 0
C22420 _0234_ _0762_/a_297_297# 0.00464f
C22421 _0251_ _0831_/a_285_297# 0.00158f
C22422 _0249_ net92 0
C22423 net53 _1024_/a_193_47# 0
C22424 net123 net28 0
C22425 _0476_ _0955_/a_304_297# 0
C22426 pp[2] _0827_/a_109_297# 0
C22427 hold70/a_49_47# hold81/a_285_47# 0
C22428 _0297_ net41 0
C22429 _0465_ net47 0.00273f
C22430 _0229_ _0228_ 0.1134f
C22431 net160 _0210_ 0.21702f
C22432 _0118_ _0586_/a_27_47# 0
C22433 _0358_ clknet_1_1__leaf__0462_ 0
C22434 _0081_ net165 0
C22435 _0609_/a_109_297# _0461_ 0
C22436 _1019_/a_193_47# _0345_ 0.06781f
C22437 _0985_/a_193_47# _0846_/a_51_297# 0
C22438 _0361_ _1009_/a_27_47# 0.0013f
C22439 _0574_/a_109_297# net50 0
C22440 hold69/a_391_47# _0370_ 0.00108f
C22441 _0182_ _0584_/a_373_47# 0
C22442 _1012_/a_1059_315# _0351_ 0
C22443 _1012_/a_634_159# _0110_ 0.00379f
C22444 net21 clknet_0__0464_ 0.00653f
C22445 _0713_/a_27_47# net207 0
C22446 _0343_ _0384_ 0
C22447 clknet_1_1__leaf__0459_ _0276_ 0.07886f
C22448 hold27/a_391_47# _0172_ 0.05379f
C22449 _0217_ net110 0.32036f
C22450 _0225_ _1005_/a_1059_315# 0
C22451 _0412_ net41 0
C22452 _1051_/a_27_47# _0150_ 0
C22453 _0195_ net197 0.27584f
C22454 _0578_/a_109_297# VPWR 0.19316f
C22455 _0644_/a_129_47# VPWR 0
C22456 net239 net116 0.00668f
C22457 acc0.A\[21\] clknet_1_0__leaf__0460_ 0.38144f
C22458 acc0.A\[27\] clknet_0__0460_ 0.03273f
C22459 _0583_/a_27_297# net6 0
C22460 _0140_ _1042_/a_592_47# 0
C22461 VPWR _1044_/a_592_47# 0
C22462 _0146_ _1049_/a_193_47# 0
C22463 clknet_1_0__leaf__0462_ _0228_ 0
C22464 net125 clkbuf_0__0464_/a_110_47# 0
C22465 acc0.A\[14\] _0219_ 0.43157f
C22466 _0161_ hold84/a_391_47# 0
C22467 _0313_ VPWR 1.84689f
C22468 _0349_ net96 0
C22469 _0316_ _0697_/a_217_297# 0
C22470 hold35/a_285_47# _0189_ 0.00477f
C22471 _0217_ clkbuf_1_1__f__0457_/a_110_47# 0.00315f
C22472 _0399_ _0352_ 0.05462f
C22473 _0661_/a_27_297# _0288_ 0.17538f
C22474 _0982_/a_1017_47# _0345_ 0
C22475 _0756_/a_377_297# _0379_ 0.00206f
C22476 net55 _0331_ 0
C22477 _1001_/a_592_47# _0461_ 0
C22478 clkbuf_1_1__f__0465_/a_110_47# _0422_ 0.00441f
C22479 _1027_/a_1059_315# net156 0
C22480 _0643_/a_103_199# _0274_ 0.11811f
C22481 _0643_/a_253_297# _0272_ 0
C22482 net44 _0340_ 0.00338f
C22483 _0606_/a_392_297# _0345_ 0
C22484 _0606_/a_215_297# net241 0
C22485 clknet_1_1__leaf__0460_ _0240_ 0
C22486 _0697_/a_80_21# _0739_/a_79_21# 0
C22487 net179 net47 0
C22488 net1 _1014_/a_27_47# 0.00215f
C22489 _1030_/a_1059_315# _0707_/a_75_199# 0
C22490 _1030_/a_466_413# _0707_/a_201_297# 0
C22491 net239 hold92/a_285_47# 0.00983f
C22492 clknet_1_1__leaf__0460_ _0369_ 0.0014f
C22493 VPWR net202 0.25302f
C22494 _0293_ _0986_/a_27_47# 0
C22495 comp0.B\[2\] _0560_/a_150_297# 0
C22496 _0747_/a_79_21# net52 0.01829f
C22497 _0749_/a_81_21# _0248_ 0.06164f
C22498 _0710_/a_381_47# VPWR 0
C22499 hold22/a_49_47# acc0.A\[8\] 0
C22500 output66/a_27_47# pp[8] 0.38099f
C22501 _0636_/a_59_75# net170 0
C22502 clknet_1_0__leaf__0462_ _1023_/a_561_413# 0
C22503 clknet_0__0465_ _0840_/a_150_297# 0
C22504 net204 comp0.B\[6\] 0
C22505 _0482_ _0488_ 0.03876f
C22506 VPWR clknet_1_1__leaf__0463_ 3.95279f
C22507 clknet_0__0460_ _0364_ 0
C22508 _0582_/a_27_297# _0582_/a_109_47# 0.00393f
C22509 _0751_/a_183_297# _0225_ 0.00407f
C22510 net119 _0474_ 0.00183f
C22511 net202 _1015_/a_466_413# 0.00291f
C22512 acc0.A\[20\] clknet_1_0__leaf__0457_ 0.06295f
C22513 _0478_ _1071_/a_634_159# 0
C22514 _1007_/a_27_47# _1007_/a_634_159# 0.14145f
C22515 _1052_/a_27_47# _1052_/a_1059_315# 0.04875f
C22516 _1052_/a_193_47# _1052_/a_466_413# 0.07482f
C22517 _0991_/a_975_413# clknet_1_1__leaf__0465_ 0
C22518 _1035_/a_381_47# _0133_ 0.13142f
C22519 clknet_1_0__leaf__0465_ _0255_ 0.5678f
C22520 hold87/a_285_47# _0266_ 0.0019f
C22521 _0348_ net162 0
C22522 _1012_/a_193_47# acc0.A\[30\] 0
C22523 _0358_ net242 0
C22524 net186 _1034_/a_27_47# 0.07128f
C22525 _1058_/a_193_47# _1058_/a_891_413# 0.19489f
C22526 _1058_/a_27_47# _1058_/a_381_47# 0.06222f
C22527 _1058_/a_634_159# _1058_/a_1059_315# 0
C22528 clkload4/a_268_47# _0459_ 0
C22529 clknet_1_0__leaf__0464_ hold7/a_49_47# 0
C22530 _0343_ _0781_/a_150_297# 0
C22531 net86 _0247_ 0.01048f
C22532 hold14/a_49_47# net24 0
C22533 hold14/a_285_47# B[1] 0.00153f
C22534 clk _0977_/a_75_212# 0.00124f
C22535 _0353_ _0723_/a_207_413# 0.07587f
C22536 _0172_ _1045_/a_592_47# 0.00112f
C22537 VPWR net8 0.5836f
C22538 net69 _0849_/a_215_47# 0
C22539 net185 _1035_/a_27_47# 0
C22540 hold41/a_285_47# acc0.A\[12\] 0
C22541 net134 acc0.A\[15\] 0
C22542 _1050_/a_466_413# _0527_/a_27_297# 0
C22543 _1050_/a_634_159# _0527_/a_109_297# 0
C22544 _1010_/a_1059_315# _0333_ 0
C22545 VPWR net32 0.97923f
C22546 _0718_/a_129_47# _0349_ 0
C22547 _0343_ pp[28] 0.3777f
C22548 net44 acc0.A\[16\] 0.0191f
C22549 _0462_ _0773_/a_285_297# 0
C22550 _1011_/a_466_413# _0355_ 0.00645f
C22551 _1011_/a_634_159# net227 0
C22552 VPWR _1013_/a_634_159# 0.17799f
C22553 _0167_ control0.count\[0\] 0
C22554 _1002_/a_27_47# VPWR 0.6324f
C22555 _0182_ _1015_/a_891_413# 0
C22556 _1052_/a_466_413# net12 0.00298f
C22557 _1052_/a_193_47# _0194_ 0
C22558 _0642_/a_382_47# _0434_ 0
C22559 _0831_/a_35_297# clknet_1_1__leaf__0458_ 0.0046f
C22560 _0328_ _1007_/a_193_47# 0
C22561 clkbuf_1_1__f__0460_/a_110_47# _0319_ 0
C22562 _0812_/a_297_297# _0345_ 0
C22563 _0174_ _1061_/a_466_413# 0
C22564 net149 hold60/a_285_47# 0
C22565 _0607_/a_27_297# clkbuf_0__0461_/a_110_47# 0
C22566 clkbuf_0__0464_/a_110_47# _0473_ 0.01285f
C22567 acc0.A\[22\] _0120_ 0.41362f
C22568 comp0.B\[10\] _1061_/a_891_413# 0
C22569 _0195_ _1018_/a_975_413# 0
C22570 _1027_/a_1059_315# acc0.A\[26\] 0
C22571 hold68/a_285_47# _0380_ 0
C22572 _0174_ net171 0.44161f
C22573 net58 _0988_/a_975_413# 0
C22574 _0300_ _0405_ 0.01901f
C22575 net208 net209 0.02185f
C22576 _0786_/a_80_21# _0786_/a_472_297# 0.01636f
C22577 _0181_ _0184_ 0.00967f
C22578 _0855_/a_81_21# hold18/a_49_47# 0
C22579 acc0.A\[31\] net162 0
C22580 _0462_ _0350_ 0.0982f
C22581 _0239_ _0181_ 0
C22582 _1038_/a_891_413# _0176_ 0.00573f
C22583 _0575_/a_27_297# _0216_ 0.17601f
C22584 _0461_ _0294_ 0.00794f
C22585 _1021_/a_193_47# acc0.A\[20\] 0
C22586 _0974_/a_79_199# _0974_/a_222_93# 0.22112f
C22587 _0530_/a_81_21# _1048_/a_1059_315# 0.01733f
C22588 _1039_/a_27_47# _0497_/a_150_297# 0
C22589 net205 _1034_/a_634_159# 0
C22590 hold11/a_49_47# _1049_/a_27_47# 0
C22591 clknet_1_0__leaf__0462_ _0323_ 0
C22592 _0984_/a_27_47# VPWR 0.71113f
C22593 _0985_/a_634_159# _0260_ 0
C22594 net12 _0194_ 0.26309f
C22595 _0880_/a_27_47# clknet_1_0__leaf__0457_ 0.19969f
C22596 net9 _0148_ 0.03823f
C22597 _0994_/a_634_159# _0218_ 0.00552f
C22598 _0550_/a_51_297# net152 0
C22599 net59 _1012_/a_891_413# 0.00429f
C22600 _0195_ net1 0.05049f
C22601 _1010_/a_27_47# net98 0
C22602 acc0.A\[30\] clknet_1_1__leaf__0461_ 0
C22603 hold75/a_49_47# _0269_ 0
C22604 comp0.B\[12\] net19 0.00714f
C22605 _0869_/a_27_47# clknet_1_0__leaf__0461_ 0.00399f
C22606 net89 net159 0.00504f
C22607 hold13/a_391_47# _1039_/a_27_47# 0
C22608 net111 _1026_/a_27_47# 0.00866f
C22609 _0995_/a_891_413# pp[14] 0.02479f
C22610 _0413_ _0400_ 0
C22611 _0520_/a_27_297# _0186_ 0.08933f
C22612 clknet_1_0__leaf__0465_ A[7] 0.2645f
C22613 _0520_/a_373_47# net14 0.00164f
C22614 _0798_/a_199_47# _0219_ 0
C22615 net68 net36 0.23709f
C22616 _1002_/a_27_47# net48 0
C22617 VPWR _1042_/a_1059_315# 0.40683f
C22618 _1056_/a_634_159# acc0.A\[9\] 0.00145f
C22619 _0982_/a_193_47# _0346_ 0.02622f
C22620 _0195_ clkbuf_1_1__f__0461_/a_110_47# 0
C22621 _1028_/a_466_413# _1008_/a_27_47# 0
C22622 _0179_ net134 0.04353f
C22623 _0518_/a_109_47# net65 0
C22624 _0201_ comp0.B\[10\] 0
C22625 pp[26] _0572_/a_27_297# 0
C22626 _1043_/a_381_47# _1042_/a_891_413# 0
C22627 _1043_/a_891_413# _1042_/a_381_47# 0
C22628 clknet_1_1__leaf__0464_ net18 0.02078f
C22629 _1030_/a_193_47# acc0.A\[30\] 0.05642f
C22630 _0642_/a_215_297# _0252_ 0.15345f
C22631 net207 _0399_ 0.05041f
C22632 _0328_ _0599_/a_113_47# 0
C22633 _0857_/a_27_47# clknet_1_0__leaf__0457_ 0.00422f
C22634 hold89/a_285_47# _0488_ 0.00111f
C22635 hold89/a_49_47# _0466_ 0.03129f
C22636 _0233_ _0369_ 0
C22637 pp[27] _1030_/a_561_413# 0
C22638 _0988_/a_634_159# _0988_/a_466_413# 0.23992f
C22639 _0988_/a_193_47# _0988_/a_1059_315# 0.03405f
C22640 _0988_/a_27_47# _0988_/a_891_413# 0.03224f
C22641 _1039_/a_466_413# _0174_ 0
C22642 _0984_/a_891_413# _0983_/a_193_47# 0
C22643 _0368_ _0366_ 0.06688f
C22644 VPWR net10 3.12424f
C22645 net43 _0097_ 0.00215f
C22646 _0730_/a_297_297# _0358_ 0
C22647 _0730_/a_215_47# _0357_ 0.05635f
C22648 clknet_1_1__leaf__0460_ _1010_/a_381_47# 0.00704f
C22649 _0165_ clknet_1_0__leaf__0460_ 0.05728f
C22650 net63 _0836_/a_150_297# 0.00134f
C22651 _0216_ net60 0
C22652 _0953_/a_32_297# _0953_/a_304_297# 0.00167f
C22653 hold20/a_391_47# net167 0.13057f
C22654 hold28/a_285_47# _0465_ 0
C22655 _0478_ _0978_/a_27_297# 0.01145f
C22656 _0312_ _0694_/a_113_47# 0
C22657 _0695_/a_80_21# _0326_ 0.08596f
C22658 _0542_/a_245_297# _0542_/a_240_47# 0
C22659 _0346_ _0410_ 0.03751f
C22660 net63 _0437_ 0.24479f
C22661 hold96/a_391_47# _0575_/a_27_297# 0.00545f
C22662 hold96/a_285_47# _0575_/a_109_297# 0.00207f
C22663 _0485_ _1064_/a_592_47# 0
C22664 _0162_ _1064_/a_381_47# 0.12138f
C22665 clkbuf_1_0__f__0463_/a_110_47# control0.sh 0
C22666 net216 _0219_ 0.00173f
C22667 net171 _0208_ 0.02497f
C22668 _0982_/a_193_47# _0629_/a_59_75# 0
C22669 _1001_/a_193_47# clknet_1_0__leaf__0457_ 0.04545f
C22670 acc0.A\[2\] hold28/a_285_47# 0.00618f
C22671 _0465_ _1047_/a_1017_47# 0
C22672 _0225_ _0592_/a_68_297# 0.05504f
C22673 _0999_/a_27_47# _0097_ 0.13799f
C22674 _0346_ net62 0.0314f
C22675 _0089_ _0842_/a_59_75# 0
C22676 _0999_/a_634_159# _0396_ 0
C22677 _1003_/a_193_47# net240 0
C22678 clknet_1_0__leaf__0457_ _1062_/a_27_47# 0
C22679 _0472_ _1061_/a_1017_47# 0
C22680 _0346_ _0450_ 0
C22681 _0817_/a_368_297# _0424_ 0.0025f
C22682 clknet_1_1__leaf__0460_ _1009_/a_561_413# 0
C22683 net56 hold95/a_285_47# 0.08481f
C22684 _1035_/a_193_47# net27 0.03722f
C22685 clknet_1_0__leaf__0459_ net202 0
C22686 output67/a_27_47# output37/a_27_47# 0.0033f
C22687 clkbuf_1_1__f__0459_/a_110_47# hold91/a_49_47# 0
C22688 _0853_/a_150_297# _0218_ 0
C22689 _0981_/a_373_47# _0484_ 0
C22690 net46 _0616_/a_292_297# 0
C22691 _0452_ _0264_ 0.02818f
C22692 _0982_/a_466_413# hold60/a_285_47# 0
C22693 comp0.B\[9\] _1040_/a_27_47# 0
C22694 hold48/a_49_47# net195 0
C22695 _0787_/a_209_297# _0787_/a_303_47# 0
C22696 _0279_ _0994_/a_27_47# 0
C22697 _0795_/a_81_21# acc0.A\[13\] 0
C22698 net24 _0208_ 0.27813f
C22699 _0230_ _0219_ 0.08548f
C22700 _0404_ _0405_ 0.28144f
C22701 _0792_/a_209_47# _0345_ 0.00176f
C22702 _0315_ _0181_ 0
C22703 clkload2/Y VPWR 0.44772f
C22704 _0399_ _0849_/a_79_21# 0.12786f
C22705 _1037_/a_27_47# _0135_ 0.09849f
C22706 _1037_/a_1059_315# _1037_/a_1017_47# 0
C22707 _0997_/a_466_413# _0218_ 0
C22708 VPWR hold70/a_391_47# 0.1689f
C22709 _0195_ _0998_/a_1059_315# 0.04577f
C22710 _0305_ _0309_ 0.03517f
C22711 _0502_/a_27_47# comp0.B\[15\] 0.00545f
C22712 net231 _0951_/a_209_311# 0.08694f
C22713 _0465_ _0848_/a_109_297# 0
C22714 pp[30] _1030_/a_466_413# 0.00686f
C22715 clknet_1_0__leaf__0462_ net237 0.0015f
C22716 _0779_/a_79_21# clknet_1_1__leaf__0461_ 0
C22717 _0608_/a_27_47# _0397_ 0
C22718 net44 output56/a_27_47# 0
C22719 VPWR _1005_/a_592_47# 0.00317f
C22720 net42 _0406_ 0.03835f
C22721 _0690_/a_68_297# _0318_ 0.16904f
C22722 _0310_ clknet_1_1__leaf__0461_ 0
C22723 hold89/a_285_47# _1064_/a_27_47# 0
C22724 _0985_/a_27_47# _0448_ 0
C22725 _0121_ _1023_/a_1059_315# 0
C22726 net204 net26 0
C22727 _1001_/a_27_47# _1001_/a_891_413# 0.03224f
C22728 _1001_/a_193_47# _1001_/a_1059_315# 0.03225f
C22729 _1001_/a_634_159# _1001_/a_466_413# 0.23992f
C22730 _0430_ acc0.A\[6\] 0.70313f
C22731 net150 _0181_ 0
C22732 _0621_/a_285_47# acc0.A\[6\] 0.0025f
C22733 _0440_ net148 0
C22734 _0343_ _0825_/a_150_297# 0
C22735 _0607_/a_109_47# clknet_1_0__leaf__0459_ 0
C22736 control0.add hold73/a_49_47# 0
C22737 VPWR _0232_ 0.27725f
C22738 hold76/a_285_47# net223 0.01031f
C22739 hold76/a_49_47# _0391_ 0
C22740 _0176_ net196 0.09954f
C22741 net189 A[11] 0
C22742 _0553_/a_240_47# _0957_/a_32_297# 0
C22743 _1062_/a_27_47# _1062_/a_466_413# 0.27314f
C22744 _1062_/a_193_47# _1062_/a_634_159# 0.12603f
C22745 _0708_/a_68_297# output60/a_27_47# 0
C22746 _0239_ _0677_/a_377_297# 0
C22747 _0183_ hold40/a_391_47# 0.00141f
C22748 _0341_ _0567_/a_27_297# 0.0071f
C22749 _0254_ net47 0
C22750 _0217_ _0486_ 0
C22751 hold38/a_391_47# _0951_/a_109_93# 0
C22752 hold38/a_285_47# _0951_/a_209_311# 0
C22753 acc0.A\[5\] acc0.A\[6\] 0
C22754 _0149_ net13 0
C22755 output55/a_27_47# _0354_ 0
C22756 hold90/a_49_47# hold90/a_285_47# 0.22264f
C22757 _0575_/a_109_297# _1024_/a_27_47# 0
C22758 _0575_/a_27_297# _1024_/a_193_47# 0.00116f
C22759 clkbuf_1_1__f__0465_/a_110_47# _0423_ 0
C22760 _0198_ net175 0.18544f
C22761 _1049_/a_891_413# _1048_/a_634_159# 0.0021f
C22762 _1049_/a_1059_315# _1048_/a_466_413# 0.0028f
C22763 _0227_ hold94/a_49_47# 0.04404f
C22764 hold14/a_391_47# _1037_/a_193_47# 0
C22765 hold14/a_49_47# _1037_/a_466_413# 0
C22766 _0376_ _0383_ 0.00259f
C22767 _0572_/a_109_297# VPWR 0.1958f
C22768 VPWR _1006_/a_561_413# 0.003f
C22769 _0459_ _1060_/a_27_47# 0
C22770 _0222_ hold29/a_391_47# 0
C22771 _0285_ _0787_/a_80_21# 0.0579f
C22772 _1000_/a_634_159# _0217_ 0
C22773 _1000_/a_27_47# _0183_ 0
C22774 hold43/a_285_47# _1029_/a_27_47# 0
C22775 _0343_ net229 0
C22776 _0481_ _1069_/a_1059_315# 0.00137f
C22777 _0963_/a_35_297# clknet_1_0__leaf_clk 0.04231f
C22778 net194 _0538_/a_240_47# 0
C22779 _0195_ _1030_/a_592_47# 0.00307f
C22780 _0216_ _1030_/a_561_413# 0
C22781 net48 _1005_/a_592_47# 0
C22782 VPWR _0986_/a_561_413# 0.00296f
C22783 _1039_/a_193_47# comp0.B\[8\] 0
C22784 hold52/a_391_47# _0347_ 0
C22785 net101 comp0.B\[15\] 0
C22786 _0714_/a_149_47# _0219_ 0.00356f
C22787 pp[9] _1058_/a_891_413# 0
C22788 _0663_/a_27_413# _0399_ 0
C22789 _0343_ _0797_/a_27_413# 0.0015f
C22790 _1070_/a_193_47# _0978_/a_27_297# 0
C22791 _0185_ _0505_/a_373_47# 0
C22792 _1031_/a_193_47# net209 0
C22793 hold26/a_285_47# _0546_/a_51_297# 0
C22794 _0244_ _0462_ 0.00158f
C22795 _1004_/a_1059_315# _0216_ 0
C22796 _0460_ clknet_1_0__leaf__0461_ 0.00553f
C22797 clknet_1_0__leaf__0457_ net107 0.00879f
C22798 hold66/a_285_47# _0374_ 0
C22799 hold78/a_391_47# _0714_/a_51_297# 0.00864f
C22800 clknet_1_1__leaf__0459_ _0369_ 0.02454f
C22801 _0554_/a_68_297# _0552_/a_68_297# 0
C22802 acc0.A\[5\] _0523_/a_384_47# 0
C22803 _0561_/a_51_297# _0561_/a_149_47# 0.02487f
C22804 VPWR _0616_/a_493_297# 0.00297f
C22805 _1072_/a_193_47# _1068_/a_1059_315# 0
C22806 _1072_/a_27_47# _1068_/a_891_413# 0
C22807 _0476_ _1065_/a_193_47# 0
C22808 _0251_ _0833_/a_79_21# 0
C22809 _0114_ net6 0
C22810 hold13/a_391_47# _1037_/a_27_47# 0
C22811 _0662_/a_81_21# _0294_ 0.15052f
C22812 hold41/a_49_47# _0179_ 0.04594f
C22813 net246 _0345_ 0
C22814 net36 A[1] 0
C22815 _1001_/a_891_413# _0459_ 0
C22816 _0957_/a_32_297# _0213_ 0
C22817 _0259_ _0186_ 0
C22818 _1036_/a_27_47# clknet_1_1__leaf__0463_ 0.06863f
C22819 VPWR _0707_/a_75_199# 0.14297f
C22820 _0836_/a_68_297# clkbuf_1_0__f__0465_/a_110_47# 0.00511f
C22821 _0457_ clknet_1_0__leaf__0461_ 0.27365f
C22822 _0293_ _0288_ 0.00133f
C22823 hold67/a_49_47# acc0.A\[10\] 0.00101f
C22824 _1001_/a_27_47# _0586_/a_27_47# 0
C22825 net61 _0434_ 0
C22826 _0133_ _0561_/a_149_47# 0.0092f
C22827 _1035_/a_1059_315# _0132_ 0.00504f
C22828 _1035_/a_381_47# _0208_ 0
C22829 hold87/a_285_47# _0399_ 0
C22830 _0236_ _0219_ 0.00324f
C22831 net212 clkbuf_1_0__f__0465_/a_110_47# 0
C22832 clknet_1_0__leaf__0463_ acc0.A\[15\] 0.00117f
C22833 net23 _0213_ 0
C22834 _1047_/a_193_47# _1047_/a_381_47# 0.09503f
C22835 _1047_/a_634_159# _1047_/a_891_413# 0.03684f
C22836 _1047_/a_27_47# _1047_/a_561_413# 0.0027f
C22837 _0181_ control0.add 0.02053f
C22838 _1030_/a_466_413# _0339_ 0.00604f
C22839 _1030_/a_1059_315# _0338_ 0.00144f
C22840 _0206_ _1040_/a_975_413# 0.002f
C22841 comp0.B\[8\] _1040_/a_592_47# 0
C22842 clknet_1_1__leaf__0465_ net37 0.30041f
C22843 _0504_/a_27_47# _1014_/a_193_47# 0
C22844 _0322_ _0352_ 0
C22845 _0957_/a_304_297# _0472_ 0.01365f
C22846 hold1/a_285_47# _0987_/a_1059_315# 0.01504f
C22847 hold1/a_49_47# _0987_/a_891_413# 0.00773f
C22848 _0957_/a_220_297# _0475_ 0.00174f
C22849 _0632_/a_113_47# acc0.A\[18\] 0
C22850 _0714_/a_51_297# net163 0
C22851 clkbuf_1_1__f__0460_/a_110_47# _0333_ 0
C22852 _0573_/a_27_47# net1 0
C22853 _1041_/a_381_47# _0174_ 0
C22854 _0327_ _0352_ 0
C22855 _0664_/a_79_21# _0284_ 0.09304f
C22856 _0664_/a_382_297# _0285_ 0.00222f
C22857 _0343_ clknet_0__0458_ 0
C22858 _0582_/a_109_47# _0115_ 0
C22859 net58 _0833_/a_79_21# 0.01015f
C22860 hold98/a_49_47# pp[31] 0
C22861 hold52/a_49_47# _0574_/a_27_297# 0.00134f
C22862 net234 _1014_/a_1059_315# 0
C22863 _0456_ _1014_/a_193_47# 0
C22864 hold20/a_49_47# net89 0
C22865 net202 _0113_ 0
C22866 _1052_/a_891_413# _1052_/a_1017_47# 0.00617f
C22867 _1007_/a_381_47# _1007_/a_561_413# 0.00123f
C22868 _1007_/a_27_47# net93 0.22242f
C22869 _1007_/a_891_413# _1007_/a_975_413# 0.00851f
C22870 hold96/a_49_47# _1004_/a_381_47# 0.00167f
C22871 VPWR _0321_ 1.22493f
C22872 _0525_/a_81_21# _0522_/a_109_297# 0
C22873 _0476_ net33 0.28325f
C22874 _0113_ clknet_1_1__leaf__0463_ 0
C22875 _0432_ _0835_/a_215_47# 0.08478f
C22876 _0837_/a_81_21# _0440_ 0.12357f
C22877 hold39/a_285_47# comp0.B\[2\] 0
C22878 net240 hold93/a_391_47# 0.1316f
C22879 _0172_ _1044_/a_975_413# 0
C22880 hold69/a_285_47# _1006_/a_1059_315# 0.0054f
C22881 VPWR clkbuf_0__0460_/a_110_47# 1.4101f
C22882 _0292_ _0369_ 0.00156f
C22883 _1020_/a_891_413# _0352_ 0.04599f
C22884 _0179_ _1052_/a_975_413# 0
C22885 _0209_ net28 0
C22886 net190 _1027_/a_193_47# 0
C22887 _1021_/a_466_413# clknet_1_0__leaf__0461_ 0
C22888 _1021_/a_193_47# net107 0.01325f
C22889 _0983_/a_27_47# _0852_/a_35_297# 0
C22890 VPWR _0498_/a_245_297# 0.00593f
C22891 _0986_/a_27_47# _0840_/a_150_297# 0
C22892 _0986_/a_193_47# _0840_/a_68_297# 0
C22893 _0309_ _0181_ 0
C22894 _0223_ _0617_/a_68_297# 0
C22895 _0557_/a_512_297# VPWR 0.00628f
C22896 net189 net66 0
C22897 _0731_/a_299_297# _0462_ 0
C22898 _0734_/a_47_47# _0734_/a_377_297# 0.00899f
C22899 _0550_/a_240_47# clkbuf_1_0__f__0463_/a_110_47# 0
C22900 hold74/a_391_47# _0305_ 0.01474f
C22901 _0212_ net23 0
C22902 VPWR _0351_ 0.22658f
C22903 _0239_ clknet_1_1__leaf__0461_ 0
C22904 _1003_/a_1059_315# _0487_ 0
C22905 control0.state\[0\] _0951_/a_296_53# 0
C22906 control0.state\[1\] _0951_/a_209_311# 0.00874f
C22907 acc0.A\[12\] net4 0.42772f
C22908 _0669_/a_183_297# net41 0
C22909 comp0.B\[11\] net198 0.02648f
C22910 B[14] net22 0.0049f
C22911 _1011_/a_1017_47# _0109_ 0.002f
C22912 net97 net227 0
C22913 input6/a_75_212# net6 0.10848f
C22914 hold78/a_49_47# net41 0
C22915 _0216_ _0726_/a_149_47# 0
C22916 _0294_ _0582_/a_27_297# 0.00856f
C22917 _1033_/a_891_413# control0.reset 0
C22918 net69 clknet_1_0__leaf__0458_ 0.11053f
C22919 _1061_/a_466_413# comp0.B\[9\] 0
C22920 _0179_ net75 0.0109f
C22921 net61 acc0.A\[7\] 0
C22922 output42/a_27_47# pp[14] 0
C22923 pp[15] output41/a_27_47# 0.01115f
C22924 net61 _0989_/a_1059_315# 0.031f
C22925 _0243_ _0616_/a_215_47# 0
C22926 clknet_0__0462_ hold90/a_49_47# 0.00338f
C22927 _0983_/a_27_47# _0081_ 0.08952f
C22928 hold40/a_285_47# hold40/a_391_47# 0.41909f
C22929 hold75/a_49_47# _0082_ 0
C22930 _0983_/a_466_413# _0454_ 0
C22931 _0983_/a_634_159# _0455_ 0
C22932 _0368_ acc0.A\[24\] 0.02406f
C22933 _0286_ hold70/a_285_47# 0
C22934 _0283_ hold70/a_391_47# 0
C22935 net21 comp0.B\[14\] 0.06586f
C22936 _0369_ _0435_ 0.0033f
C22937 _1059_/a_1059_315# _0277_ 0
C22938 _1063_/a_634_159# _1063_/a_1059_315# 0
C22939 _1063_/a_27_47# _1063_/a_381_47# 0.05761f
C22940 _1063_/a_193_47# _1063_/a_891_413# 0.19226f
C22941 _0645_/a_285_47# acc0.A\[15\] 0.00396f
C22942 _0183_ _0374_ 0
C22943 clkbuf_0_clk/a_110_47# net159 0.01893f
C22944 clkbuf_1_1__f__0458_/a_110_47# _0826_/a_27_53# 0
C22945 _1019_/a_466_413# _0346_ 0.00617f
C22946 hold86/a_285_47# _0465_ 0.00673f
C22947 _0179_ _0513_/a_299_297# 0.11984f
C22948 acc0.A\[8\] _0830_/a_79_21# 0
C22949 hold19/a_49_47# net221 0
C22950 _1037_/a_466_413# _0208_ 0
C22951 net159 _1063_/a_634_159# 0
C22952 _0218_ _0869_/a_27_47# 0.00151f
C22953 _0195_ acc0.A\[3\] 0.05631f
C22954 _1063_/a_891_413# _0460_ 0.00323f
C22955 _0786_/a_300_47# _0402_ 0
C22956 _0462_ _1006_/a_634_159# 0.00424f
C22957 acc0.A\[1\] acc0.A\[18\] 0
C22958 net36 clkbuf_0__0463_/a_110_47# 0
C22959 hold86/a_49_47# net58 0.04371f
C22960 hold86/a_285_47# acc0.A\[2\] 0
C22961 net46 _1022_/a_27_47# 0
C22962 _0172_ _0180_ 0.0245f
C22963 B[1] B[2] 0.00498f
C22964 _1039_/a_891_413# _0177_ 0
C22965 _0183_ _0507_/a_27_297# 0.09619f
C22966 _0195_ control0.sh 0
C22967 hold52/a_391_47# _1025_/a_27_47# 0
C22968 _0200_ clkbuf_0__0464_/a_110_47# 0
C22969 net63 _0252_ 0.09555f
C22970 net63 _0989_/a_381_47# 0.00911f
C22971 B[12] comp0.B\[10\] 0
C22972 _0172_ net152 0.09564f
C22973 hold74/a_285_47# net43 0.00186f
C22974 _0820_/a_215_47# net66 0
C22975 _0820_/a_79_21# _0291_ 0
C22976 _0760_/a_377_297# _0219_ 0
C22977 _0663_/a_27_413# _0295_ 0
C22978 _1004_/a_381_47# net90 0
C22979 _1011_/a_381_47# acc0.A\[29\] 0.00155f
C22980 _1004_/a_193_47# _1024_/a_1059_315# 0
C22981 _1004_/a_27_47# _1024_/a_891_413# 0
C22982 _0183_ net165 0.03339f
C22983 _0306_ _0352_ 0.0586f
C22984 _0576_/a_27_297# _0352_ 0
C22985 A[14] _0797_/a_27_413# 0
C22986 _1060_/a_634_159# _1060_/a_1059_315# 0
C22987 _1060_/a_27_47# _1060_/a_381_47# 0.06222f
C22988 _1060_/a_193_47# _1060_/a_891_413# 0.19489f
C22989 _0179_ net138 0.24444f
C22990 net198 _0202_ 0.00305f
C22991 _0513_/a_81_21# _0513_/a_299_297# 0.08213f
C22992 _1051_/a_27_47# _0527_/a_27_297# 0
C22993 _0733_/a_79_199# _0319_ 0.17021f
C22994 net114 _1008_/a_193_47# 0
C22995 _1028_/a_193_47# net94 0
C22996 _0510_/a_373_47# acc0.A\[10\] 0.00321f
C22997 _1070_/a_27_47# _0480_ 0.00313f
C22998 hold43/a_391_47# _1028_/a_1059_315# 0.01554f
C22999 net126 _1040_/a_27_47# 0.22171f
C23000 pp[26] _0124_ 0
C23001 _0734_/a_47_47# clknet_0__0462_ 0
C23002 _1053_/a_27_47# net11 0.00457f
C23003 _0432_ _0172_ 0.01238f
C23004 _0143_ _1050_/a_466_413# 0
C23005 _1039_/a_466_413# comp0.B\[9\] 0
C23006 _0805_/a_181_47# clknet_1_1__leaf__0459_ 0
C23007 _1039_/a_1059_315# _0555_/a_51_297# 0
C23008 clknet_1_1__leaf__0463_ comp0.B\[3\] 0.08589f
C23009 _0343_ net178 0.02244f
C23010 _0467_ _0971_/a_384_47# 0
C23011 _0988_/a_466_413# net74 0
C23012 net175 net247 0
C23013 _0553_/a_51_297# _0174_ 0.09878f
C23014 _1067_/a_634_159# clknet_1_1__leaf_clk 0
C23015 pp[29] _0355_ 0
C23016 _0787_/a_80_21# _0218_ 0.00276f
C23017 net70 _0983_/a_1059_315# 0
C23018 _0984_/a_1059_315# net69 0
C23019 _0181_ clknet_1_1__leaf__0457_ 0.36081f
C23020 _0968_/a_109_297# net34 0
C23021 _0968_/a_193_297# control0.state\[1\] 0.00332f
C23022 net56 _1011_/a_193_47# 0
C23023 pp[27] _0568_/a_109_297# 0
C23024 VPWR _1009_/a_27_47# 0.69985f
C23025 _1053_/a_891_413# _0252_ 0
C23026 net84 _0781_/a_68_297# 0.0012f
C23027 _0366_ clknet_0__0460_ 0
C23028 clknet_1_0__leaf__0460_ _0757_/a_150_297# 0
C23029 _0312_ _0350_ 0.02553f
C23030 _0183_ acc0.A\[19\] 0.11998f
C23031 _1041_/a_1059_315# comp0.B\[8\] 0
C23032 _1041_/a_466_413# _0206_ 0
C23033 _0217_ _0242_ 0.00222f
C23034 _0347_ _0301_ 0
C23035 VPWR _0146_ 0.38475f
C23036 _0982_/a_561_413# _0465_ 0
C23037 _0195_ _0851_/a_113_47# 0
C23038 net45 net99 0.02398f
C23039 _0753_/a_465_47# _0378_ 0
C23040 _0233_ _0756_/a_47_47# 0
C23041 _0504_/a_27_47# clknet_0__0457_ 0
C23042 _1071_/a_27_47# _0168_ 0
C23043 VPWR _1014_/a_891_413# 0.17569f
C23044 _1071_/a_634_159# VPWR 0.18497f
C23045 net58 acc0.A\[14\] 0.01692f
C23046 _0326_ clknet_1_0__leaf__0460_ 0
C23047 _0678_/a_68_297# _0397_ 0.02076f
C23048 _0203_ net195 0
C23049 net53 _0319_ 0.00773f
C23050 VPWR _0492_/a_27_47# 0.23518f
C23051 _0856_/a_79_21# _0452_ 0
C23052 clknet_1_0__leaf__0457_ _0772_/a_297_297# 0
C23053 _0984_/a_193_47# hold75/a_49_47# 0
C23054 _0984_/a_27_47# hold75/a_285_47# 0
C23055 hold28/a_49_47# clknet_1_0__leaf__0464_ 0
C23056 acc0.A\[15\] _0507_/a_27_297# 0.01027f
C23057 _0329_ hold95/a_391_47# 0
C23058 net82 _1060_/a_1059_315# 0.00146f
C23059 _0172_ _1042_/a_466_413# 0.002f
C23060 clknet_0__0457_ _0456_ 0
C23061 acc0.A\[27\] _0569_/a_27_297# 0
C23062 hold59/a_49_47# acc0.A\[1\] 0
C23063 _0195_ net157 0.00188f
C23064 _1021_/a_561_413# _0460_ 0
C23065 net121 B[4] 0
C23066 _1021_/a_592_47# clknet_1_0__leaf__0457_ 0
C23067 _0361_ _0685_/a_68_297# 0
C23068 net193 clkbuf_0__0464_/a_110_47# 0
C23069 _0253_ _0186_ 0.0123f
C23070 _0680_/a_217_297# _0250_ 0
C23071 _0716_/a_27_47# acc0.A\[15\] 0
C23072 net36 hold71/a_49_47# 0
C23073 _0080_ hold60/a_285_47# 0
C23074 _0891_/a_27_47# _0352_ 0
C23075 net153 net174 0
C23076 _1067_/a_466_413# clkbuf_1_1__f_clk/a_110_47# 0
C23077 _0257_ _0271_ 0.09301f
C23078 _0258_ _0270_ 0
C23079 net165 acc0.A\[15\] 0.00772f
C23080 _0309_ _0677_/a_377_297# 0.00188f
C23081 hold35/a_49_47# acc0.A\[9\] 0.00307f
C23082 _0992_/a_634_159# net143 0
C23083 clkbuf_0__0464_/a_110_47# _1046_/a_466_413# 0.00635f
C23084 _0535_/a_150_297# _0473_ 0
C23085 hold79/a_49_47# control0.count\[0\] 0.00271f
C23086 output54/a_27_47# _1027_/a_193_47# 0
C23087 hold67/a_285_47# _0181_ 0
C23088 _0144_ _0465_ 0
C23089 _1008_/a_193_47# _0365_ 0.03876f
C23090 _0313_ _0697_/a_80_21# 0.14039f
C23091 clknet_1_1__leaf__0465_ _0505_/a_27_297# 0.04202f
C23092 _0228_ _0382_ 0.00555f
C23093 _0718_/a_47_47# _1030_/a_466_413# 0
C23094 net175 _1048_/a_466_413# 0
C23095 net9 _1048_/a_27_47# 0.0253f
C23096 _0370_ _0219_ 0.00275f
C23097 VPWR input28/a_75_212# 0.25724f
C23098 _0179_ _0442_ 0
C23099 hold25/a_285_47# _1038_/a_466_413# 0.00377f
C23100 hold25/a_391_47# _1038_/a_634_159# 0.00125f
C23101 hold25/a_49_47# _1038_/a_1059_315# 0
C23102 clknet_1_0__leaf__0457_ _0208_ 0.19644f
C23103 _0958_/a_27_47# _1062_/a_193_47# 0
C23104 _0538_/a_51_297# _1045_/a_1059_315# 0
C23105 _0538_/a_240_47# _1045_/a_27_47# 0
C23106 _0538_/a_149_47# _1045_/a_193_47# 0
C23107 net44 _0779_/a_297_297# 0.00561f
C23108 net22 _0544_/a_51_297# 0
C23109 net149 _1047_/a_193_47# 0.03785f
C23110 output66/a_27_47# A[10] 0.0066f
C23111 hold74/a_391_47# _0181_ 0
C23112 hold13/a_49_47# _0473_ 0.03566f
C23113 VPWR _1022_/a_193_47# 0.32103f
C23114 clknet_1_1__leaf__0460_ _0680_/a_300_47# 0
C23115 _0285_ _0402_ 0.3843f
C23116 hold75/a_49_47# clkbuf_0__0458_/a_110_47# 0
C23117 net23 _0161_ 0
C23118 _0553_/a_51_297# _0208_ 0.16074f
C23119 net85 _0790_/a_117_297# 0
C23120 clknet_1_1__leaf__0459_ _0993_/a_27_47# 0.00145f
C23121 _0993_/a_634_159# net38 0
C23122 _0999_/a_27_47# _0999_/a_634_159# 0.14145f
C23123 _0820_/a_79_21# _0290_ 0.01314f
C23124 hold13/a_391_47# _0133_ 0
C23125 _0083_ _0447_ 0.02491f
C23126 VPWR _0771_/a_27_413# 0.25648f
C23127 _1017_/a_193_47# net221 0
C23128 clknet_1_0__leaf__0462_ _0320_ 0
C23129 A[0] rst 0.11142f
C23130 hold24/a_49_47# control0.sh 0
C23131 _1001_/a_466_413# _0772_/a_215_47# 0.00141f
C23132 hold32/a_49_47# _0179_ 0
C23133 clknet_1_0__leaf__0465_ _0989_/a_27_47# 0
C23134 clknet_1_0__leaf__0465_ hold1/a_49_47# 0.03597f
C23135 net120 _1034_/a_27_47# 0.23081f
C23136 _0991_/a_891_413# _0345_ 0
C23137 hold58/a_285_47# VPWR 0.30039f
C23138 hold47/a_391_47# clknet_1_0__leaf__0464_ 0
C23139 acc0.A\[16\] net102 0
C23140 _1035_/a_1059_315# net25 0.02777f
C23141 hold86/a_49_47# _0262_ 0
C23142 net185 _0959_/a_80_21# 0
C23143 _1062_/a_27_47# _0160_ 0.07749f
C23144 _1062_/a_1059_315# _1062_/a_1017_47# 0
C23145 net55 _0729_/a_150_297# 0
C23146 clknet_1_1__leaf__0465_ _0506_/a_81_21# 0.01507f
C23147 _0679_/a_68_297# clkbuf_0__0461_/a_110_47# 0
C23148 _1011_/a_1059_315# _0353_ 0
C23149 input19/a_75_212# B[11] 0.19715f
C23150 _0738_/a_68_297# hold50/a_285_47# 0
C23151 net39 _0647_/a_377_297# 0.00586f
C23152 acc0.A\[12\] _0647_/a_47_47# 0.10358f
C23153 acc0.A\[9\] A[9] 0.21264f
C23154 _0459_ net149 0
C23155 _1021_/a_634_159# _1021_/a_975_413# 0
C23156 _1021_/a_466_413# _1021_/a_561_413# 0.00772f
C23157 net199 _1024_/a_1059_315# 0.0016f
C23158 _0454_ _0452_ 0
C23159 _1017_/a_466_413# _0459_ 0.00164f
C23160 clkbuf_1_0__f__0459_/a_110_47# net229 0
C23161 _0147_ _1048_/a_1059_315# 0.00459f
C23162 _1049_/a_891_413# net134 0
C23163 net144 pp[10] 0
C23164 _0476_ _0563_/a_149_47# 0
C23165 _0222_ net50 0.05646f
C23166 _0732_/a_209_297# _0742_/a_299_297# 0
C23167 _0732_/a_80_21# _0742_/a_384_47# 0
C23168 net35 _0161_ 0
C23169 hold15/a_391_47# net60 0
C23170 net162 _0708_/a_68_297# 0
C23171 control0.state\[1\] _0181_ 0.02581f
C23172 _0329_ acc0.A\[28\] 0.02368f
C23173 _0179_ net165 0
C23174 _0733_/a_79_199# _0733_/a_448_47# 0.04614f
C23175 _0853_/a_68_297# _0347_ 0
C23176 _0963_/a_117_297# clk 0
C23177 hold65/a_285_47# _0274_ 0.00183f
C23178 net62 _0988_/a_634_159# 0.00506f
C23179 _0181_ _0583_/a_109_47# 0
C23180 _0346_ _0352_ 0.05208f
C23181 _0556_/a_68_297# VPWR 0.15406f
C23182 hold98/a_391_47# net42 0
C23183 _1011_/a_193_47# _0345_ 0.03268f
C23184 hold87/a_391_47# net36 0.08616f
C23185 net48 _1022_/a_193_47# 0.03437f
C23186 clkbuf_1_0__f__0465_/a_110_47# _0989_/a_891_413# 0
C23187 _1031_/a_466_413# _1013_/a_193_47# 0
C23188 _1031_/a_193_47# _1013_/a_466_413# 0
C23189 _1031_/a_634_159# _1013_/a_634_159# 0
C23190 net34 _0486_ 0.33173f
C23191 _0434_ _0431_ 0
C23192 clknet_1_1__leaf__0464_ _1043_/a_1017_47# 0.00109f
C23193 _0234_ _0378_ 0.00334f
C23194 _0216_ _0568_/a_109_297# 0.01141f
C23195 _1046_/a_634_159# net147 0
C23196 _0248_ _0242_ 0.14556f
C23197 clknet_1_1__leaf__0459_ _0409_ 0
C23198 hold57/a_49_47# VPWR 0.26974f
C23199 _0953_/a_114_297# comp0.B\[8\] 0.01459f
C23200 _0953_/a_32_297# _0206_ 0
C23201 net45 _0396_ 0.00343f
C23202 VPWR _0978_/a_27_297# 0.23033f
C23203 _1034_/a_1059_315# clknet_0__0463_ 0.00602f
C23204 VPWR _0795_/a_81_21# 0.2143f
C23205 hold97/a_49_47# net54 0.32403f
C23206 hold19/a_49_47# _1017_/a_27_47# 0
C23207 hold85/a_49_47# hold85/a_285_47# 0.22264f
C23208 _0780_/a_35_297# _0780_/a_117_297# 0.00641f
C23209 clknet_1_0__leaf__0465_ _0538_/a_51_297# 0.00237f
C23210 hold17/a_49_47# _1071_/a_466_413# 0
C23211 hold78/a_391_47# net225 0.13583f
C23212 hold78/a_49_47# _0111_ 0
C23213 comp0.B\[5\] _0562_/a_150_297# 0
C23214 _0259_ net62 0.02529f
C23215 _0352_ hold94/a_49_47# 0
C23216 _0750_/a_181_47# _0460_ 0
C23217 hold49/a_285_47# _0174_ 0
C23218 _0221_ acc0.A\[28\] 0.18519f
C23219 _0561_/a_149_47# _0208_ 0.01788f
C23220 _0561_/a_245_297# _0132_ 0.00161f
C23221 VPWR _1067_/a_466_413# 0.2627f
C23222 _0717_/a_209_297# pp[17] 0
C23223 clknet_0__0460_ _0689_/a_68_297# 0
C23224 _1050_/a_193_47# _0186_ 0.02714f
C23225 net53 _0733_/a_448_47# 0
C23226 net17 _1062_/a_634_159# 0
C23227 _0498_/a_51_297# _0913_/a_27_47# 0
C23228 _1033_/a_193_47# clknet_1_0__leaf__0461_ 0
C23229 _0228_ _1005_/a_634_159# 0
C23230 _0982_/a_1059_315# _0263_ 0
C23231 _1021_/a_27_47# net17 0
C23232 _0381_ clknet_1_0__leaf__0460_ 0.00193f
C23233 hold88/a_391_47# net58 0
C23234 _0640_/a_392_297# _0271_ 0
C23235 net149 _0265_ 0.00176f
C23236 _1020_/a_891_413# net106 0
C23237 _0372_ clkbuf_1_0__f__0460_/a_110_47# 0
C23238 net188 _0181_ 0
C23239 _0527_/a_27_297# _0085_ 0
C23240 hold14/a_285_47# hold14/a_391_47# 0.41909f
C23241 VPWR _0338_ 0.45226f
C23242 _0243_ _0771_/a_215_297# 0.14931f
C23243 _0389_ _0771_/a_298_297# 0.04274f
C23244 _0390_ _0771_/a_27_413# 0.25154f
C23245 _0348_ _1030_/a_1059_315# 0.0014f
C23246 _0555_/a_51_297# _1037_/a_1059_315# 0.01354f
C23247 _0555_/a_240_47# _1037_/a_27_47# 0
C23248 _0586_/a_27_47# _0772_/a_79_21# 0
C23249 _0683_/a_113_47# _0219_ 0
C23250 _0313_ _0345_ 0.17444f
C23251 _0401_ _0814_/a_181_47# 0.00242f
C23252 _0746_/a_81_21# _0370_ 0.01759f
C23253 _0309_ clknet_1_1__leaf__0461_ 0.00477f
C23254 _0458_ _0640_/a_215_297# 0
C23255 hold69/a_49_47# _0679_/a_68_297# 0
C23256 _0372_ _0250_ 0
C23257 _0179_ hold83/a_285_47# 0
C23258 _1041_/a_592_47# net153 0.00116f
C23259 _1041_/a_381_47# comp0.B\[9\] 0
C23260 net47 net146 0
C23261 _1047_/a_1059_315# _0145_ 0
C23262 _0573_/a_27_47# control0.sh 0
C23263 net45 _0790_/a_117_297# 0
C23264 A[5] net11 0.03972f
C23265 _1003_/a_1059_315# _0760_/a_47_47# 0.00115f
C23266 hold12/a_285_47# _0382_ 0
C23267 _0111_ _0129_ 0
C23268 clknet_1_0__leaf_clk _0484_ 0.00121f
C23269 net157 _1048_/a_193_47# 0
C23270 comp0.B\[1\] _0214_ 0.00394f
C23271 net185 _0173_ 0.08588f
C23272 pp[28] _0109_ 0
C23273 _0216_ net176 0
C23274 _0567_/a_27_297# acc0.A\[30\] 0.06619f
C23275 _0953_/a_32_297# _1046_/a_1059_315# 0
C23276 _0217_ _1018_/a_1017_47# 0
C23277 _0458_ _0465_ 0.01279f
C23278 _0536_/a_240_47# _0472_ 0
C23279 net243 _1004_/a_1017_47# 0
C23280 output44/a_27_47# hold15/a_285_47# 0.00395f
C23281 _0123_ _1007_/a_193_47# 0
C23282 _0441_ _0442_ 0.14354f
C23283 _0231_ _0183_ 0
C23284 _0518_/a_109_297# _0186_ 0.02631f
C23285 _0994_/a_27_47# net246 0
C23286 _0451_ _0263_ 0
C23287 net197 net156 0.06731f
C23288 _0119_ clknet_1_0__leaf__0461_ 0.00655f
C23289 _0544_/a_51_297# _0544_/a_245_297# 0.01218f
C23290 clkbuf_1_0__f__0461_/a_110_47# _0611_/a_68_297# 0.00543f
C23291 _0643_/a_103_199# _0433_ 0
C23292 _0733_/a_222_93# _0317_ 0
C23293 hold7/a_285_47# _0987_/a_381_47# 0
C23294 acc0.A\[2\] _0458_ 0.02649f
C23295 _0134_ VPWR 0.31932f
C23296 _0956_/a_32_297# control0.reset 0.01469f
C23297 _0734_/a_285_47# _0362_ 0.04448f
C23298 _0183_ net1 1.2325f
C23299 _0514_/a_373_47# net142 0
C23300 _1034_/a_27_47# _1034_/a_466_413# 0.26005f
C23301 _1034_/a_193_47# _1034_/a_634_159# 0.12729f
C23302 _0536_/a_51_297# _0536_/a_512_297# 0.0116f
C23303 _1021_/a_27_47# acc0.A\[21\] 0
C23304 net168 _1053_/a_634_159# 0
C23305 _0559_/a_51_297# hold58/a_391_47# 0
C23306 hold10/a_391_47# comp0.B\[15\] 0
C23307 _0430_ _0826_/a_219_297# 0.04404f
C23308 _0294_ _0115_ 0.03683f
C23309 net104 _0580_/a_109_297# 0
C23310 comp0.B\[7\] VPWR 0.88969f
C23311 _1057_/a_975_413# net67 0
C23312 hold25/a_285_47# _0550_/a_240_47# 0
C23313 _0982_/a_1059_315# clknet_1_0__leaf__0461_ 0
C23314 _0459_ _0094_ 0.00198f
C23315 _1038_/a_891_413# net28 0
C23316 _0217_ _0855_/a_81_21# 0.05858f
C23317 _0516_/a_27_297# acc0.A\[9\] 0.06665f
C23318 net69 _0455_ 0.08361f
C23319 net39 _0802_/a_59_75# 0.0682f
C23320 clkbuf_0__0464_/a_110_47# _1045_/a_193_47# 0.00244f
C23321 clkbuf_0__0463_/a_110_47# _0563_/a_149_47# 0
C23322 _1063_/a_466_413# _0161_ 0.0345f
C23323 clknet_0__0460_ acc0.A\[24\] 0.00948f
C23324 net235 _0988_/a_193_47# 0.00112f
C23325 _0218_ _0796_/a_79_21# 0
C23326 net205 control0.sh 0
C23327 _0746_/a_299_297# _0350_ 0
C23328 VPWR _1026_/a_27_47# 0.64275f
C23329 _0854_/a_297_297# acc0.A\[18\] 0.00129f
C23330 _0525_/a_81_21# _0150_ 0
C23331 _0573_/a_27_47# net157 0.02135f
C23332 control0.count\[3\] _1072_/a_193_47# 0.05485f
C23333 net207 _0346_ 0.37846f
C23334 _0712_/a_79_21# _1013_/a_1059_315# 0
C23335 net78 _0992_/a_193_47# 0.00678f
C23336 net194 clkbuf_1_1__f__0464_/a_110_47# 0.00584f
C23337 _0135_ _0208_ 0.02322f
C23338 _0182_ hold2/a_391_47# 0.00568f
C23339 _0230_ _0101_ 0
C23340 VPWR _1024_/a_1059_315# 0.41434f
C23341 _0959_/a_217_297# _0470_ 0.01042f
C23342 hold13/a_49_47# hold13/a_285_47# 0.22264f
C23343 _0257_ clknet_1_0__leaf__0465_ 0.30149f
C23344 VPWR net99 0.41411f
C23345 _0462_ net92 0.0221f
C23346 _0172_ _0498_/a_51_297# 0.14732f
C23347 _0585_/a_109_297# net149 0.00305f
C23348 net203 _0563_/a_512_297# 0
C23349 clkbuf_1_1__f__0462_/a_110_47# _0319_ 0.00552f
C23350 _0402_ _0218_ 0.00681f
C23351 _0982_/a_891_413# net47 0.00359f
C23352 acc0.A\[17\] _0674_/a_113_47# 0
C23353 net36 _0264_ 0.33457f
C23354 _0446_ _0186_ 0
C23355 VPWR _1048_/a_381_47# 0.07678f
C23356 pp[30] _0567_/a_109_47# 0
C23357 net18 _0542_/a_240_47# 0.00222f
C23358 acc0.A\[4\] hold7/a_285_47# 0.00795f
C23359 _0183_ _0185_ 0
C23360 input2/a_75_212# _0186_ 0.01058f
C23361 _0144_ clknet_0__0464_ 0
C23362 net232 _1062_/a_381_47# 0
C23363 _0731_/a_299_297# _0312_ 0.06059f
C23364 _1028_/a_1017_47# clknet_1_1__leaf__0462_ 0
C23365 _1017_/a_27_47# _1017_/a_193_47# 0.96574f
C23366 net45 acc0.A\[31\] 0.10653f
C23367 output55/a_27_47# _0353_ 0
C23368 output64/a_27_47# net141 0
C23369 _0361_ _0368_ 0
C23370 _0427_ clknet_0__0465_ 0.13535f
C23371 net194 _0186_ 0
C23372 hold13/a_391_47# _0174_ 0
C23373 _0472_ _1046_/a_27_47# 0
C23374 _0473_ _1046_/a_634_159# 0.00647f
C23375 _0984_/a_27_47# _0345_ 0
C23376 _0343_ _0675_/a_68_297# 0
C23377 net57 acc0.A\[29\] 0.50929f
C23378 hold101/a_49_47# _0255_ 0
C23379 net194 hold49/a_49_47# 0
C23380 net197 acc0.A\[26\] 0.02118f
C23381 VPWR _1010_/a_1017_47# 0
C23382 _1000_/a_634_159# _1000_/a_975_413# 0
C23383 _1000_/a_466_413# _1000_/a_561_413# 0.00772f
C23384 _1000_/a_193_47# _1000_/a_592_47# 0
C23385 _0600_/a_103_199# clknet_1_0__leaf__0460_ 0.01381f
C23386 _0993_/a_193_47# _0281_ 0.00378f
C23387 _1060_/a_466_413# _0158_ 0.00473f
C23388 _1060_/a_1059_315# net146 0
C23389 VPWR _0797_/a_297_47# 0
C23390 _0271_ clknet_1_1__leaf__0458_ 0.08283f
C23391 control0.count\[1\] _0979_/a_109_297# 0.0011f
C23392 hold43/a_49_47# acc0.A\[28\] 0.33385f
C23393 _0459_ _0508_/a_299_297# 0
C23394 _0305_ _0998_/a_27_47# 0
C23395 _0399_ acc0.A\[9\] 0.0216f
C23396 _0457_ _0112_ 0
C23397 hold55/a_49_47# clknet_1_0__leaf__0457_ 0
C23398 _1072_/a_1059_315# VPWR 0.39768f
C23399 _0277_ hold91/a_49_47# 0
C23400 _0640_/a_215_297# clkbuf_1_1__f__0458_/a_110_47# 0
C23401 clkbuf_0__0463_/a_110_47# _1061_/a_27_47# 0.0012f
C23402 clknet_1_1__leaf__0458_ _0987_/a_891_413# 0.00101f
C23403 _0554_/a_68_297# VPWR 0.15912f
C23404 clknet_0__0458_ _0842_/a_59_75# 0.00483f
C23405 _0953_/a_304_297# comp0.B\[9\] 0.01441f
C23406 hold56/a_285_47# control0.reset 0.00899f
C23407 _0269_ _0434_ 0
C23408 acc0.A\[12\] _0287_ 0
C23409 _0399_ _0986_/a_592_47# 0
C23410 _0661_/a_27_297# _0424_ 0
C23411 _0292_ _0817_/a_81_21# 0
C23412 net240 _1063_/a_193_47# 0
C23413 _0346_ _0849_/a_79_21# 0
C23414 _0136_ comp0.B\[10\] 0
C23415 _0399_ _0670_/a_79_21# 0
C23416 _0736_/a_56_297# _1009_/a_193_47# 0
C23417 _0457_ _1033_/a_891_413# 0.00905f
C23418 _0343_ _0618_/a_79_21# 0.02192f
C23419 _1002_/a_1059_315# _0228_ 0
C23420 _0583_/a_27_297# _0114_ 0.11527f
C23421 net240 _0460_ 0.02498f
C23422 _0459_ _0393_ 0.01019f
C23423 _1072_/a_27_47# clkbuf_1_0__f_clk/a_110_47# 0.0071f
C23424 _1050_/a_27_47# _1050_/a_466_413# 0.27314f
C23425 _1050_/a_193_47# _1050_/a_634_159# 0.12497f
C23426 hold59/a_285_47# _0854_/a_79_21# 0
C23427 _1056_/a_381_47# net178 0
C23428 _0465_ clkbuf_1_1__f__0458_/a_110_47# 0.0013f
C23429 _0253_ net62 0
C23430 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# 1.66474f
C23431 hold37/a_391_47# clknet_0__0464_ 0.03083f
C23432 _0959_/a_300_47# _0160_ 0
C23433 _1019_/a_193_47# clknet_1_0__leaf__0457_ 0
C23434 _0557_/a_51_297# comp0.B\[5\] 0.01671f
C23435 _0985_/a_592_47# _0179_ 0.00253f
C23436 _0443_ _0826_/a_219_297# 0
C23437 _1032_/a_193_47# control0.reset 0
C23438 hold85/a_285_47# net17 0.05926f
C23439 net224 _1010_/a_27_47# 0
C23440 acc0.A\[15\] _0185_ 0.04549f
C23441 hold74/a_391_47# clknet_1_1__leaf__0461_ 0.08187f
C23442 _0221_ _1011_/a_634_159# 0.01531f
C23443 clknet_1_1__leaf__0460_ _0780_/a_117_297# 0
C23444 clknet_1_1__leaf__0463_ _1065_/a_1059_315# 0.00892f
C23445 acc0.A\[27\] _0127_ 0
C23446 _0179_ _1049_/a_381_47# 0.00461f
C23447 _1018_/a_1059_315# _0181_ 0
C23448 _0819_/a_384_47# _0401_ 0.00954f
C23449 net232 net185 0
C23450 _1059_/a_975_413# _0219_ 0
C23451 _1036_/a_27_47# input28/a_75_212# 0
C23452 _0778_/a_68_297# _0352_ 0.03704f
C23453 _0999_/a_466_413# _1012_/a_193_47# 0
C23454 _0999_/a_634_159# _1012_/a_634_159# 0
C23455 _0999_/a_193_47# _1012_/a_466_413# 0
C23456 _0499_/a_59_75# _0208_ 0
C23457 _0365_ _0318_ 0
C23458 clknet_0__0464_ _1046_/a_592_47# 0.00282f
C23459 _0997_/a_1059_315# pp[14] 0
C23460 _0997_/a_381_47# net41 0.01647f
C23461 _0359_ _0460_ 0
C23462 _1054_/a_27_47# _1052_/a_27_47# 0.0011f
C23463 net54 _1027_/a_592_47# 0.00131f
C23464 _1008_/a_1017_47# _0106_ 0
C23465 _0670_/a_297_297# _0277_ 0
C23466 clknet_1_1__leaf__0465_ _0184_ 0.22363f
C23467 hold13/a_391_47# _0208_ 0.00194f
C23468 net224 _1009_/a_193_47# 0
C23469 hold33/a_49_47# VPWR 0.25714f
C23470 net85 net43 0
C23471 _1039_/a_27_47# clkbuf_0__0463_/a_110_47# 0.00644f
C23472 _0538_/a_51_297# _1044_/a_466_413# 0
C23473 _0538_/a_149_47# _1044_/a_27_47# 0
C23474 _0178_ _1047_/a_381_47# 0.01234f
C23475 output38/a_27_47# VPWR 0.27531f
C23476 _0577_/a_373_47# VPWR 0
C23477 comp0.B\[11\] _1043_/a_592_47# 0
C23478 hold25/a_285_47# net172 0.01095f
C23479 net46 _0756_/a_285_47# 0.00644f
C23480 acc0.A\[14\] _1060_/a_466_413# 0
C23481 _0477_ _1062_/a_193_47# 0.03338f
C23482 pp[28] _0725_/a_80_21# 0.00741f
C23483 hold46/a_49_47# hold46/a_391_47# 0.00188f
C23484 control0.state\[2\] _1068_/a_1059_315# 0
C23485 _0486_ _1068_/a_466_413# 0.0372f
C23486 hold27/a_49_47# net174 0
C23487 _0200_ _0535_/a_150_297# 0
C23488 net21 _1045_/a_891_413# 0.00412f
C23489 _0143_ _1045_/a_634_159# 0
C23490 hold58/a_285_47# _1036_/a_27_47# 0
C23491 hold58/a_49_47# _1036_/a_193_47# 0
C23492 net46 _0749_/a_299_297# 0
C23493 _0399_ _0449_ 0
C23494 _0606_/a_109_53# _0460_ 0.00198f
C23495 _0973_/a_27_297# _0973_/a_109_297# 0.17136f
C23496 clknet_1_0__leaf__0465_ net11 0.0394f
C23497 _0531_/a_27_297# clknet_1_1__leaf__0457_ 0.00169f
C23498 hold70/a_391_47# _0345_ 0.00252f
C23499 pp[30] net208 0.00799f
C23500 _1033_/a_634_159# _0173_ 0
C23501 _0343_ _1000_/a_634_159# 0.00515f
C23502 _0328_ net216 0.00183f
C23503 _0179_ _0426_ 0
C23504 VPWR _0396_ 0.22323f
C23505 _0537_/a_68_297# net20 0
C23506 _0999_/a_891_413# _0999_/a_975_413# 0.00851f
C23507 _0999_/a_27_47# net85 0.22381f
C23508 _0999_/a_381_47# _0999_/a_561_413# 0.00123f
C23509 acc0.A\[17\] _0307_ 0.10197f
C23510 net17 _1063_/a_592_47# 0.00259f
C23511 _0339_ _0567_/a_109_47# 0
C23512 net239 _0347_ 0
C23513 _1001_/a_193_47# _1019_/a_1059_315# 0
C23514 _1001_/a_27_47# _1019_/a_891_413# 0
C23515 _0772_/a_215_47# _0772_/a_510_47# 0.00529f
C23516 _0754_/a_512_297# _0103_ 0
C23517 VPWR _0993_/a_1059_315# 0.41898f
C23518 _1001_/a_381_47# _0099_ 0.13563f
C23519 _0535_/a_68_297# _0206_ 0
C23520 hold76/a_285_47# _0350_ 0
C23521 _1021_/a_27_47# _0165_ 0.00105f
C23522 _0601_/a_68_297# _0360_ 0
C23523 _0752_/a_27_413# _0752_/a_300_297# 0.00737f
C23524 _0663_/a_27_413# _0346_ 0.02895f
C23525 _0565_/a_240_47# comp0.B\[0\] 0.00136f
C23526 hold68/a_285_47# _1024_/a_27_47# 0.00861f
C23527 clknet_1_0__leaf__0462_ _1007_/a_1059_315# 0.00475f
C23528 _0298_ hold91/a_49_47# 0
C23529 _0404_ hold91/a_285_47# 0
C23530 hold24/a_391_47# net29 0
C23531 _0697_/a_80_21# _0321_ 0.02835f
C23532 VPWR _0580_/a_27_297# 0.2054f
C23533 _0131_ _0957_/a_32_297# 0
C23534 _0983_/a_27_47# _0183_ 0
C23535 _0983_/a_634_159# _0217_ 0
C23536 _0346_ _0237_ 0.00213f
C23537 hold88/a_285_47# net47 0.031f
C23538 pp[28] _0128_ 0
C23539 clkbuf_1_1__f__0465_/a_110_47# _0369_ 0.01465f
C23540 _0186_ _0987_/a_193_47# 0
C23541 net67 _0304_ 0
C23542 _0179_ _0185_ 0.10907f
C23543 _1043_/a_27_47# _0542_/a_149_47# 0
C23544 _0556_/a_68_297# _1036_/a_27_47# 0
C23545 _0232_ _0345_ 0
C23546 _0695_/a_217_297# clkbuf_0__0460_/a_110_47# 0.0028f
C23547 hold100/a_391_47# _0267_ 0
C23548 net245 net43 0.00166f
C23549 _1021_/a_561_413# _0119_ 0
C23550 _1001_/a_27_47# net206 0
C23551 net188 _0187_ 0
C23552 _0209_ clknet_0__0463_ 0
C23553 hold34/a_49_47# acc0.A\[11\] 0
C23554 _0648_/a_27_297# _0279_ 0.05771f
C23555 _0577_/a_373_47# net48 0
C23556 hold17/a_49_47# _0480_ 0
C23557 _0547_/a_68_297# net127 0.0045f
C23558 clknet_1_1__leaf__0460_ _0317_ 0.06207f
C23559 clknet_1_0__leaf__0465_ hold7/a_391_47# 0.01146f
C23560 _1017_/a_1059_315# _0218_ 0
C23561 _1072_/a_27_47# control0.count\[2\] 0
C23562 hold48/a_49_47# VPWR 0.35889f
C23563 _0237_ hold94/a_49_47# 0.00657f
C23564 VPWR _0790_/a_117_297# 0.00872f
C23565 net62 net74 0
C23566 _0958_/a_27_47# net17 0
C23567 _0691_/a_68_297# clknet_0__0460_ 0.03981f
C23568 _1002_/a_193_47# clknet_1_0__leaf__0460_ 0.00988f
C23569 net126 _1041_/a_381_47# 0
C23570 _0294_ net146 0.15485f
C23571 _1006_/a_466_413# _0219_ 0
C23572 _0086_ net47 0
C23573 _0221_ _0702_/a_113_47# 0
C23574 _0174_ _0206_ 0.14544f
C23575 output39/a_27_47# A[13] 0
C23576 _0800_/a_240_47# net81 0.00278f
C23577 hold87/a_285_47# _0346_ 0
C23578 hold41/a_285_47# acc0.A\[11\] 0.04863f
C23579 _0467_ _1068_/a_891_413# 0
C23580 _0518_/a_27_297# _0518_/a_373_47# 0.01338f
C23581 _0183_ _0225_ 0
C23582 hold83/a_49_47# hold83/a_285_47# 0.22264f
C23583 _0985_/a_193_47# _0985_/a_891_413# 0.19489f
C23584 _0985_/a_27_47# _0985_/a_381_47# 0.06222f
C23585 _0985_/a_634_159# _0985_/a_1059_315# 0
C23586 _0295_ acc0.A\[9\] 0
C23587 _0217_ hold29/a_49_47# 0
C23588 hold46/a_391_47# comp0.B\[14\] 0.06027f
C23589 _0217_ _0566_/a_27_47# 0.00135f
C23590 hold38/a_49_47# comp0.B\[2\] 0
C23591 _0973_/a_109_297# net17 0.00194f
C23592 _0780_/a_285_47# _0397_ 0.00283f
C23593 _0998_/a_27_47# _0181_ 0
C23594 _1018_/a_27_47# _1018_/a_1059_315# 0.04875f
C23595 _1018_/a_193_47# _1018_/a_466_413# 0.07482f
C23596 _0086_ _0831_/a_285_47# 0
C23597 net70 _0399_ 0
C23598 control0.count\[2\] _1071_/a_592_47# 0.00258f
C23599 net46 _0122_ 0
C23600 _0404_ _0670_/a_215_47# 0
C23601 net50 _1022_/a_466_413# 0
C23602 hold28/a_49_47# clkbuf_1_0__f__0464_/a_110_47# 0.00152f
C23603 output47/a_27_47# clknet_1_1__leaf__0465_ 0.0065f
C23604 net61 _0186_ 0.13374f
C23605 _0818_/a_193_47# clknet_0__0465_ 0
C23606 _0982_/a_27_47# _0982_/a_193_47# 0.96469f
C23607 net160 control0.sh 0.27029f
C23608 _0353_ _0707_/a_208_47# 0
C23609 _1010_/a_1059_315# acc0.A\[29\] 0.00177f
C23610 B[11] net18 0.00164f
C23611 _0983_/a_27_47# acc0.A\[15\] 0.00282f
C23612 clknet_1_1__leaf_clk _0951_/a_209_311# 0.01484f
C23613 _0216_ acc0.A\[18\] 0.12352f
C23614 _0348_ VPWR 0.51574f
C23615 _0228_ net91 0.06932f
C23616 net45 net43 0.10231f
C23617 net221 net219 0.01782f
C23618 _0645_/a_47_47# _0671_/a_113_297# 0
C23619 _1019_/a_891_413# _0459_ 0
C23620 _0359_ _1007_/a_1017_47# 0
C23621 hold99/a_285_47# VPWR 0.31752f
C23622 _0753_/a_297_297# _0343_ 0.06718f
C23623 _0130_ clknet_1_0__leaf__0461_ 0.29231f
C23624 _0530_/a_81_21# _0197_ 0.16587f
C23625 hold44/a_391_47# _0195_ 0
C23626 hold44/a_49_47# _0216_ 0.00622f
C23627 _0780_/a_285_297# acc0.A\[17\] 0
C23628 _0397_ _0677_/a_47_47# 0
C23629 _0276_ _0669_/a_111_297# 0.00357f
C23630 _1054_/a_193_47# input15/a_75_212# 0
C23631 _1019_/a_27_47# _0586_/a_27_47# 0
C23632 VPWR _1027_/a_975_413# 0.00497f
C23633 hold98/a_49_47# hold98/a_285_47# 0.22264f
C23634 hold79/a_285_47# hold79/a_391_47# 0.41909f
C23635 _0369_ _0673_/a_253_47# 0.00249f
C23636 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# 1.62775f
C23637 _0473_ _1045_/a_27_47# 0
C23638 VPWR _0749_/a_384_47# 0
C23639 _0693_/a_68_297# _0315_ 0
C23640 net89 _0760_/a_129_47# 0
C23641 net45 _0999_/a_27_47# 0.01203f
C23642 VPWR _1052_/a_193_47# 0.29982f
C23643 _0339_ net208 0.02745f
C23644 _1023_/a_193_47# _1022_/a_27_47# 0
C23645 _1023_/a_27_47# _1022_/a_193_47# 0.00785f
C23646 _1056_/a_1059_315# acc0.A\[10\] 0.10631f
C23647 net8 _1040_/a_27_47# 0
C23648 _0459_ net206 0.02224f
C23649 clk _0485_ 0.03115f
C23650 _0251_ acc0.A\[8\] 0.1753f
C23651 _0174_ _1046_/a_1059_315# 0
C23652 acc0.A\[25\] _1008_/a_1059_315# 0
C23653 hold100/a_49_47# _0446_ 0.0072f
C23654 _0134_ _1036_/a_27_47# 0
C23655 hold3/a_285_47# _0460_ 0
C23656 _0743_/a_240_47# _0360_ 0.03602f
C23657 net152 _1040_/a_193_47# 0
C23658 net32 _1040_/a_27_47# 0
C23659 _0487_ _1063_/a_1059_315# 0.00315f
C23660 clknet_0__0459_ _0183_ 0.02155f
C23661 _0342_ _0219_ 0.07067f
C23662 clkbuf_1_1__f__0464_/a_110_47# _1045_/a_27_47# 0
C23663 clkbuf_0__0460_/a_110_47# _0743_/a_149_47# 0
C23664 clknet_1_0__leaf__0465_ clknet_1_1__leaf__0458_ 0.14208f
C23665 hold58/a_285_47# comp0.B\[3\] 0.00296f
C23666 net55 _0358_ 0.1086f
C23667 acc0.A\[8\] _0989_/a_592_47# 0.00281f
C23668 _0233_ _0374_ 0
C23669 _0155_ _0187_ 0
C23670 VPWR _0332_ 0.54987f
C23671 _0804_/a_79_21# _0279_ 0.08081f
C23672 _0416_ _0648_/a_27_297# 0
C23673 pp[17] net162 0.00329f
C23674 _0346_ _0991_/a_561_413# 0.0015f
C23675 net159 _0487_ 0.20616f
C23676 _0994_/a_891_413# net80 0
C23677 hold78/a_391_47# _0340_ 0
C23678 clknet_1_0__leaf__0464_ _0987_/a_561_413# 0
C23679 _0544_/a_149_47# net198 0.00653f
C23680 _0544_/a_512_297# net18 0
C23681 _0811_/a_81_21# net37 0
C23682 _0345_ _0321_ 0.1085f
C23683 acc0.A\[31\] VPWR 0.83913f
C23684 VPWR _0685_/a_68_297# 0.17071f
C23685 pp[15] _0341_ 0
C23686 _0357_ _0347_ 0.29608f
C23687 _0519_/a_299_297# _0989_/a_27_47# 0
C23688 clkbuf_0__0460_/a_110_47# _0345_ 0
C23689 net43 _0587_/a_27_47# 0
C23690 _0334_ _0219_ 0.02352f
C23691 VPWR net12 0.72292f
C23692 _1034_/a_1059_315# _1034_/a_1017_47# 0
C23693 _0536_/a_51_297# _0144_ 0.10228f
C23694 _0513_/a_384_47# acc0.A\[11\] 0
C23695 hold6/a_49_47# _0204_ 0
C23696 net238 _0410_ 0.1534f
C23697 output65/a_27_47# _0989_/a_27_47# 0
C23698 _0343_ _0507_/a_109_47# 0
C23699 net168 net139 0
C23700 input25/a_75_212# net27 0.14375f
C23701 net25 input27/a_75_212# 0
C23702 _0440_ _0834_/a_109_297# 0.01129f
C23703 net58 acc0.A\[8\] 0.02374f
C23704 hold6/a_49_47# hold6/a_391_47# 0.00188f
C23705 clknet_1_1__leaf__0460_ net197 0
C23706 acc0.A\[23\] _1006_/a_193_47# 0
C23707 _0728_/a_59_75# _0334_ 0
C23708 clkbuf_0__0464_/a_110_47# _1044_/a_27_47# 0
C23709 _0640_/a_465_297# clknet_0__0465_ 0
C23710 _0627_/a_369_297# VPWR 0
C23711 _0499_/a_145_75# _0178_ 0
C23712 hold85/a_49_47# _0477_ 0.0135f
C23713 _1013_/a_592_47# _0219_ 0
C23714 _0190_ acc0.A\[9\] 0
C23715 _0999_/a_27_47# _0587_/a_27_47# 0
C23716 _0570_/a_27_297# _0126_ 0.10883f
C23717 _0570_/a_373_47# net190 0.00265f
C23718 clknet_0__0464_ _1045_/a_561_413# 0
C23719 _0534_/a_81_21# _1047_/a_27_47# 0.00171f
C23720 hold10/a_391_47# _0176_ 0
C23721 _0481_ hold79/a_285_47# 0.00839f
C23722 _0179_ _0289_ 0.46952f
C23723 clknet_1_0__leaf__0459_ _0580_/a_27_297# 0
C23724 net163 _0340_ 0
C23725 comp0.B\[14\] net153 0
C23726 net149 _0178_ 0.00537f
C23727 net36 _0856_/a_79_21# 0
C23728 _0446_ _0450_ 0.28875f
C23729 _0848_/a_27_47# _0451_ 0.052f
C23730 net206 _0265_ 0.01743f
C23731 net243 net50 0.45872f
C23732 _0344_ _1013_/a_466_413# 0
C23733 VPWR _0817_/a_585_47# 0
C23734 pp[30] _1031_/a_193_47# 0.00266f
C23735 _1001_/a_634_159# _0352_ 0
C23736 _0793_/a_240_47# net42 0.09349f
C23737 _1058_/a_27_47# net2 0
C23738 _0218_ _0451_ 0.03289f
C23739 _1058_/a_1059_315# A[11] 0
C23740 _0626_/a_68_297# _0432_ 0
C23741 clknet_0__0459_ acc0.A\[15\] 0.16072f
C23742 pp[15] _1013_/a_891_413# 0.0012f
C23743 clknet_0_clk _0972_/a_250_297# 0
C23744 net180 _0159_ 0
C23745 _0232_ net52 0
C23746 _1050_/a_27_47# _0270_ 0
C23747 _1018_/a_891_413# _0242_ 0
C23748 _0080_ _0265_ 0
C23749 _1071_/a_1059_315# _0466_ 0.003f
C23750 _1071_/a_891_413# _0488_ 0
C23751 net21 input21/a_75_212# 0.10848f
C23752 _0993_/a_466_413# _0286_ 0
C23753 net81 _0995_/a_466_413# 0
C23754 hold77/a_391_47# _1009_/a_193_47# 0
C23755 hold8/a_391_47# _0352_ 0
C23756 clknet_1_0__leaf__0460_ _1005_/a_1017_47# 0
C23757 _0476_ _1062_/a_27_47# 0.00109f
C23758 _1017_/a_466_413# _1017_/a_592_47# 0.00553f
C23759 _1017_/a_634_159# _1017_/a_1017_47# 0
C23760 _0343_ _0242_ 0.05593f
C23761 _0353_ acc0.A\[30\] 0
C23762 _0487_ _1062_/a_975_413# 0
C23763 net211 _0216_ 0.04224f
C23764 _1058_/a_193_47# net3 0
C23765 _0753_/a_465_47# _0375_ 0.00141f
C23766 _0231_ _0752_/a_27_413# 0
C23767 _0753_/a_297_297# _0376_ 0.00565f
C23768 _0723_/a_207_413# hold80/a_391_47# 0.00121f
C23769 net64 _0251_ 0.02793f
C23770 control0.sh acc0.A\[15\] 0
C23771 _1052_/a_381_47# net9 0.01915f
C23772 _0786_/a_217_297# _0422_ 0.00111f
C23773 hold24/a_391_47# _0137_ 0
C23774 net10 _1040_/a_27_47# 0
C23775 _0473_ net132 0.0018f
C23776 _0361_ clknet_0__0460_ 0.02632f
C23777 _0126_ hold50/a_49_47# 0.00838f
C23778 clknet_0__0458_ acc0.A\[6\] 0.0104f
C23779 _0507_/a_109_297# net5 0.00987f
C23780 _1000_/a_1059_315# net45 0.1295f
C23781 _1056_/a_891_413# hold34/a_391_47# 0
C23782 _0172_ A[15] 0
C23783 net137 net11 0
C23784 _0514_/a_27_297# _0186_ 0.12572f
C23785 _0804_/a_79_21# _0416_ 0.10798f
C23786 _0804_/a_297_297# _0415_ 0.00314f
C23787 _0254_ clkbuf_1_1__f__0458_/a_110_47# 0.02221f
C23788 net204 _0553_/a_149_47# 0
C23789 _0555_/a_240_47# _0174_ 0
C23790 _0402_ net228 0.01833f
C23791 _0714_/a_51_297# _0220_ 0
C23792 _0476_ _0561_/a_51_297# 0.08179f
C23793 _0521_/a_299_297# _0521_/a_384_47# 0
C23794 _1033_/a_634_159# _1033_/a_1059_315# 0
C23795 _1033_/a_27_47# _1033_/a_381_47# 0.05761f
C23796 _1033_/a_193_47# _1033_/a_891_413# 0.19685f
C23797 _0457_ _0956_/a_32_297# 0
C23798 _0655_/a_109_93# acc0.A\[15\] 0
C23799 _0329_ net97 0
C23800 _0259_ _0659_/a_150_297# 0.00149f
C23801 _0985_/a_381_47# _0197_ 0
C23802 VPWR _0951_/a_296_53# 0
C23803 _0758_/a_79_21# net51 0
C23804 _1012_/a_634_159# _1012_/a_1059_315# 0
C23805 _1012_/a_27_47# _1012_/a_381_47# 0.06222f
C23806 _1012_/a_193_47# _1012_/a_891_413# 0.19685f
C23807 _0196_ _0527_/a_109_297# 0.00859f
C23808 _0293_ _0424_ 0.16549f
C23809 _0401_ _0992_/a_561_413# 0
C23810 _0758_/a_215_47# net93 0
C23811 _0352_ _1007_/a_381_47# 0
C23812 _1056_/a_1059_315# _0510_/a_109_297# 0
C23813 _0260_ _0399_ 0
C23814 _0512_/a_109_297# _0186_ 0.01116f
C23815 _0216_ _1031_/a_891_413# 0
C23816 _0107_ _1009_/a_634_159# 0.00165f
C23817 _0399_ _0795_/a_384_47# 0
C23818 _0233_ _0249_ 0
C23819 net64 net58 0.41482f
C23820 VPWR acc0.A\[10\] 1.05307f
C23821 net58 _0621_/a_117_297# 0
C23822 _1002_/a_27_47# hold93/a_49_47# 0
C23823 VPWR _0738_/a_68_297# 0.15249f
C23824 _1072_/a_975_413# clknet_0_clk 0
C23825 _1050_/a_193_47# net136 0.01325f
C23826 _1050_/a_1059_315# _1050_/a_1017_47# 0
C23827 _0274_ VPWR 0.48309f
C23828 _0305_ _0996_/a_27_47# 0
C23829 _0476_ _0133_ 0.02379f
C23830 _0343_ _1030_/a_27_47# 0.02143f
C23831 _0990_/a_891_413# _0181_ 0.01453f
C23832 hold31/a_49_47# _0399_ 0
C23833 net36 _0454_ 0.00224f
C23834 _0325_ _0460_ 0.0138f
C23835 hold26/a_49_47# _0540_/a_51_297# 0
C23836 _1041_/a_891_413# _0546_/a_51_297# 0
C23837 _1041_/a_193_47# _0546_/a_240_47# 0
C23838 net132 _0186_ 0
C23839 _1024_/a_381_47# net50 0.00567f
C23840 clknet_1_0__leaf__0464_ _1051_/a_1059_315# 0
C23841 _0221_ net97 0.17809f
C23842 _0179_ acc0.A\[3\] 0.18038f
C23843 input10/a_75_212# net10 0.10863f
C23844 VPWR _0837_/a_266_47# 0.01827f
C23845 _0149_ hold7/a_285_47# 0
C23846 _0764_/a_299_297# _0462_ 0.00643f
C23847 clkbuf_1_0__f__0463_/a_110_47# _0549_/a_68_297# 0
C23848 _0218_ _0373_ 0
C23849 _0565_/a_51_297# net201 0.08461f
C23850 hold11/a_285_47# hold26/a_49_47# 0
C23851 comp0.B\[0\] _0171_ 0.00423f
C23852 _0730_/a_79_21# _0350_ 0.00288f
C23853 _0231_ clknet_1_1__leaf__0460_ 0
C23854 net157 acc0.A\[15\] 0.33608f
C23855 _0544_/a_51_297# _1043_/a_193_47# 0
C23856 _0461_ _0388_ 0.00448f
C23857 acc0.A\[21\] _0227_ 0.11461f
C23858 _0369_ _0830_/a_79_21# 0.10514f
C23859 _0998_/a_1017_47# net43 0
C23860 _0762_/a_79_21# clknet_1_0__leaf__0460_ 0.00338f
C23861 _0229_ net51 0.01207f
C23862 _1017_/a_27_47# net219 0
C23863 _1054_/a_381_47# _1052_/a_891_413# 0
C23864 _0181_ clknet_1_1__leaf_clk 0
C23865 net76 clknet_1_1__leaf__0458_ 0.10241f
C23866 acc0.A\[27\] _0322_ 0.12005f
C23867 hold65/a_285_47# _0828_/a_113_297# 0
C23868 _0252_ _0180_ 0
C23869 _1014_/a_891_413# hold2/a_49_47# 0
C23870 _0179_ _1054_/a_1059_315# 0.08092f
C23871 net21 _1044_/a_1059_315# 0
C23872 _0143_ _1044_/a_193_47# 0
C23873 acc0.A\[27\] _0327_ 0.02707f
C23874 _0343_ _0153_ 0
C23875 acc0.A\[14\] _0158_ 0.02646f
C23876 clkbuf_0__0463_/a_110_47# _0953_/a_32_297# 0
C23877 _0182_ control0.reset 0.00236f
C23878 net56 _0338_ 0
C23879 _0098_ _1018_/a_1059_315# 0
C23880 net45 _1018_/a_193_47# 0
C23881 _0719_/a_27_47# _0238_ 0
C23882 _0357_ hold95/a_49_47# 0
C23883 output59/a_27_47# _0219_ 0.00333f
C23884 _1056_/a_891_413# _0181_ 0
C23885 _0486_ _0166_ 0.07024f
C23886 _0143_ net131 0
C23887 _1031_/a_193_47# _0339_ 0.03407f
C23888 _0750_/a_181_47# _0373_ 0.00168f
C23889 net205 _1036_/a_891_413# 0
C23890 _1020_/a_27_47# clknet_0__0457_ 0
C23891 _0973_/a_109_297# _0165_ 0.00498f
C23892 _0555_/a_240_47# _0208_ 0.09042f
C23893 _0238_ _0460_ 0.04728f
C23894 _1024_/a_27_47# _1023_/a_1059_315# 0
C23895 _0820_/a_297_297# _0369_ 0
C23896 _0256_ _0638_/a_109_297# 0
C23897 comp0.B\[13\] _1046_/a_1059_315# 0.02763f
C23898 net193 _1046_/a_634_159# 0
C23899 acc0.A\[29\] _0700_/a_113_47# 0
C23900 VPWR pp[5] 0.53724f
C23901 acc0.A\[1\] _0465_ 0.07764f
C23902 net234 _0181_ 0.15541f
C23903 _0182_ _1061_/a_891_413# 0
C23904 net8 _1061_/a_466_413# 0
C23905 _0180_ _1061_/a_1059_315# 0
C23906 _0343_ net86 0
C23907 net119 _0173_ 0.00982f
C23908 _0131_ _0213_ 0.00234f
C23909 _0445_ _0840_/a_68_297# 0.10566f
C23910 comp0.B\[15\] _1047_/a_193_47# 0
C23911 _1012_/a_891_413# clknet_1_1__leaf__0461_ 0
C23912 _1012_/a_466_413# net98 0
C23913 clkbuf_0__0460_/a_110_47# net52 0.00396f
C23914 _1046_/a_634_159# _1046_/a_466_413# 0.23992f
C23915 _1046_/a_193_47# _1046_/a_1059_315# 0.03138f
C23916 _1046_/a_27_47# _1046_/a_891_413# 0.03024f
C23917 net39 _0414_ 0.31148f
C23918 pp[30] _0712_/a_297_297# 0
C23919 _0978_/a_109_47# _0466_ 0.00309f
C23920 _0475_ _0956_/a_32_297# 0.36842f
C23921 net40 acc0.A\[13\] 0.67094f
C23922 _1058_/a_1059_315# net66 0
C23923 _1019_/a_891_413# _0772_/a_79_21# 0
C23924 acc0.A\[21\] _0759_/a_113_47# 0
C23925 clknet_1_1__leaf__0463_ net24 0.00203f
C23926 clknet_1_0__leaf__0462_ net51 0.03475f
C23927 _0271_ _0218_ 0.1536f
C23928 net54 _0570_/a_27_297# 0.0031f
C23929 _0716_/a_27_47# clknet_1_1__leaf__0459_ 0
C23930 net8 net171 0.38998f
C23931 acc0.A\[2\] acc0.A\[1\] 0
C23932 _1032_/a_466_413# clknet_1_0__leaf__0457_ 0.00209f
C23933 _1016_/a_975_413# net221 0.00176f
C23934 _1016_/a_466_413# _0115_ 0.00682f
C23935 net166 _0582_/a_27_297# 0
C23936 _0432_ _0252_ 0
C23937 _0234_ _0375_ 0.0098f
C23938 _0221_ _0707_/a_201_297# 0.0376f
C23939 net215 _1024_/a_891_413# 0
C23940 _1051_/a_27_47# _1050_/a_27_47# 0
C23941 _0322_ _0364_ 0.00151f
C23942 VPWR _0117_ 0.2188f
C23943 _0207_ net152 0
C23944 net178 acc0.A\[6\] 0.01049f
C23945 _0724_/a_113_297# _0219_ 0.00241f
C23946 VPWR _0203_ 0.32069f
C23947 _0775_/a_510_47# _0393_ 0.00189f
C23948 pp[8] net2 0.00107f
C23949 _0996_/a_891_413# net42 0.01001f
C23950 _0996_/a_1059_315# acc0.A\[15\] 0.03105f
C23951 net123 _1038_/a_27_47# 0
C23952 clknet_1_0__leaf__0463_ _1038_/a_634_159# 0.00114f
C23953 VPWR net43 0.98581f
C23954 _0172_ comp0.B\[12\] 0.08054f
C23955 hold64/a_285_47# acc0.A\[18\] 0
C23956 _0211_ _1036_/a_1059_315# 0
C23957 hold33/a_285_47# net180 0.01509f
C23958 acc0.A\[12\] hold42/a_285_47# 0.00139f
C23959 net196 _0542_/a_51_297# 0.0591f
C23960 hold38/a_285_47# _0215_ 0
C23961 _0186_ _0431_ 0
C23962 VPWR _0701_/a_209_47# 0
C23963 acc0.A\[12\] _1057_/a_1059_315# 0.05262f
C23964 _0998_/a_27_47# clknet_1_1__leaf__0461_ 0.00264f
C23965 _0662_/a_299_297# _0423_ 0.00414f
C23966 _0662_/a_81_21# _0290_ 0.04037f
C23967 hold27/a_391_47# _0472_ 0.00199f
C23968 _0723_/a_207_413# _0336_ 0
C23969 _0328_ _0370_ 0
C23970 VPWR hold73/a_285_47# 0.28743f
C23971 clkload1/a_110_47# net248 0
C23972 clkload1/Y hold101/a_285_47# 0
C23973 _1016_/a_1017_47# _0459_ 0
C23974 _0457_ _1032_/a_193_47# 0.01767f
C23975 _0279_ _0280_ 0
C23976 _0179_ net157 0
C23977 net44 _0999_/a_1059_315# 0.08557f
C23978 net59 hold16/a_285_47# 0.00265f
C23979 _0230_ _0750_/a_27_47# 0
C23980 _0226_ _0750_/a_109_47# 0.00231f
C23981 _0206_ comp0.B\[9\] 0.0372f
C23982 clkbuf_1_1__f__0460_/a_110_47# acc0.A\[29\] 0.00123f
C23983 hold54/a_49_47# net23 0.01271f
C23984 net168 acc0.A\[8\] 0
C23985 _0261_ _0350_ 0.04417f
C23986 _0181_ _0584_/a_109_47# 0.00324f
C23987 _1016_/a_27_47# _0218_ 0
C23988 _0294_ _1016_/a_193_47# 0
C23989 VPWR _0999_/a_27_47# 0.61606f
C23990 hold37/a_391_47# comp0.B\[14\] 0.0015f
C23991 hold27/a_49_47# _0536_/a_51_297# 0
C23992 _0667_/a_113_47# _0297_ 0
C23993 _0477_ net17 0.02447f
C23994 _0459_ _0773_/a_35_297# 0
C23995 hold20/a_49_47# _0487_ 0
C23996 net162 _0567_/a_109_297# 0.01052f
C23997 clknet_0__0459_ _0645_/a_129_47# 0.00222f
C23998 net45 _0708_/a_68_297# 0.0011f
C23999 _0598_/a_297_47# _0227_ 0.05465f
C24000 comp0.B\[2\] _0565_/a_51_297# 0
C24001 net61 net62 0.0271f
C24002 _0243_ _0311_ 0
C24003 _0518_/a_373_47# _0191_ 0.00217f
C24004 net61 _0450_ 0
C24005 net4 acc0.A\[11\] 0.1786f
C24006 _1038_/a_891_413# clknet_0__0463_ 0
C24007 _1039_/a_466_413# net8 0.01294f
C24008 _0985_/a_466_413# _0083_ 0.02202f
C24009 _0195_ _0728_/a_145_75# 0
C24010 net186 comp0.B\[6\] 0
C24011 pp[28] hold16/a_391_47# 0
C24012 clkbuf_1_0__f__0463_/a_110_47# _1040_/a_891_413# 0.01835f
C24013 VPWR _0510_/a_109_297# 0.19199f
C24014 _0464_ _0138_ 0
C24015 _1018_/a_891_413# _1018_/a_1017_47# 0.00617f
C24016 _1018_/a_634_159# net104 0
C24017 hold67/a_285_47# clknet_1_1__leaf__0465_ 0.04545f
C24018 _0343_ _0990_/a_27_47# 0.02624f
C24019 comp0.B\[14\] _1046_/a_592_47# 0
C24020 clkbuf_0__0461_/a_110_47# _0675_/a_68_297# 0.01049f
C24021 net50 net151 0.00142f
C24022 _0970_/a_27_297# _0484_ 0.18701f
C24023 _0789_/a_315_47# _0409_ 0.00146f
C24024 _0795_/a_81_21# _0345_ 0.00248f
C24025 _1053_/a_27_47# net15 0
C24026 _0982_/a_634_159# _0982_/a_1017_47# 0
C24027 _0982_/a_466_413# _0982_/a_592_47# 0.00553f
C24028 VPWR _0368_ 0.38976f
C24029 hold88/a_391_47# _0833_/a_79_21# 0
C24030 _1011_/a_381_47# clknet_1_1__leaf__0462_ 0
C24031 _1049_/a_634_159# _1049_/a_592_47# 0
C24032 _0157_ _0346_ 0
C24033 _0457_ _0721_/a_27_47# 0.02482f
C24034 _0869_/a_27_47# clkbuf_1_0__f__0461_/a_110_47# 0.01201f
C24035 hold65/a_285_47# _0433_ 0.00296f
C24036 _0304_ _0302_ 0
C24037 _0240_ _0219_ 0.00476f
C24038 net66 net47 0
C24039 pp[10] A[11] 0.58018f
C24040 net39 _0300_ 0.00519f
C24041 _0747_/a_79_21# _0747_/a_510_47# 0.00844f
C24042 _0747_/a_297_297# _0747_/a_215_47# 0
C24043 _0233_ _0231_ 0.41304f
C24044 net48 hold73/a_285_47# 0.08915f
C24045 control0.count\[3\] control0.state\[2\] 0
C24046 _0369_ _0219_ 0.25722f
C24047 VPWR _0618_/a_215_47# 0.00164f
C24048 net10 _1061_/a_466_413# 0
C24049 _1052_/a_193_47# _0523_/a_81_21# 0.00297f
C24050 _0339_ _0395_ 0
C24051 _1053_/a_27_47# _1053_/a_1059_315# 0.04875f
C24052 _1053_/a_193_47# _1053_/a_466_413# 0.08301f
C24053 _0575_/a_27_297# _0575_/a_373_47# 0.01338f
C24054 _0637_/a_139_47# _0267_ 0
C24055 _0269_ _0635_/a_109_297# 0
C24056 _0093_ net6 0
C24057 _0714_/a_245_297# _0218_ 0
C24058 _1019_/a_381_47# _0218_ 0
C24059 clknet_1_1__leaf__0462_ acc0.A\[25\] 0.01833f
C24060 net40 net245 0.00397f
C24061 _0195_ _1008_/a_466_413# 0
C24062 _0996_/a_27_47# _0181_ 0
C24063 hold39/a_391_47# _1065_/a_193_47# 0
C24064 _0748_/a_81_21# _0326_ 0
C24065 _0129_ _0195_ 0.0777f
C24066 _1066_/a_634_159# _1066_/a_592_47# 0
C24067 _0627_/a_109_93# acc0.A\[6\] 0.00191f
C24068 _0831_/a_285_297# acc0.A\[8\] 0
C24069 _0338_ _0345_ 0
C24070 _1046_/a_1059_315# comp0.B\[9\] 0.00221f
C24071 _0441_ acc0.A\[3\] 0
C24072 _0327_ _1010_/a_193_47# 0
C24073 _0991_/a_27_47# net47 0.03381f
C24074 hold34/a_49_47# A[12] 0
C24075 _0849_/a_510_47# _0263_ 0
C24076 control0.reset _0562_/a_150_297# 0
C24077 _1034_/a_27_47# _0175_ 0.03308f
C24078 _1056_/a_27_47# _0343_ 0
C24079 _0201_ _1042_/a_634_159# 0
C24080 net31 _1040_/a_634_159# 0
C24081 _0680_/a_472_297# _0462_ 0.00163f
C24082 _1068_/a_634_159# _1068_/a_592_47# 0
C24083 acc0.A\[23\] _0103_ 0
C24084 _0222_ hold94/a_49_47# 0.00178f
C24085 _1030_/a_634_159# _1030_/a_1059_315# 0
C24086 _1030_/a_27_47# _1030_/a_381_47# 0.06222f
C24087 _1030_/a_193_47# _1030_/a_891_413# 0.19226f
C24088 _0254_ _0291_ 0
C24089 _1041_/a_634_159# _0176_ 0
C24090 _0712_/a_297_297# _0339_ 0.03958f
C24091 net207 _0782_/a_27_47# 0
C24092 net71 _0447_ 0
C24093 clkbuf_1_1__f__0465_/a_110_47# _0817_/a_81_21# 0
C24094 _0283_ acc0.A\[10\] 0.09131f
C24095 _1017_/a_27_47# _0352_ 0
C24096 _1034_/a_193_47# control0.sh 0
C24097 hold41/a_285_47# A[12] 0
C24098 net205 _0474_ 0
C24099 _0476_ _0959_/a_300_47# 0.00152f
C24100 _0183_ _0462_ 0
C24101 _0752_/a_27_413# _0225_ 0
C24102 _0330_ _0726_/a_512_297# 0
C24103 pp[9] net3 0.17445f
C24104 _0416_ _0280_ 0
C24105 hold9/a_285_47# hold9/a_391_47# 0.41909f
C24106 _0429_ _0519_/a_299_297# 0
C24107 _0312_ _1009_/a_381_47# 0
C24108 _0571_/a_27_297# clknet_1_1__leaf__0462_ 0.00102f
C24109 _1035_/a_381_47# clknet_1_1__leaf__0463_ 0.00322f
C24110 _1035_/a_1059_315# net122 0
C24111 _0753_/a_381_47# net46 0
C24112 _0992_/a_634_159# net37 0
C24113 _0804_/a_297_297# _0347_ 0.00165f
C24114 _0786_/a_217_297# _0423_ 0
C24115 _0786_/a_80_21# _0290_ 0
C24116 _0216_ _0611_/a_150_297# 0
C24117 _0429_ output65/a_27_47# 0
C24118 net18 _0140_ 0
C24119 _0110_ _0306_ 0
C24120 _0598_/a_79_21# _0229_ 0.15394f
C24121 _1015_/a_1059_315# _0181_ 0.01079f
C24122 _0320_ _0737_/a_35_297# 0.01996f
C24123 _0987_/a_193_47# _0987_/a_634_159# 0.11897f
C24124 _0987_/a_27_47# _0987_/a_466_413# 0.27314f
C24125 _0152_ acc0.A\[7\] 0.12434f
C24126 _0217_ net102 0
C24127 hold64/a_285_47# net211 0.01139f
C24128 _0946_/a_30_53# _0946_/a_184_297# 0.00863f
C24129 net47 _0350_ 0.23411f
C24130 _1034_/a_975_413# comp0.B\[2\] 0.00186f
C24131 net194 _1045_/a_193_47# 0.01021f
C24132 net220 _0346_ 0
C24133 acc0.A\[27\] _1008_/a_561_413# 0
C24134 clknet_0_clk _0971_/a_81_21# 0
C24135 _0992_/a_1059_315# net67 0.02821f
C24136 _1000_/a_1059_315# VPWR 0.38172f
C24137 VPWR _0188_ 0.15921f
C24138 net40 net45 0
C24139 hold16/a_49_47# _0338_ 0
C24140 net164 _0466_ 0.16185f
C24141 clknet_0__0464_ _1044_/a_381_47# 0
C24142 _1072_/a_381_47# _0466_ 0
C24143 _0151_ _1053_/a_193_47# 0.27429f
C24144 B[12] B[13] 0.28164f
C24145 hold77/a_49_47# net96 0.00128f
C24146 _0750_/a_27_47# _0236_ 0
C24147 _0346_ _1006_/a_592_47# 0
C24148 _0346_ acc0.A\[9\] 0.02599f
C24149 _0378_ net50 0.03093f
C24150 _1029_/a_27_47# _1029_/a_466_413# 0.27314f
C24151 _1029_/a_193_47# _1029_/a_634_159# 0.12729f
C24152 _0304_ net6 0
C24153 _0399_ _0097_ 0
C24154 _0352_ _0772_/a_215_47# 0.06822f
C24155 _0255_ _0445_ 0
C24156 clkbuf_0__0464_/a_110_47# _0196_ 0
C24157 clknet_1_0__leaf__0459_ net43 0.30465f
C24158 _0844_/a_79_21# _0219_ 0.00271f
C24159 _1032_/a_975_413# clknet_1_0__leaf__0461_ 0
C24160 clknet_0_clk _0164_ 0
C24161 net39 _0404_ 0.20256f
C24162 _0387_ _0459_ 0
C24163 net188 clknet_1_1__leaf__0465_ 0.05423f
C24164 _0637_/a_56_297# _0446_ 0
C24165 _0343_ _0998_/a_381_47# 0.0011f
C24166 _0581_/a_373_47# _0393_ 0
C24167 _0722_/a_215_47# clknet_1_1__leaf__0462_ 0
C24168 _0346_ _0670_/a_79_21# 0.00643f
C24169 clkload0/a_27_47# _1072_/a_27_47# 0.00921f
C24170 _0430_ _0831_/a_35_297# 0.0035f
C24171 net64 _0831_/a_285_297# 0
C24172 comp0.B\[13\] _1045_/a_634_159# 0.00233f
C24173 _1050_/a_193_47# net73 0
C24174 _1050_/a_27_47# _0085_ 0
C24175 net136 _0987_/a_193_47# 0
C24176 hold33/a_391_47# hold26/a_49_47# 0
C24177 net99 _0345_ 0.04253f
C24178 _0383_ net109 0
C24179 _1015_/a_193_47# _0565_/a_51_297# 0
C24180 _1015_/a_27_47# _0565_/a_245_297# 0
C24181 clknet_1_0__leaf__0465_ _0536_/a_149_47# 0
C24182 clknet_1_0__leaf__0463_ _0550_/a_149_47# 0.02897f
C24183 pp[30] _0221_ 0
C24184 _0520_/a_373_47# _0180_ 0.00162f
C24185 _1017_/a_1059_315# _1016_/a_1059_315# 0
C24186 _1017_/a_466_413# _1016_/a_891_413# 0
C24187 _0783_/a_79_21# net43 0.00248f
C24188 _0269_ _0186_ 0
C24189 clknet_1_0__leaf__0460_ _0771_/a_215_297# 0
C24190 hold30/a_391_47# net51 0
C24191 _0998_/a_891_413# acc0.A\[17\] 0
C24192 _0254_ _0621_/a_285_297# 0
C24193 net219 _0245_ 0
C24194 B[2] net25 0.00405f
C24195 _0643_/a_253_47# _0255_ 0
C24196 control0.reset _0495_/a_68_297# 0.18859f
C24197 _1037_/a_466_413# clknet_1_1__leaf__0463_ 0
C24198 _0464_ net134 0.02107f
C24199 _1033_/a_193_47# _0956_/a_32_297# 0
C24200 _0998_/a_466_413# clkbuf_1_1__f__0461_/a_110_47# 0.00703f
C24201 _1028_/a_27_47# _1028_/a_634_159# 0.13601f
C24202 _0555_/a_245_297# _0555_/a_240_47# 0
C24203 net201 _0493_/a_27_47# 0
C24204 _0606_/a_109_53# _0373_ 0.02201f
C24205 input4/a_75_212# _0188_ 0
C24206 hold41/a_285_47# _1057_/a_193_47# 0
C24207 clknet_1_0__leaf__0465_ _0218_ 0.12728f
C24208 _0189_ _0186_ 0.01892f
C24209 net44 _0397_ 0.02465f
C24210 net58 _0986_/a_466_413# 0.00544f
C24211 net225 _0220_ 0
C24212 _0476_ _0208_ 0.45161f
C24213 _0999_/a_27_47# _0783_/a_79_21# 0
C24214 _0394_ _1009_/a_27_47# 0
C24215 _0308_ _1009_/a_466_413# 0
C24216 net230 _0151_ 0.48936f
C24217 _1033_/a_27_47# comp0.B\[1\] 0.00149f
C24218 _1033_/a_466_413# _0131_ 0.00337f
C24219 _0985_/a_634_159# VPWR 0.17892f
C24220 net63 _0987_/a_1059_315# 0.11457f
C24221 _0965_/a_129_47# _0478_ 0.00236f
C24222 VPWR _1018_/a_193_47# 0.29698f
C24223 _1039_/a_1017_47# _0176_ 0.00227f
C24224 _0148_ net11 0.23743f
C24225 _0130_ _1033_/a_891_413# 0
C24226 net182 acc0.A\[10\] 0
C24227 _0343_ net44 0.02083f
C24228 _0856_/a_215_47# hold60/a_49_47# 0
C24229 _0846_/a_240_47# _0219_ 0.04681f
C24230 _0985_/a_891_413# _0636_/a_59_75# 0
C24231 _0197_ _0147_ 0.00213f
C24232 _1056_/a_891_413# _0187_ 0
C24233 hold55/a_285_47# hold55/a_391_47# 0.41909f
C24234 net76 _0988_/a_1017_47# 0
C24235 _0243_ _1000_/a_891_413# 0
C24236 _0743_/a_51_297# _0315_ 0
C24237 hold22/a_285_47# _0179_ 0.0073f
C24238 hold4/a_285_47# _1005_/a_891_413# 0
C24239 _1009_/a_561_413# _0219_ 0
C24240 _1050_/a_975_413# acc0.A\[4\] 0
C24241 _0191_ _0987_/a_466_413# 0
C24242 _0981_/a_27_297# _1072_/a_27_47# 0
C24243 hold54/a_391_47# _0457_ 0.00196f
C24244 _1041_/a_466_413# _0139_ 0.00115f
C24245 _0519_/a_299_297# clknet_1_1__leaf__0458_ 0
C24246 acc0.A\[24\] net50 0
C24247 hold37/a_49_47# hold37/a_391_47# 0.00188f
C24248 _0946_/a_30_53# _0162_ 0
C24249 _0946_/a_184_297# _0487_ 0
C24250 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0461_/a_110_47# 0
C24251 _0297_ acc0.A\[15\] 0
C24252 _0508_/a_384_47# net228 0.01f
C24253 _0229_ _0606_/a_297_297# 0
C24254 _0226_ _0606_/a_215_297# 0.00136f
C24255 _0993_/a_466_413# net79 0
C24256 net67 _0421_ 0
C24257 _0517_/a_81_21# _0088_ 0
C24258 VPWR _1034_/a_381_47# 0.06961f
C24259 hold42/a_49_47# _0179_ 0.04063f
C24260 clknet_1_0__leaf__0460_ _1067_/a_1059_315# 0.0942f
C24261 net18 _1043_/a_634_159# 0.00551f
C24262 net198 _1043_/a_466_413# 0.01216f
C24263 VPWR hold6/a_49_47# 0.29425f
C24264 _0155_ clknet_1_1__leaf__0465_ 0.01832f
C24265 _0343_ _0983_/a_634_159# 0.00691f
C24266 clknet_1_0__leaf__0462_ _0324_ 0
C24267 VPWR _0816_/a_68_297# 0.16026f
C24268 _0348_ net56 0.00278f
C24269 _0578_/a_109_297# clknet_1_0__leaf__0457_ 0.0045f
C24270 _0174_ clkbuf_0__0463_/a_110_47# 0.00148f
C24271 _1053_/a_1059_315# A[5] 0
C24272 _0398_ _0309_ 0
C24273 _1002_/a_466_413# acc0.A\[20\] 0
C24274 _0998_/a_193_47# _0998_/a_381_47# 0.09503f
C24275 _0998_/a_634_159# _0998_/a_891_413# 0.03684f
C24276 _0998_/a_27_47# _0998_/a_561_413# 0.00163f
C24277 _0195_ hold61/a_285_47# 0
C24278 _0305_ _0673_/a_103_199# 0.07726f
C24279 net126 _0206_ 0.20542f
C24280 _0779_/a_79_21# _0308_ 0
C24281 _1003_/a_466_413# _0369_ 0
C24282 _0498_/a_149_47# _1061_/a_193_47# 0
C24283 _0498_/a_240_47# _1061_/a_27_47# 0.00129f
C24284 VPWR _0708_/a_68_297# 0.16735f
C24285 net110 _1023_/a_634_159# 0
C24286 _0122_ _1023_/a_193_47# 0
C24287 hold56/a_49_47# _1033_/a_634_159# 0.00115f
C24288 hold56/a_391_47# _1033_/a_27_47# 0.00127f
C24289 hold56/a_285_47# _1033_/a_193_47# 0.00118f
C24290 _0662_/a_81_21# _0986_/a_1059_315# 0
C24291 _0310_ _0308_ 0.09984f
C24292 net169 net75 0
C24293 _0174_ _1044_/a_193_47# 0
C24294 _1019_/a_634_159# _1019_/a_466_413# 0.23992f
C24295 _1019_/a_193_47# _1019_/a_1059_315# 0.03405f
C24296 _1019_/a_27_47# _1019_/a_891_413# 0.03089f
C24297 _0717_/a_80_21# _0221_ 0.10788f
C24298 _1046_/a_466_413# net132 0
C24299 pp[30] _0344_ 0
C24300 hold42/a_49_47# _0513_/a_81_21# 0
C24301 _1000_/a_1059_315# clknet_1_0__leaf__0459_ 0
C24302 hold89/a_49_47# net17 0
C24303 net54 _0126_ 0.02646f
C24304 _1056_/a_381_47# _0153_ 0
C24305 net62 _0431_ 0.02462f
C24306 net123 B[6] 0.0184f
C24307 _0340_ net116 0
C24308 acc0.A\[21\] _0352_ 0.06538f
C24309 clknet_1_1__leaf__0458_ _0986_/a_193_47# 0
C24310 _0837_/a_368_297# _0172_ 0.00134f
C24311 net202 clknet_1_0__leaf__0457_ 0.08415f
C24312 VPWR _1012_/a_634_159# 0.18714f
C24313 net166 _0115_ 0.06397f
C24314 _0221_ _0339_ 0
C24315 _0218_ _0400_ 0
C24316 _0233_ _0225_ 0.2151f
C24317 _1051_/a_891_413# _1050_/a_381_47# 0
C24318 _1051_/a_381_47# _1050_/a_891_413# 0
C24319 _0783_/a_510_47# _0307_ 0.00172f
C24320 _0565_/a_245_297# _0215_ 0.00118f
C24321 hold52/a_285_47# _1024_/a_1059_315# 0
C24322 _0684_/a_145_75# _0316_ 0
C24323 clknet_1_1__leaf__0463_ clknet_1_0__leaf__0457_ 0.00735f
C24324 _0472_ _0496_/a_27_47# 0.02428f
C24325 _0985_/a_1017_47# net175 0
C24326 _1050_/a_27_47# net131 0
C24327 _0642_/a_215_297# clknet_0__0465_ 0
C24328 net56 _0332_ 0.02141f
C24329 net70 _0346_ 0.21468f
C24330 _0902_/a_27_47# hold73/a_49_47# 0.00794f
C24331 clknet_1_0__leaf__0463_ net124 0.19426f
C24332 _0580_/a_27_297# _0345_ 0.01616f
C24333 net9 _1049_/a_1059_315# 0.00625f
C24334 _0292_ _0426_ 0
C24335 net248 _0434_ 0
C24336 clknet_1_1__leaf__0459_ _0998_/a_1059_315# 0.01039f
C24337 control0.sh _0565_/a_240_47# 0
C24338 net160 _0474_ 0.0221f
C24339 _0393_ _0347_ 0.13555f
C24340 hold15/a_391_47# _1031_/a_891_413# 0.00323f
C24341 net162 _1031_/a_27_47# 0.02482f
C24342 _0974_/a_222_93# _0468_ 0.11357f
C24343 clkbuf_0_clk/a_110_47# _0950_/a_75_212# 0.00552f
C24344 hold3/a_285_47# _0373_ 0
C24345 _0982_/a_27_47# net207 0
C24346 net34 clknet_0_clk 0
C24347 _0098_ net46 0
C24348 net101 _0217_ 0
C24349 _0568_/a_109_297# _0333_ 0
C24350 _0758_/a_79_21# _0347_ 0.1323f
C24351 _1024_/a_634_159# pp[24] 0
C24352 _1024_/a_1059_315# net52 0.03101f
C24353 hold32/a_285_47# A[12] 0
C24354 _1052_/a_1017_47# acc0.A\[6\] 0
C24355 _1052_/a_891_413# _0193_ 0
C24356 clknet_0__0458_ _0826_/a_219_297# 0.00945f
C24357 _0294_ _0991_/a_27_47# 0.01203f
C24358 _0984_/a_975_413# _0465_ 0
C24359 _0581_/a_27_297# _0116_ 0.15817f
C24360 _0581_/a_373_47# net206 0.00122f
C24361 _0234_ VPWR 1.39806f
C24362 _0245_ _0352_ 0.14328f
C24363 _0990_/a_634_159# _0990_/a_1059_315# 0
C24364 _0990_/a_27_47# _0990_/a_381_47# 0.05761f
C24365 _0990_/a_193_47# _0990_/a_891_413# 0.18949f
C24366 clkbuf_0__0463_/a_110_47# _0208_ 0.00141f
C24367 _0463_ _0173_ 0
C24368 _0732_/a_303_47# VPWR 0
C24369 _0292_ _0185_ 0
C24370 _0179_ net13 0.03161f
C24371 _0313_ hold90/a_391_47# 0
C24372 net9 net18 0.00158f
C24373 _1002_/a_27_47# clknet_1_0__leaf__0457_ 0.00233f
C24374 _0553_/a_51_297# net8 0
C24375 _0350_ net93 0
C24376 clkbuf_0__0461_/a_110_47# _0242_ 0.02079f
C24377 _0747_/a_297_297# _0352_ 0.00274f
C24378 _0217_ _0228_ 0
C24379 _0985_/a_975_413# acc0.A\[3\] 0
C24380 _0457_ _0182_ 0
C24381 _0967_/a_109_93# _0967_/a_297_297# 0
C24382 _0967_/a_403_297# _0485_ 0.00189f
C24383 _0967_/a_109_93# _0162_ 0
C24384 acc0.A\[25\] _1007_/a_466_413# 0
C24385 _0487_ _0162_ 0.13114f
C24386 _0488_ _0975_/a_59_75# 0.11494f
C24387 hold97/a_49_47# _0329_ 0
C24388 _0409_ _0219_ 0
C24389 clkbuf_1_0__f__0465_/a_110_47# _0270_ 0
C24390 _0805_/a_27_47# _0992_/a_27_47# 0
C24391 hold53/a_391_47# _1025_/a_27_47# 0
C24392 hold53/a_285_47# _1025_/a_193_47# 0.01463f
C24393 net57 clknet_1_1__leaf__0462_ 0
C24394 _1049_/a_891_413# acc0.A\[3\] 0.00342f
C24395 _1034_/a_193_47# _0955_/a_32_297# 0
C24396 VPWR clknet_0__0460_ 2.24212f
C24397 _0273_ clkbuf_1_1__f__0458_/a_110_47# 0
C24398 _1011_/a_1059_315# hold80/a_391_47# 0.01554f
C24399 hold9/a_285_47# _0739_/a_215_47# 0.00236f
C24400 _0848_/a_109_297# _0350_ 0
C24401 clknet_1_0__leaf__0459_ _1018_/a_193_47# 0
C24402 _0461_ _0216_ 0.03441f
C24403 net243 _0576_/a_27_297# 0.00196f
C24404 _0229_ hold3/a_391_47# 0.00106f
C24405 _0226_ hold3/a_49_47# 0.00472f
C24406 net248 _0989_/a_1059_315# 0
C24407 _0294_ _0350_ 0
C24408 _1070_/a_634_159# _1070_/a_592_47# 0
C24409 _1045_/a_27_47# _1045_/a_193_47# 0.97453f
C24410 _0348_ _0345_ 0
C24411 _1052_/a_1059_315# _0150_ 0.00358f
C24412 _1053_/a_891_413# _1053_/a_1017_47# 0.00617f
C24413 net40 VPWR 1.54707f
C24414 pp[17] _1030_/a_1059_315# 0.00284f
C24415 net44 _1030_/a_381_47# 0.02055f
C24416 _1057_/a_592_47# acc0.A\[10\] 0
C24417 clknet_1_0__leaf__0465_ _1050_/a_592_47# 0
C24418 _0198_ _0465_ 0.0064f
C24419 net45 _0998_/a_975_413# 0
C24420 _0577_/a_27_297# net177 0
C24421 _0183_ _1023_/a_891_413# 0
C24422 acc0.A\[22\] _1023_/a_381_47# 0
C24423 _1066_/a_891_413# control0.sh 0.02956f
C24424 hold21/a_285_47# _0518_/a_27_297# 0
C24425 _0584_/a_109_297# net201 0
C24426 _1062_/a_634_159# _0468_ 0
C24427 hold37/a_391_47# acc0.A\[4\] 0
C24428 VPWR _1030_/a_634_159# 0.17634f
C24429 clknet_1_1__leaf__0463_ _0561_/a_149_47# 0.00187f
C24430 _0314_ _1007_/a_592_47# 0
C24431 _1043_/a_27_47# _1043_/a_193_47# 0.96639f
C24432 net7 _1040_/a_634_159# 0
C24433 _0234_ net48 0.06514f
C24434 _0768_/a_27_47# _0308_ 0
C24435 acc0.A\[2\] _0198_ 0.00229f
C24436 _1061_/a_466_413# _0492_/a_27_47# 0
C24437 _1017_/a_193_47# hold72/a_49_47# 0.00957f
C24438 _1017_/a_27_47# hold72/a_285_47# 0
C24439 net109 _1022_/a_1017_47# 0
C24440 _0749_/a_384_47# _0345_ 0
C24441 _0647_/a_47_47# _0303_ 0
C24442 _0997_/a_1059_315# net83 0
C24443 _1038_/a_27_47# _0209_ 0.00331f
C24444 _0344_ _0339_ 0.02018f
C24445 _1030_/a_27_47# _0568_/a_27_297# 0
C24446 hold67/a_49_47# _0399_ 0.00586f
C24447 _1021_/a_193_47# _1002_/a_27_47# 0.0116f
C24448 _1021_/a_27_47# _1002_/a_193_47# 0.00846f
C24449 clknet_1_0__leaf__0462_ _0347_ 0.03555f
C24450 clknet_1_0__leaf__0458_ _1047_/a_193_47# 0
C24451 comp0.B\[7\] _1040_/a_27_47# 0
C24452 _0551_/a_27_47# net17 0
C24453 _0330_ _0109_ 0
C24454 hold27/a_391_47# _1046_/a_891_413# 0
C24455 A[12] net4 0.01914f
C24456 hold100/a_49_47# _0269_ 0.06221f
C24457 _0125_ clknet_1_1__leaf__0462_ 0.04366f
C24458 _1056_/a_634_159# _1056_/a_1059_315# 0
C24459 _1056_/a_27_47# _1056_/a_381_47# 0.06222f
C24460 _1056_/a_193_47# _1056_/a_891_413# 0.19489f
C24461 _1032_/a_891_413# net17 0.02372f
C24462 _0402_ _0401_ 0.01648f
C24463 A[15] _1040_/a_193_47# 0
C24464 net194 _1044_/a_27_47# 0.13501f
C24465 _0947_/a_109_297# _0466_ 0.00217f
C24466 _0332_ _0345_ 0.00692f
C24467 _0987_/a_1059_315# _0987_/a_1017_47# 0
C24468 _0987_/a_193_47# net73 0.01355f
C24469 _0987_/a_27_47# _0085_ 0.09906f
C24470 clknet_1_1__leaf__0459_ _0289_ 0.01234f
C24471 hold74/a_391_47# _0398_ 0
C24472 hold55/a_285_47# _0352_ 0
C24473 pp[17] net45 0.00994f
C24474 _0323_ _0367_ 0
C24475 _0833_/a_79_21# acc0.A\[8\] 0.08416f
C24476 _0348_ hold16/a_49_47# 0
C24477 _0855_/a_299_297# net234 0.05724f
C24478 _0661_/a_205_297# VPWR 0
C24479 _0199_ _1047_/a_466_413# 0.00703f
C24480 _0182_ _1047_/a_561_413# 0.00162f
C24481 _0239_ _0308_ 0
C24482 acc0.A\[31\] _0345_ 0
C24483 _0180_ _0472_ 0
C24484 acc0.A\[20\] _0385_ 0.07411f
C24485 _1041_/a_27_47# _0548_/a_245_297# 0
C24486 clknet_1_0__leaf__0465_ net15 0.00131f
C24487 _1004_/a_634_159# _1004_/a_592_47# 0
C24488 net242 net57 0.05754f
C24489 _0557_/a_149_47# _1035_/a_891_413# 0
C24490 _0557_/a_240_47# _1035_/a_1059_315# 0
C24491 _1027_/a_634_159# _1008_/a_1059_315# 0
C24492 _1027_/a_1059_315# _1008_/a_634_159# 0
C24493 net157 _1049_/a_891_413# 0
C24494 _0403_ _0399_ 0.22455f
C24495 net162 _0712_/a_79_21# 0.02584f
C24496 acc0.A\[31\] _0712_/a_381_47# 0
C24497 _1067_/a_466_413# hold93/a_49_47# 0
C24498 _1067_/a_634_159# hold93/a_285_47# 0
C24499 _1067_/a_193_47# hold93/a_391_47# 0
C24500 comp0.B\[2\] clkbuf_1_1__f_clk/a_110_47# 0
C24501 _0680_/a_472_297# _0312_ 0
C24502 net86 clkbuf_0__0461_/a_110_47# 0.02188f
C24503 clknet_1_0__leaf__0463_ _0464_ 0
C24504 clknet_1_1__leaf__0464_ net154 0.00688f
C24505 _1029_/a_27_47# net191 0.0968f
C24506 _1029_/a_193_47# net115 0.0065f
C24507 _1029_/a_1059_315# _1029_/a_1017_47# 0
C24508 _1019_/a_634_159# _0352_ 0
C24509 input24/a_75_212# net28 0.13421f
C24510 net24 input28/a_75_212# 0
C24511 VPWR net201 0.78471f
C24512 VPWR _0828_/a_113_297# 0.18693f
C24513 comp0.B\[15\] _0178_ 0.04744f
C24514 net62 _0269_ 0.03327f
C24515 comp0.B\[13\] _1044_/a_193_47# 0
C24516 hold69/a_285_47# _0250_ 0
C24517 VPWR _0531_/a_109_297# 0.19582f
C24518 _0269_ _0450_ 0.01104f
C24519 _0268_ _0451_ 0
C24520 _0328_ _0737_/a_285_47# 0
C24521 _0817_/a_585_47# _0345_ 0
C24522 _0260_ _0346_ 0
C24523 _0718_/a_47_47# _0221_ 0
C24524 comp0.B\[13\] net131 0
C24525 acc0.A\[4\] _0987_/a_975_413# 0
C24526 _0216_ _0465_ 0
C24527 _1000_/a_193_47# acc0.A\[18\] 0
C24528 _1004_/a_891_413# _0225_ 0
C24529 _1020_/a_193_47# _0183_ 0.02231f
C24530 _1020_/a_466_413# _0217_ 0
C24531 acc0.A\[16\] _0459_ 0.04991f
C24532 net103 _1016_/a_381_47# 0.00171f
C24533 _0292_ _0289_ 0.11909f
C24534 net206 _0347_ 0
C24535 hold15/a_49_47# _0129_ 0
C24536 net106 net17 0.00324f
C24537 _0382_ net51 0
C24538 _1016_/a_27_47# _1016_/a_1059_315# 0.04672f
C24539 _1016_/a_193_47# _1016_/a_466_413# 0.07482f
C24540 hold101/a_49_47# clknet_1_1__leaf__0458_ 0.00287f
C24541 A[10] net2 0.02802f
C24542 _0343_ _0829_/a_109_297# 0
C24543 _0251_ _0369_ 0.05721f
C24544 hold11/a_285_47# _1061_/a_193_47# 0
C24545 _0135_ clknet_1_1__leaf__0463_ 0
C24546 _0756_/a_129_47# net109 0
C24547 _0512_/a_27_297# net143 0
C24548 _0478_ _0976_/a_505_21# 0
C24549 _1028_/a_891_413# _1028_/a_975_413# 0.00851f
C24550 _1028_/a_27_47# net114 0.22448f
C24551 _1028_/a_381_47# _1028_/a_561_413# 0.00123f
C24552 _0249_ _0617_/a_150_297# 0
C24553 hold25/a_285_47# _1041_/a_27_47# 0
C24554 _0238_ _0373_ 0
C24555 hold17/a_49_47# _1070_/a_27_47# 0
C24556 hold87/a_285_47# _0982_/a_27_47# 0
C24557 _0343_ _0996_/a_381_47# 0
C24558 hold87/a_49_47# _0982_/a_193_47# 0
C24559 _1067_/a_193_47# control0.reset 0
C24560 _0369_ _0989_/a_592_47# 0
C24561 _0440_ _0255_ 0.08254f
C24562 _1057_/a_193_47# net4 0
C24563 clknet_1_0__leaf__0458_ _0265_ 0.01498f
C24564 clknet_0__0459_ clknet_1_1__leaf__0459_ 0.00418f
C24565 _0331_ _0701_/a_80_21# 0
C24566 _0765_/a_510_47# _0460_ 0
C24567 VPWR _0990_/a_634_159# 0.20197f
C24568 _0812_/a_215_47# _0812_/a_510_47# 0.00529f
C24569 _0999_/a_193_47# _0096_ 0
C24570 _0999_/a_634_159# _0399_ 0
C24571 clkbuf_1_1__f__0460_/a_110_47# _0686_/a_219_297# 0
C24572 clkbuf_1_0__f__0462_/a_110_47# _0737_/a_35_297# 0.01336f
C24573 _0245_ _0613_/a_109_297# 0.0124f
C24574 _0514_/a_27_297# _0514_/a_109_297# 0.17136f
C24575 net64 _0833_/a_79_21# 0
C24576 output67/a_27_47# net37 0.02411f
C24577 pp[12] net80 0
C24578 _0557_/a_51_297# _1037_/a_891_413# 0
C24579 VPWR _1049_/a_1017_47# 0
C24580 _0135_ net8 0
C24581 _0473_ _0560_/a_68_297# 0
C24582 _0556_/a_68_297# net24 0.04408f
C24583 net237 _0367_ 0.06078f
C24584 net140 hold83/a_391_47# 0
C24585 _0516_/a_373_47# _0181_ 0.00122f
C24586 _1041_/a_975_413# net31 0
C24587 _1017_/a_193_47# clknet_0__0461_ 0
C24588 _0647_/a_285_47# VPWR 0.00241f
C24589 net20 hold51/a_391_47# 0.05379f
C24590 _0460_ _1006_/a_891_413# 0.01316f
C24591 net120 comp0.B\[6\] 0
C24592 VPWR _1066_/a_1017_47# 0
C24593 net58 _0369_ 0.17893f
C24594 _0623_/a_109_297# acc0.A\[8\] 0
C24595 net167 _1072_/a_466_413# 0.00225f
C24596 _0170_ _1072_/a_27_47# 0.14208f
C24597 _0086_ clkbuf_1_1__f__0458_/a_110_47# 0.00213f
C24598 _1010_/a_1059_315# clknet_1_1__leaf__0462_ 0.02408f
C24599 acc0.A\[10\] _0345_ 0
C24600 control0.state\[1\] _0488_ 0.04299f
C24601 control0.state\[0\] _0466_ 0.12644f
C24602 _0738_/a_68_297# _0345_ 0.04112f
C24603 _0783_/a_297_297# clknet_1_1__leaf__0461_ 0
C24604 _0241_ clknet_0__0461_ 0
C24605 _0730_/a_297_297# net57 0
C24606 net123 comp0.B\[5\] 0
C24607 _0730_/a_79_21# _0195_ 0
C24608 clknet_1_0__leaf__0462_ _1025_/a_27_47# 0.05151f
C24609 clknet_1_1__leaf__0460_ _0462_ 0.11585f
C24610 _1056_/a_634_159# VPWR 0.18848f
C24611 _0993_/a_381_47# _0091_ 0.11658f
C24612 _0993_/a_1017_47# _0417_ 0
C24613 clknet_1_1__leaf__0459_ _0655_/a_109_93# 0
C24614 _0770_/a_382_297# _0770_/a_297_47# 0
C24615 _0512_/a_27_297# _0512_/a_373_47# 0.01338f
C24616 hold87/a_285_47# _0446_ 0
C24617 _0435_ _0436_ 0.07397f
C24618 hold86/a_285_47# _0350_ 0.00926f
C24619 VPWR comp0.B\[2\] 1.87454f
C24620 _0244_ _0294_ 0.00528f
C24621 net18 net129 0
C24622 _0179_ net189 0.0671f
C24623 net198 net196 0
C24624 _0695_/a_217_297# _0368_ 0
C24625 clknet_1_0__leaf__0465_ _1046_/a_1017_47# 0
C24626 clknet_1_1__leaf__0465_ hold81/a_49_47# 0
C24627 _0446_ _0529_/a_27_297# 0.00202f
C24628 _0343_ net69 0
C24629 _0322_ _0689_/a_68_297# 0
C24630 hold85/a_285_47# _0468_ 0
C24631 net175 net9 0
C24632 _0170_ _1071_/a_592_47# 0
C24633 _1028_/a_27_47# _0365_ 0
C24634 _0616_/a_78_199# _0460_ 0
C24635 _0996_/a_891_413# net5 0.02805f
C24636 _0996_/a_466_413# _0185_ 0
C24637 hold57/a_49_47# _1039_/a_466_413# 0
C24638 _0680_/a_300_47# _0219_ 0
C24639 clknet_0_clk _1068_/a_466_413# 0.00863f
C24640 _0227_ _0381_ 0
C24641 acc0.A\[21\] _0237_ 0.69892f
C24642 _0327_ _0689_/a_68_297# 0
C24643 control0.sh _0171_ 1.00042f
C24644 pp[6] output58/a_27_47# 0.01226f
C24645 VPWR _0433_ 0.51967f
C24646 _0259_ acc0.A\[9\] 0.09226f
C24647 output46/a_27_47# VPWR 0.31039f
C24648 _0100_ acc0.A\[20\] 0
C24649 _0340_ _0220_ 0.17729f
C24650 _0998_/a_891_413# net84 0.00162f
C24651 _1020_/a_1059_315# control0.add 0
C24652 net178 _1055_/a_634_159# 0
C24653 clknet_1_1__leaf__0459_ _0418_ 0.01396f
C24654 _0374_ _0754_/a_51_297# 0.02195f
C24655 net247 _0465_ 0.24799f
C24656 _0097_ _0306_ 0
C24657 _0101_ _0369_ 0.26145f
C24658 _0159_ _1061_/a_634_159# 0
C24659 net247 _1061_/a_381_47# 0
C24660 _1024_/a_592_47# acc0.A\[23\] 0
C24661 net203 _1033_/a_381_47# 0.00341f
C24662 hold56/a_49_47# net119 0.00524f
C24663 VPWR _0806_/a_113_297# 0.18964f
C24664 _0984_/a_381_47# net47 0.01405f
C24665 _0799_/a_209_297# _0409_ 0
C24666 control0.state\[0\] net236 0.02528f
C24667 net231 _1065_/a_193_47# 0
C24668 _1019_/a_466_413# net105 0.00222f
C24669 _1019_/a_634_159# net207 0.00325f
C24670 acc0.A\[2\] net247 0.00205f
C24671 _0267_ _0986_/a_27_47# 0
C24672 net51 _1005_/a_634_159# 0
C24673 _0271_ _0268_ 0
C24674 _0172_ _0544_/a_240_47# 0.02787f
C24675 _0725_/a_209_297# _0333_ 0.0396f
C24676 _1051_/a_891_413# acc0.A\[4\] 0
C24677 _0381_ _0759_/a_113_47# 0.0095f
C24678 hold52/a_391_47# _0122_ 0
C24679 _0949_/a_145_75# _0161_ 0
C24680 _0548_/a_149_47# net174 0
C24681 _0726_/a_245_297# _0354_ 0
C24682 _0726_/a_51_297# _0355_ 0.09161f
C24683 acc0.A\[12\] _0992_/a_27_47# 0
C24684 _0961_/a_113_297# clkbuf_1_0__f_clk/a_110_47# 0
C24685 _1058_/a_592_47# net67 0
C24686 comp0.B\[7\] net171 0.00965f
C24687 _0535_/a_68_297# _0139_ 0.00667f
C24688 net119 _1032_/a_27_47# 0
C24689 net36 clknet_1_1__leaf__0457_ 0.08542f
C24690 _0533_/a_109_47# _0178_ 0
C24691 net8 _0499_/a_59_75# 0
C24692 net242 _1010_/a_1059_315# 0.00572f
C24693 _0117_ _0345_ 0.0168f
C24694 _0465_ _0844_/a_382_297# 0
C24695 control0.state\[0\] _1064_/a_193_47# 0
C24696 control0.state\[1\] _1064_/a_27_47# 0
C24697 _0178_ hold71/a_285_47# 0
C24698 _0402_ hold70/a_49_47# 0.00105f
C24699 _0996_/a_27_47# clkbuf_1_1__f__0459_/a_110_47# 0
C24700 _0130_ _1032_/a_193_47# 0.00145f
C24701 hold64/a_285_47# _0461_ 0
C24702 _1015_/a_193_47# _0584_/a_109_297# 0
C24703 _1015_/a_634_159# _0584_/a_27_297# 0
C24704 _1050_/a_27_47# net170 0
C24705 _1050_/a_193_47# _0196_ 0
C24706 _1050_/a_381_47# _0528_/a_81_21# 0
C24707 _1001_/a_27_47# _0247_ 0
C24708 hold38/a_391_47# _1065_/a_27_47# 0
C24709 hold13/a_391_47# net8 0
C24710 net43 _0345_ 0.02661f
C24711 _0536_/a_240_47# _0176_ 0
C24712 _0180_ net149 0
C24713 net58 _0844_/a_79_21# 0.03658f
C24714 acc0.A\[2\] _0844_/a_382_297# 0
C24715 _0739_/a_79_21# _0739_/a_510_47# 0.00844f
C24716 _0739_/a_297_297# _0739_/a_215_47# 0
C24717 VPWR _0998_/a_975_413# 0.00418f
C24718 net149 net218 0.00307f
C24719 clkbuf_1_0__f__0457_/a_110_47# _1001_/a_27_47# 0
C24720 _1020_/a_27_47# hold40/a_391_47# 0
C24721 _1020_/a_193_47# hold40/a_285_47# 0
C24722 _0127_ hold50/a_285_47# 0
C24723 clknet_1_0__leaf__0465_ _0987_/a_592_47# 0
C24724 _0352_ _0739_/a_297_297# 0
C24725 _0990_/a_891_413# clknet_1_1__leaf__0465_ 0
C24726 _0731_/a_299_297# _0294_ 0
C24727 _0465_ _1048_/a_466_413# 0.00133f
C24728 _0999_/a_193_47# _0395_ 0
C24729 _0965_/a_129_47# VPWR 0
C24730 _1006_/a_27_47# net51 0
C24731 net33 net231 0.0013f
C24732 net157 _0171_ 0.1779f
C24733 _0751_/a_29_53# net51 0
C24734 _0990_/a_466_413# _0088_ 0.02982f
C24735 _0216_ _1007_/a_27_47# 0
C24736 _0108_ _0334_ 0
C24737 net125 _0498_/a_512_297# 0
C24738 input13/a_75_212# net13 0.10988f
C24739 _1002_/a_592_47# _0460_ 0
C24740 _0152_ _0186_ 0
C24741 _0999_/a_27_47# _0345_ 0
C24742 _1032_/a_891_413# _0165_ 0
C24743 acc0.A\[2\] _1048_/a_466_413# 0
C24744 _0793_/a_245_297# _0793_/a_240_47# 0
C24745 net67 _0186_ 0
C24746 _0205_ _0543_/a_68_297# 0
C24747 acc0.A\[27\] hold8/a_391_47# 0.00236f
C24748 _0273_ _0621_/a_285_297# 0
C24749 clknet_1_1__leaf__0459_ _0996_/a_1059_315# 0
C24750 net45 _0567_/a_109_297# 0
C24751 input31/a_75_212# comp0.B\[10\] 0
C24752 net59 net239 0.10781f
C24753 net46 hold29/a_285_47# 0.0329f
C24754 _0598_/a_79_21# _0382_ 0
C24755 _0598_/a_297_47# _0237_ 0.00594f
C24756 hold65/a_285_47# _0399_ 0.05077f
C24757 _0107_ _0691_/a_68_297# 0
C24758 _0228_ _0755_/a_109_297# 0
C24759 _0174_ _0139_ 0.02375f
C24760 _0564_/a_68_297# _0215_ 0.10647f
C24761 _1050_/a_1059_315# _0180_ 0.01627f
C24762 _0743_/a_149_47# _0368_ 0.00797f
C24763 clknet_1_0__leaf__0458_ _0267_ 0.05329f
C24764 _0958_/a_27_47# _0468_ 0.14405f
C24765 _0130_ _0721_/a_27_47# 0
C24766 _0465_ _0841_/a_79_21# 0
C24767 comp0.B\[7\] _1039_/a_466_413# 0
C24768 _0327_ acc0.A\[24\] 0
C24769 clknet_1_1__leaf__0463_ _0160_ 0
C24770 _0123_ _1025_/a_975_413# 0
C24771 net213 clknet_1_0__leaf__0460_ 0.00318f
C24772 net200 _1025_/a_381_47# 0.13012f
C24773 _0995_/a_27_47# acc0.A\[13\] 0.00107f
C24774 _1034_/a_193_47# _0474_ 0
C24775 _1034_/a_466_413# comp0.B\[6\] 0.00587f
C24776 _1034_/a_1059_315# comp0.B\[5\] 0
C24777 hold21/a_391_47# net63 0
C24778 net57 hold80/a_49_47# 0.35228f
C24779 _0777_/a_47_47# clknet_1_1__leaf__0461_ 0.01032f
C24780 _0699_/a_68_297# clkbuf_1_1__f__0462_/a_110_47# 0.00521f
C24781 _1051_/a_634_159# _1051_/a_381_47# 0
C24782 pp[17] VPWR 0.46335f
C24783 _1045_/a_27_47# _1044_/a_27_47# 0
C24784 comp0.B\[14\] _1042_/a_193_47# 0.00161f
C24785 clknet_1_1__leaf_clk _0215_ 0.02223f
C24786 _1056_/a_891_413# clknet_1_1__leaf__0465_ 0
C24787 _0347_ _0774_/a_150_297# 0
C24788 acc0.A\[21\] _1005_/a_27_47# 0
C24789 hold15/a_285_47# hold61/a_49_47# 0
C24790 _0368_ _0345_ 0
C24791 _0992_/a_27_47# _0650_/a_68_297# 0
C24792 pp[27] _0705_/a_145_75# 0
C24793 _1070_/a_891_413# control0.count\[1\] 0.01092f
C24794 _1070_/a_1017_47# VPWR 0
C24795 _1045_/a_466_413# _1045_/a_592_47# 0.00553f
C24796 _1045_/a_634_159# _1045_/a_1017_47# 0
C24797 _0195_ _0509_/a_27_47# 0.02621f
C24798 _0343_ net102 0
C24799 hold55/a_285_47# net106 0.06356f
C24800 acc0.A\[22\] acc0.A\[23\] 0.00313f
C24801 _0120_ net177 0.0145f
C24802 VPWR _1043_/a_891_413# 0.18631f
C24803 _0309_ _0308_ 0.33159f
C24804 _0852_/a_35_297# _0261_ 0
C24805 net44 _0568_/a_27_297# 0
C24806 clkbuf_0__0460_/a_110_47# hold90/a_391_47# 0
C24807 net100 _0465_ 0
C24808 _0209_ B[6] 0
C24809 clknet_0__0457_ net23 0
C24810 _0218_ _0986_/a_193_47# 0
C24811 _0356_ _0347_ 0
C24812 _1018_/a_466_413# _0399_ 0
C24813 _1038_/a_193_47# _0175_ 0
C24814 _0733_/a_448_47# _0697_/a_300_47# 0
C24815 _1043_/a_466_413# _1043_/a_592_47# 0.00553f
C24816 _1043_/a_634_159# _1043_/a_1017_47# 0
C24817 hold18/a_49_47# _0265_ 0
C24818 hold18/a_391_47# net47 0.00165f
C24819 VPWR _1015_/a_193_47# 0.30764f
C24820 clknet_0__0459_ _0655_/a_215_53# 0
C24821 hold58/a_49_47# _1037_/a_1059_315# 0
C24822 _0574_/a_27_297# _0352_ 0
C24823 hold88/a_391_47# acc0.A\[8\] 0.06578f
C24824 clkbuf_0__0464_/a_110_47# _0540_/a_51_297# 0.01224f
C24825 _0459_ _0247_ 0.0301f
C24826 input11/a_75_212# A[4] 0.19676f
C24827 _0554_/a_68_297# net24 0.04039f
C24828 _0734_/a_47_47# acc0.A\[27\] 0.01375f
C24829 _0176_ _1046_/a_27_47# 0
C24830 _1042_/a_27_47# net127 0
C24831 _0961_/a_113_297# control0.count\[2\] 0.00758f
C24832 _1030_/a_27_47# _0128_ 0
C24833 net216 _0370_ 0.0535f
C24834 _0384_ _0460_ 0.00366f
C24835 clknet_0__0464_ clknet_1_1__leaf__0464_ 0.19376f
C24836 _1004_/a_1017_47# VPWR 0
C24837 VPWR A[2] 0.20481f
C24838 _1054_/a_193_47# _1054_/a_381_47# 0.09503f
C24839 _1054_/a_634_159# _1054_/a_891_413# 0.03684f
C24840 _1054_/a_27_47# _1054_/a_561_413# 0.0027f
C24841 _0786_/a_217_297# _0369_ 0.00179f
C24842 hold11/a_285_47# clkbuf_0__0464_/a_110_47# 0
C24843 net187 _0218_ 0.00253f
C24844 _1071_/a_634_159# control0.count\[0\] 0
C24845 _1071_/a_381_47# clknet_1_0__leaf_clk 0
C24846 _1015_/a_27_47# _1015_/a_1059_315# 0.04875f
C24847 _1015_/a_193_47# _1015_/a_466_413# 0.07402f
C24848 _0983_/a_1059_315# VPWR 0.40484f
C24849 _0375_ net50 0
C24850 _0814_/a_109_47# _0181_ 0
C24851 _0982_/a_891_413# acc0.A\[1\] 0
C24852 input8/a_75_212# A[1] 0.19873f
C24853 _0347_ _0773_/a_35_297# 0
C24854 clknet_1_1__leaf__0462_ _1027_/a_634_159# 0.00543f
C24855 net113 _1027_/a_27_47# 0.23641f
C24856 net35 _0369_ 0
C24857 _0792_/a_209_297# _0405_ 0.09039f
C24858 _0792_/a_80_21# _0400_ 0.04345f
C24859 acc0.A\[30\] hold92/a_391_47# 0
C24860 _0195_ net47 0.00507f
C24861 _1020_/a_27_47# comp0.B\[0\] 0
C24862 _1038_/a_634_159# _1038_/a_466_413# 0.23992f
C24863 _1038_/a_193_47# _1038_/a_1059_315# 0.03405f
C24864 _1038_/a_27_47# _1038_/a_891_413# 0.03224f
C24865 _0556_/a_68_297# _1037_/a_466_413# 0
C24866 _0245_ _0392_ 0.03908f
C24867 _0472_ _0498_/a_51_297# 0.0025f
C24868 _0082_ _0450_ 0
C24869 net222 _0451_ 0.1352f
C24870 _0411_ _0797_/a_297_47# 0
C24871 _0199_ _0145_ 0.04021f
C24872 _0319_ _1008_/a_193_47# 0
C24873 _0655_/a_215_53# _0655_/a_109_93# 0.13675f
C24874 _0469_ net17 0
C24875 _0442_ _0830_/a_79_21# 0
C24876 _0343_ _0300_ 0
C24877 control0.state\[1\] _1065_/a_193_47# 0.00147f
C24878 clknet_0__0465_ _0347_ 0.00183f
C24879 hold2/a_285_47# _0181_ 0
C24880 net194 _0196_ 0
C24881 net61 _0529_/a_27_297# 0.00526f
C24882 _0157_ _1060_/a_975_413# 0
C24883 _1059_/a_975_413# _0158_ 0
C24884 _0983_/a_634_159# _0983_/a_975_413# 0
C24885 _0983_/a_466_413# _0983_/a_561_413# 0.00772f
C24886 _0983_/a_193_47# _0983_/a_592_47# 0
C24887 _0990_/a_27_47# acc0.A\[6\] 0
C24888 clknet_1_0__leaf__0465_ _1051_/a_381_47# 0.00265f
C24889 net41 pp[14] 0.01789f
C24890 _0217_ hold60/a_285_47# 0.01979f
C24891 _0700_/a_113_47# clknet_1_1__leaf__0462_ 0
C24892 clknet_1_0__leaf__0465_ _1045_/a_975_413# 0
C24893 _0352_ _0757_/a_150_297# 0
C24894 _0758_/a_510_47# _0380_ 0.00225f
C24895 _0262_ _0844_/a_79_21# 0.00173f
C24896 net40 _0995_/a_634_159# 0.00395f
C24897 net245 _0995_/a_27_47# 0.0337f
C24898 net234 _0452_ 0.01712f
C24899 hold29/a_391_47# VPWR 0.18948f
C24900 _0574_/a_27_297# _0574_/a_109_297# 0.17136f
C24901 net105 _0352_ 0
C24902 _0985_/a_466_413# net71 0
C24903 _0659_/a_68_297# _0659_/a_150_297# 0.00477f
C24904 _0143_ _0954_/a_32_297# 0
C24905 _0201_ comp0.B\[11\] 0
C24906 _0399_ acc0.A\[13\] 0.02044f
C24907 _0326_ _0352_ 0.01458f
C24908 pp[28] _0705_/a_59_75# 0
C24909 output56/a_27_47# _0220_ 0
C24910 _0389_ VPWR 0.46813f
C24911 _0386_ _0391_ 0
C24912 _1026_/a_1059_315# _0320_ 0
C24913 net8 _0206_ 0
C24914 net71 _1049_/a_27_47# 0
C24915 net219 hold72/a_49_47# 0.00105f
C24916 _0371_ _0350_ 0.02022f
C24917 _0206_ net32 0
C24918 _0742_/a_384_47# acc0.A\[23\] 0
C24919 _0466_ _1068_/a_193_47# 0.03679f
C24920 _1056_/a_466_413# hold35/a_285_47# 0.00145f
C24921 net90 _1007_/a_634_159# 0
C24922 net45 _0612_/a_59_75# 0.18325f
C24923 _0113_ net201 0
C24924 _0118_ _0217_ 0
C24925 _1048_/a_27_47# _1047_/a_27_47# 0
C24926 _0637_/a_56_297# _0269_ 0.00416f
C24927 _0831_/a_285_297# _0369_ 0.00413f
C24928 _1003_/a_1059_315# _0183_ 0.01266f
C24929 net64 hold88/a_391_47# 0
C24930 _1004_/a_193_47# net50 0
C24931 _0343_ _0827_/a_27_47# 0
C24932 _0852_/a_35_297# net47 0.10111f
C24933 _0698_/a_113_297# _0322_ 0.06797f
C24934 _0785_/a_299_297# _0785_/a_384_47# 0
C24935 _1016_/a_891_413# _1016_/a_1017_47# 0.00617f
C24936 _1016_/a_193_47# net166 0.19755f
C24937 hold10/a_49_47# acc0.A\[15\] 0.01203f
C24938 clkload2/Y _1050_/a_466_413# 0
C24939 _0331_ _0330_ 0.0495f
C24940 VPWR _0355_ 0.50476f
C24941 clknet_0__0459_ _0996_/a_466_413# 0.00151f
C24942 net158 _1061_/a_381_47# 0
C24943 control0.state\[1\] net33 0
C24944 _0379_ acc0.A\[23\] 0.03807f
C24945 comp0.B\[1\] comp0.B\[15\] 0.45992f
C24946 net113 _1026_/a_466_413# 0
C24947 clknet_1_1__leaf__0462_ _1026_/a_891_413# 0.00775f
C24948 clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0462_ 0.0073f
C24949 _0478_ _0466_ 0.16528f
C24950 _0998_/a_27_47# _0398_ 0.02102f
C24951 _0329_ _0701_/a_303_47# 0
C24952 clkbuf_1_1__f__0465_/a_110_47# _0426_ 0
C24953 _0458_ _0350_ 0.02817f
C24954 _0555_/a_51_297# _0176_ 0.01689f
C24955 _1057_/a_1017_47# _0187_ 0.00172f
C24956 _0107_ _0361_ 0
C24957 _0313_ _0687_/a_145_75# 0
C24958 net19 hold51/a_49_47# 0
C24959 net195 hold51/a_285_47# 0
C24960 net85 _0399_ 0
C24961 control0.state\[1\] hold12/a_391_47# 0
C24962 _0471_ _0951_/a_109_93# 0
C24963 _0227_ _0468_ 0
C24964 _0455_ _0265_ 0
C24965 _0081_ net47 0.00303f
C24966 _0514_/a_109_297# _0189_ 0.00169f
C24967 _0514_/a_373_47# net2 0
C24968 _0179_ _0511_/a_384_47# 0
C24969 _0849_/a_215_47# _0347_ 0.00683f
C24970 _0134_ _1037_/a_466_413# 0
C24971 _0984_/a_193_47# _0450_ 0
C24972 _1059_/a_975_413# acc0.A\[14\] 0
C24973 hold54/a_49_47# _0131_ 0
C24974 _0201_ _0202_ 0.00514f
C24975 _0538_/a_240_47# net20 0.00374f
C24976 _0538_/a_245_297# _0142_ 0
C24977 hold42/a_285_47# acc0.A\[11\] 0.03342f
C24978 _1041_/a_975_413# net7 0.00201f
C24979 net160 _1035_/a_27_47# 0
C24980 clknet_1_1__leaf__0459_ _1057_/a_466_413# 0
C24981 _1057_/a_1059_315# acc0.A\[11\] 0.08745f
C24982 _0403_ _0091_ 0.01183f
C24983 net82 _0781_/a_68_297# 0
C24984 _0978_/a_27_297# control0.count\[0\] 0
C24985 _0413_ net5 0.02158f
C24986 hold54/a_391_47# _0130_ 0.00114f
C24987 _0368_ net52 0.02731f
C24988 _1015_/a_1059_315# _0215_ 0
C24989 _0378_ hold94/a_49_47# 0
C24990 VPWR _0693_/a_150_297# 0.00224f
C24991 comp0.B\[4\] _1034_/a_27_47# 0
C24992 _1036_/a_27_47# comp0.B\[2\] 0
C24993 _1048_/a_193_47# _0509_/a_27_47# 0
C24994 _0322_ _0691_/a_68_297# 0.10235f
C24995 _1052_/a_27_47# _0252_ 0
C24996 comp0.B\[13\] _0139_ 0
C24997 _0343_ _0404_ 0.0022f
C24998 hold76/a_285_47# _0183_ 0
C24999 _0343_ _0754_/a_149_47# 0
C25000 _0233_ _0754_/a_245_297# 0
C25001 _0663_/a_27_413# _0812_/a_215_47# 0
C25002 _0356_ hold95/a_49_47# 0
C25003 _1056_/a_634_159# net182 0.00212f
C25004 _0327_ _0691_/a_68_297# 0
C25005 hold18/a_49_47# _0267_ 0
C25006 _1004_/a_27_47# net215 0
C25007 _1004_/a_891_413# hold68/a_391_47# 0
C25008 _0734_/a_47_47# _1009_/a_634_159# 0
C25009 _1054_/a_975_413# VPWR 0.00488f
C25010 _0272_ _0626_/a_68_297# 0
C25011 _0643_/a_253_297# _0258_ 0
C25012 clknet_0_clk _0564_/a_150_297# 0
C25013 _0517_/a_299_297# _0190_ 0.00863f
C25014 net236 _0478_ 0
C25015 _0618_/a_215_47# net52 0
C25016 VPWR _0569_/a_27_297# 0.30306f
C25017 acc0.A\[5\] _0987_/a_891_413# 0.01743f
C25018 net137 _0987_/a_592_47# 0
C25019 hold39/a_49_47# _0473_ 0
C25020 net63 _0519_/a_81_21# 0.00407f
C25021 hold34/a_49_47# net181 0
C25022 clknet_1_0__leaf__0459_ _1015_/a_193_47# 0
C25023 _0163_ _1065_/a_466_413# 0.03747f
C25024 _0389_ _0390_ 0.02519f
C25025 clkbuf_1_1__f__0459_/a_110_47# _0794_/a_27_47# 0
C25026 _1038_/a_561_413# VPWR 0.00318f
C25027 _0697_/a_80_21# clknet_0__0460_ 0
C25028 clkbuf_0__0465_/a_110_47# clknet_0__0465_ 1.70156f
C25029 clkbuf_1_0__f__0458_/a_110_47# _0261_ 0
C25030 net154 net148 0.02346f
C25031 _1041_/a_561_413# A[15] 0
C25032 _0222_ pp[23] 0
C25033 hold39/a_391_47# _0133_ 0.00771f
C25034 comp0.B\[10\] _0548_/a_51_297# 0.00275f
C25035 _0387_ _0347_ 0.01033f
C25036 _1018_/a_592_47# acc0.A\[18\] 0.00287f
C25037 _0731_/a_81_21# _0359_ 0.12585f
C25038 net35 _1072_/a_27_47# 0.0034f
C25039 _1067_/a_466_413# clknet_1_0__leaf__0457_ 0.0107f
C25040 _0206_ net10 0
C25041 clkload3/Y _0096_ 0
C25042 _1067_/a_193_47# _0460_ 0
C25043 hold36/a_285_47# VPWR 0.28434f
C25044 _0487_ _0969_/a_109_297# 0.01446f
C25045 hold21/a_285_47# input11/a_75_212# 0
C25046 _0196_ _0987_/a_193_47# 0
C25047 net62 clkbuf_0__0458_/a_110_47# 0.00124f
C25048 clknet_0_clk _0166_ 0.01784f
C25049 _0383_ _0460_ 0.0025f
C25050 net188 _0515_/a_81_21# 0
C25051 _0983_/a_1059_315# clknet_1_0__leaf__0459_ 0
C25052 net120 _1065_/a_561_413# 0
C25053 _0450_ clkbuf_0__0458_/a_110_47# 0.00171f
C25054 comp0.B\[2\] _0113_ 0
C25055 clknet_1_0__leaf__0460_ _0618_/a_510_47# 0
C25056 _0816_/a_68_297# _0345_ 0.00583f
C25057 _0816_/a_68_297# _0814_/a_27_47# 0
C25058 net178 net141 0
C25059 _0374_ _0219_ 0.30658f
C25060 _0241_ _0616_/a_215_47# 0.02988f
C25061 clknet_0__0463_ _0563_/a_512_297# 0
C25062 _0760_/a_47_47# _0760_/a_129_47# 0.00369f
C25063 _0557_/a_51_297# net27 0.10923f
C25064 _0159_ net147 0.04157f
C25065 clknet_1_0__leaf__0462_ _0314_ 0.16077f
C25066 hold31/a_285_47# _0988_/a_193_47# 0
C25067 hold31/a_391_47# _0988_/a_27_47# 0.00179f
C25068 _0819_/a_299_297# _0181_ 0.00245f
C25069 VPWR _0266_ 0.79454f
C25070 net203 comp0.B\[1\] 0
C25071 pp[17] _0567_/a_373_47# 0
C25072 hold101/a_49_47# _0218_ 0.01301f
C25073 clkbuf_0__0459_/a_110_47# net228 0
C25074 _0487_ _0950_/a_75_212# 0
C25075 clknet_1_1__leaf__0459_ _0297_ 0.10876f
C25076 net121 net28 0
C25077 _1031_/a_27_47# _1030_/a_1059_315# 0
C25078 _1031_/a_193_47# _1030_/a_466_413# 0
C25079 _1031_/a_466_413# _1030_/a_193_47# 0
C25080 _0408_ net41 0
C25081 net105 net207 0.5473f
C25082 _0714_/a_240_47# _0111_ 0.0017f
C25083 VPWR _0567_/a_109_297# 0.1775f
C25084 clknet_1_0__leaf__0458_ _0178_ 0
C25085 _0457_ _1067_/a_193_47# 0.00251f
C25086 net35 _1071_/a_592_47# 0
C25087 _0467_ hold84/a_391_47# 0
C25088 net248 _0186_ 0
C25089 net51 net91 0
C25090 _0299_ acc0.A\[13\] 0.29675f
C25091 _1032_/a_634_159# comp0.B\[15\] 0
C25092 _0507_/a_27_297# _0219_ 0.01756f
C25093 _1038_/a_381_47# _0550_/a_51_297# 0
C25094 _1038_/a_466_413# _0550_/a_149_47# 0
C25095 clknet_1_1__leaf__0460_ _0312_ 0.46352f
C25096 net43 _0394_ 0
C25097 _0382_ hold3/a_391_47# 0.00108f
C25098 _0627_/a_215_53# _0465_ 0
C25099 _0712_/a_297_297# _0708_/a_150_297# 0
C25100 _0343_ _0995_/a_592_47# 0
C25101 _1014_/a_1017_47# clknet_1_0__leaf__0461_ 0
C25102 _1025_/a_634_159# _1025_/a_466_413# 0.23992f
C25103 _1025_/a_193_47# _1025_/a_1059_315# 0.03405f
C25104 _1025_/a_27_47# _1025_/a_891_413# 0.03224f
C25105 net199 net50 0.01419f
C25106 net49 _1005_/a_193_47# 0.00225f
C25107 net122 B[2] 0
C25108 _0359_ _1006_/a_193_47# 0
C25109 _0324_ _1006_/a_27_47# 0
C25110 _0295_ acc0.A\[13\] 0
C25111 clknet_0__0461_ net219 0.01175f
C25112 _1012_/a_634_159# _0345_ 0
C25113 _0770_/a_382_297# _0462_ 0
C25114 hold35/a_49_47# VPWR 0.27913f
C25115 _0317_ _0219_ 0
C25116 _0343_ _0228_ 0
C25117 _0179_ _1055_/a_891_413# 0
C25118 _0412_ clknet_1_1__leaf__0459_ 0.23075f
C25119 net45 _0399_ 0.03866f
C25120 net34 _1064_/a_1017_47# 0
C25121 net165 _0219_ 0
C25122 _1015_/a_561_413# net157 0
C25123 _1055_/a_193_47# _0181_ 0
C25124 hold28/a_285_47# _0195_ 0.02576f
C25125 VPWR _0522_/a_109_47# 0
C25126 acc0.A\[4\] _0528_/a_81_21# 0
C25127 _1070_/a_193_47# _0466_ 0.00264f
C25128 _1070_/a_634_159# _0488_ 0
C25129 VPWR _0976_/a_505_21# 0.17529f
C25130 net187 _0099_ 0
C25131 _0359_ acc0.A\[25\] 0.06611f
C25132 _0800_/a_245_297# VPWR 0.00648f
C25133 comp0.B\[0\] hold84/a_391_47# 0
C25134 _0432_ _0256_ 0.13999f
C25135 _0443_ _0271_ 0.22445f
C25136 _1059_/a_381_47# net228 0
C25137 clkbuf_1_0__f__0457_/a_110_47# _0772_/a_79_21# 0.00968f
C25138 _1046_/a_1059_315# net10 0.07785f
C25139 clkbuf_1_1__f__0458_/a_110_47# _0350_ 0
C25140 _0467_ _1065_/a_975_413# 0.00261f
C25141 net115 acc0.A\[28\] 0.10337f
C25142 _1021_/a_27_47# _1067_/a_1059_315# 0.00185f
C25143 _0516_/a_27_297# _0990_/a_1059_315# 0
C25144 _0195_ _1047_/a_1017_47# 0
C25145 _0097_ _0778_/a_68_297# 0
C25146 hold18/a_285_47# _0848_/a_27_47# 0
C25147 _1003_/a_634_159# control0.state\[2\] 0
C25148 _1003_/a_193_47# _0486_ 0
C25149 control0.reset clkbuf_1_1__f__0457_/a_110_47# 0
C25150 _1021_/a_891_413# _0369_ 0
C25151 _0996_/a_193_47# _0996_/a_381_47# 0.09799f
C25152 _0996_/a_634_159# _0996_/a_891_413# 0.03684f
C25153 _0996_/a_27_47# _0996_/a_561_413# 0.0027f
C25154 clknet_0__0465_ _0824_/a_59_75# 0.00734f
C25155 net140 net9 0
C25156 _0427_ _0424_ 0
C25157 _0769_/a_81_21# _0352_ 0.05903f
C25158 net45 _1031_/a_27_47# 0
C25159 _0209_ comp0.B\[5\] 0
C25160 VPWR _0835_/a_78_199# 0.2728f
C25161 _0174_ _0498_/a_240_47# 0.05995f
C25162 _0156_ acc0.A\[10\] 0.00267f
C25163 net125 _0159_ 0.00291f
C25164 _0139_ comp0.B\[9\] 0
C25165 _0835_/a_215_47# _0636_/a_59_75# 0
C25166 clknet_1_0__leaf__0464_ _1048_/a_634_159# 0
C25167 net133 _1048_/a_27_47# 0
C25168 _0276_ acc0.A\[14\] 0
C25169 clknet_1_1__leaf__0457_ _1061_/a_27_47# 0
C25170 _0793_/a_149_47# _0095_ 0
C25171 output46/a_27_47# pp[22] 0.00337f
C25172 _0329_ hold50/a_49_47# 0
C25173 _0646_/a_129_47# net5 0
C25174 _0343_ net16 0
C25175 _0234_ _0345_ 0.05259f
C25176 _0376_ _0754_/a_149_47# 0.018f
C25177 _0430_ pp[2] 0
C25178 hold56/a_391_47# net203 0.14549f
C25179 hold57/a_285_47# _0473_ 0.00226f
C25180 _0559_/a_240_47# _0175_ 0
C25181 hold8/a_285_47# _1027_/a_27_47# 0.00319f
C25182 hold8/a_49_47# _1027_/a_193_47# 0
C25183 VPWR _0996_/a_975_413# 0.00487f
C25184 acc0.A\[7\] A[8] 0.19983f
C25185 clkbuf_1_0__f__0458_/a_110_47# net47 0.00223f
C25186 _0477_ _0468_ 0.25615f
C25187 _0344_ _0999_/a_193_47# 0.00131f
C25188 _0621_/a_35_297# clkbuf_1_1__f__0458_/a_110_47# 0
C25189 comp0.B\[7\] _0553_/a_51_297# 0
C25190 _0330_ _1008_/a_27_47# 0
C25191 _0317_ _1008_/a_634_159# 0
C25192 _1065_/a_975_413# comp0.B\[0\] 0.00102f
C25193 _0726_/a_149_47# acc0.A\[29\] 0
C25194 _0672_/a_79_21# clkbuf_1_1__f__0459_/a_110_47# 0.00734f
C25195 net200 acc0.A\[25\] 0.29558f
C25196 _0483_ clkbuf_1_0__f_clk/a_110_47# 0.00217f
C25197 VPWR A[9] 0.27853f
C25198 comp0.B\[2\] comp0.B\[3\] 0
C25199 _1037_/a_1017_47# net28 0
C25200 hold33/a_391_47# _1041_/a_1059_315# 0
C25201 _1051_/a_634_159# acc0.A\[5\] 0
C25202 _1051_/a_381_47# net137 0
C25203 _1051_/a_891_413# _0149_ 0
C25204 hold22/a_391_47# _1054_/a_634_159# 0
C25205 hold22/a_49_47# _1054_/a_1059_315# 0.0037f
C25206 _0336_ acc0.A\[30\] 0.24401f
C25207 _0195_ _0294_ 0.02686f
C25208 net58 _0084_ 0.08354f
C25209 _0349_ _0729_/a_68_297# 0
C25210 clknet_0__0458_ _0831_/a_35_297# 0.0013f
C25211 _0762_/a_510_47# net51 0.00201f
C25212 _0992_/a_891_413# acc0.A\[10\] 0.06954f
C25213 _1051_/a_975_413# net131 0
C25214 _0289_ clkbuf_1_1__f__0465_/a_110_47# 0.00112f
C25215 _0805_/a_27_47# _0285_ 0.00664f
C25216 _0670_/a_79_21# net238 0
C25217 net29 _0175_ 0
C25218 clknet_0__0460_ _0345_ 0
C25219 net62 _0986_/a_975_413# 0
C25220 net22 _1040_/a_1059_315# 0
C25221 net23 _1067_/a_1017_47# 0.00226f
C25222 _0101_ hold66/a_391_47# 0.06881f
C25223 _0399_ _0990_/a_1059_315# 0.0419f
C25224 _0404_ A[14] 0
C25225 net44 _0128_ 0
C25226 _0270_ net10 0
C25227 hold47/a_285_47# clknet_1_1__leaf__0464_ 0.00283f
C25228 _0249_ _0219_ 0.02467f
C25229 _0440_ hold1/a_49_47# 0.02253f
C25230 net114 _0350_ 0
C25231 net245 _0299_ 0.00428f
C25232 _1002_/a_891_413# net240 0
C25233 _0361_ _0322_ 0.0291f
C25234 net88 _0973_/a_27_297# 0
C25235 _0984_/a_561_413# _0158_ 0
C25236 _0324_ _0737_/a_35_297# 0
C25237 _0369_ _0796_/a_215_47# 0.07382f
C25238 _1060_/a_193_47# net229 0
C25239 _0714_/a_51_297# _1013_/a_193_47# 0
C25240 acc0.A\[21\] net220 0.06857f
C25241 _1003_/a_466_413# _0467_ 0
C25242 _0713_/a_27_47# VPWR 0.50939f
C25243 clkload3/a_268_47# _0219_ 0.00152f
C25244 _0361_ _0327_ 0.0249f
C25245 _0403_ _0346_ 0
C25246 acc0.A\[14\] _0854_/a_79_21# 0
C25247 acc0.A\[20\] net150 0
C25248 _1030_/a_634_159# _0345_ 0
C25249 hold96/a_49_47# net93 0
C25250 _0972_/a_93_21# _1062_/a_27_47# 0
C25251 hold76/a_49_47# _1000_/a_27_47# 0
C25252 _0662_/a_299_297# _0817_/a_81_21# 0
C25253 clknet_1_0__leaf__0463_ _1040_/a_1059_315# 0.00781f
C25254 hold3/a_49_47# _1005_/a_1059_315# 0
C25255 hold3/a_285_47# _1005_/a_466_413# 0
C25256 hold67/a_285_47# _0428_ 0.00308f
C25257 _0984_/a_27_47# net233 0
C25258 _1039_/a_27_47# clknet_1_1__leaf__0457_ 0
C25259 control0.count\[1\] clkbuf_1_0__f_clk/a_110_47# 0.02644f
C25260 _0119_ _1002_/a_592_47# 0
C25261 A[9] output62/a_27_47# 0
C25262 _1032_/a_1059_315# _1032_/a_891_413# 0.31086f
C25263 _1032_/a_193_47# _1032_/a_975_413# 0
C25264 _1032_/a_466_413# _1032_/a_381_47# 0.03733f
C25265 _1054_/a_891_413# net140 0
C25266 net158 clknet_0__0464_ 0.06153f
C25267 output42/a_27_47# hold98/a_391_47# 0.01549f
C25268 _1015_/a_891_413# _1015_/a_1017_47# 0.00617f
C25269 _1015_/a_193_47# _0113_ 0.19374f
C25270 _1038_/a_1059_315# net29 0.01682f
C25271 hold5/a_49_47# _0176_ 0
C25272 _0569_/a_27_297# _0569_/a_109_47# 0.00393f
C25273 _0357_ _1010_/a_592_47# 0
C25274 _0108_ _1010_/a_381_47# 0.14004f
C25275 _0598_/a_297_47# _0222_ 0
C25276 _0753_/a_561_47# clknet_1_0__leaf__0460_ 0.00104f
C25277 VPWR _0612_/a_59_75# 0.21009f
C25278 hold33/a_285_47# net147 0
C25279 _1051_/a_193_47# _0180_ 0.03734f
C25280 _0376_ _0228_ 0.00306f
C25281 _0343_ _1031_/a_592_47# 0
C25282 A[12] input16/a_75_212# 0
C25283 _1014_/a_1059_315# net149 0.03217f
C25284 _0319_ _0318_ 0.01324f
C25285 _0611_/a_68_297# _0242_ 0.10185f
C25286 _1038_/a_634_159# net172 0.00257f
C25287 _1038_/a_466_413# net124 0
C25288 _0600_/a_103_199# _0352_ 0.02045f
C25289 net33 _1066_/a_634_159# 0.03714f
C25290 _0473_ _0159_ 0.00925f
C25291 _0729_/a_68_297# _0701_/a_209_297# 0
C25292 _0731_/a_299_297# _0371_ 0.00245f
C25293 _0430_ clknet_1_0__leaf__0465_ 0
C25294 _1067_/a_975_413# clknet_1_0__leaf__0461_ 0.00107f
C25295 _0290_ net217 0
C25296 _0423_ _0422_ 0.00163f
C25297 B[12] comp0.B\[11\] 0.05776f
C25298 _0661_/a_205_297# _0345_ 0
C25299 _0637_/a_56_297# _0082_ 0
C25300 _0446_ _0449_ 0.06772f
C25301 clknet_1_0__leaf__0465_ _1044_/a_561_413# 0
C25302 pp[1] net179 0
C25303 pp[16] pp[31] 0.21852f
C25304 hold16/a_285_47# _1030_/a_193_47# 0.00171f
C25305 hold16/a_391_47# _1030_/a_27_47# 0
C25306 clknet_1_0__leaf__0465_ acc0.A\[5\] 0.11567f
C25307 _1020_/a_27_47# net1 0.02659f
C25308 _0289_ _0673_/a_253_47# 0.03049f
C25309 _0350_ _0365_ 0.09977f
C25310 _0287_ _0673_/a_337_297# 0.0015f
C25311 _0997_/a_193_47# net43 0.03632f
C25312 _0227_ _0762_/a_79_21# 0.01547f
C25313 clknet_0__0461_ _0352_ 0.31821f
C25314 VPWR net50 1.11451f
C25315 VPWR _0995_/a_27_47# 0.64682f
C25316 _0983_/a_193_47# acc0.A\[18\] 0
C25317 _0483_ control0.count\[2\] 0.06805f
C25318 clknet_1_1__leaf__0458_ _0445_ 0
C25319 net45 _0712_/a_79_21# 0.0012f
C25320 _0346_ _0610_/a_59_75# 0
C25321 _0083_ net71 0.00159f
C25322 _0225_ _0754_/a_51_297# 0.01407f
C25323 net66 _0291_ 0.05721f
C25324 _0081_ _0294_ 0
C25325 net88 net17 0
C25326 clknet_1_1__leaf__0460_ _1008_/a_466_413# 0
C25327 _0511_/a_81_21# net4 0.00138f
C25328 _0347_ _0986_/a_27_47# 0
C25329 control0.sh _0494_/a_27_47# 0.04313f
C25330 _0550_/a_149_47# _0550_/a_240_47# 0.06872f
C25331 _0240_ _0775_/a_79_21# 0.05501f
C25332 net197 _1008_/a_634_159# 0.00171f
C25333 net190 _1008_/a_27_47# 0
C25334 net216 _1006_/a_466_413# 0
C25335 _0104_ _1006_/a_27_47# 0.11697f
C25336 net106 _1032_/a_1059_315# 0
C25337 _0226_ _0765_/a_215_47# 0
C25338 acc0.A\[12\] _1058_/a_891_413# 0.0369f
C25339 _0369_ _0775_/a_79_21# 0
C25340 net90 net93 0.00193f
C25341 _0174_ _0954_/a_32_297# 0.00409f
C25342 hold32/a_49_47# _1055_/a_1059_315# 0.00791f
C25343 hold32/a_391_47# _1055_/a_634_159# 0
C25344 hold31/a_49_47# _0253_ 0.01287f
C25345 _0266_ _0453_ 0.31432f
C25346 _1054_/a_381_47# acc0.A\[6\] 0
C25347 _1000_/a_193_47# _0461_ 0.01424f
C25348 _0954_/a_220_297# comp0.B\[10\] 0
C25349 clknet_1_0__leaf__0462_ _1005_/a_975_413# 0
C25350 _0520_/a_109_47# net12 0
C25351 _0578_/a_109_47# _0352_ 0.00265f
C25352 acc0.A\[20\] control0.add 0.03226f
C25353 _0546_/a_51_297# _0546_/a_245_297# 0.01218f
C25354 _0616_/a_493_297# _0246_ 0.01124f
C25355 _0240_ _0614_/a_183_297# 0.00163f
C25356 _1036_/a_466_413# _0175_ 0.00224f
C25357 _0181_ hold93/a_285_47# 0.06085f
C25358 _0534_/a_81_21# _0182_ 0.02199f
C25359 _0534_/a_299_297# acc0.A\[1\] 0.00119f
C25360 net132 _0196_ 0.00157f
C25361 _0991_/a_27_47# _0991_/a_634_159# 0.14145f
C25362 VPWR _0516_/a_27_297# 0.28806f
C25363 _0998_/a_592_47# _0096_ 0.00164f
C25364 clknet_1_0__leaf__0464_ _0138_ 0
C25365 _0263_ _0445_ 0
C25366 control0.count\[2\] control0.count\[1\] 0.07021f
C25367 input20/a_75_212# net20 0.10861f
C25368 clknet_0__0464_ net148 0
C25369 _0580_/a_27_297# clknet_1_0__leaf__0457_ 0
C25370 _0356_ _1011_/a_27_47# 0
C25371 comp0.B\[14\] clknet_1_1__leaf__0464_ 0.02207f
C25372 comp0.B\[14\] _0548_/a_149_47# 0
C25373 _0535_/a_68_297# net173 0
C25374 _0241_ _0771_/a_215_297# 0.01679f
C25375 hold23/a_285_47# _0180_ 0.04922f
C25376 hold23/a_391_47# _0182_ 0
C25377 _0243_ _0612_/a_145_75# 0
C25378 net48 net50 0
C25379 comp0.B\[1\] _0176_ 0
C25380 _0447_ _0186_ 0
C25381 _0502_/a_27_47# _0147_ 0.00111f
C25382 hold67/a_391_47# net142 0.00109f
C25383 _0210_ _0957_/a_32_297# 0.01565f
C25384 net160 _0957_/a_114_297# 0
C25385 _0183_ hold4/a_391_47# 0.0528f
C25386 _0120_ hold4/a_49_47# 0.31828f
C25387 hold86/a_285_47# hold18/a_391_47# 0
C25388 A[3] B[11] 0
C25389 _0479_ _0488_ 0.25902f
C25390 _0291_ _0350_ 0
C25391 _0982_/a_466_413# _1014_/a_1059_315# 0.00255f
C25392 _0982_/a_634_159# _1014_/a_891_413# 0.00811f
C25393 _0833_/a_79_21# _0369_ 0.10469f
C25394 _0316_ _0737_/a_35_297# 0
C25395 _0684_/a_59_75# _0321_ 0
C25396 _0195_ _1017_/a_561_413# 0.00119f
C25397 clknet_1_1__leaf__0459_ net189 0
C25398 _1001_/a_27_47# _0217_ 0.04881f
C25399 _1054_/a_27_47# _0150_ 0.00146f
C25400 net88 acc0.A\[21\] 0
C25401 clknet_1_0__leaf__0462_ _0572_/a_27_297# 0
C25402 hold6/a_49_47# _1040_/a_27_47# 0
C25403 hold39/a_49_47# _0132_ 0.30104f
C25404 _0853_/a_68_297# _0181_ 0
C25405 clknet_1_0__leaf__0458_ _0347_ 1.35731f
C25406 _1057_/a_561_413# VPWR 0.00292f
C25407 clknet_1_0__leaf__0465_ _0443_ 0
C25408 _1048_/a_561_413# _0186_ 0
C25409 clknet_0__0460_ net52 0.02722f
C25410 net176 output50/a_27_47# 0
C25411 clkbuf_1_1__f__0462_/a_110_47# _1008_/a_1059_315# 0
C25412 _0231_ _0219_ 0.05584f
C25413 _0579_/a_109_297# VPWR 0.17779f
C25414 hold35/a_49_47# hold35/a_391_47# 0.00188f
C25415 hold13/a_391_47# hold57/a_49_47# 0
C25416 _0476_ clknet_1_1__leaf__0463_ 0.04156f
C25417 _0625_/a_59_75# _0825_/a_68_297# 0.00662f
C25418 _0347_ _0737_/a_35_297# 0
C25419 _0174_ _0540_/a_245_297# 0.00318f
C25420 acc0.A\[27\] hold9/a_285_47# 0
C25421 _0784_/a_113_47# _0400_ 0.00951f
C25422 net43 _0411_ 0
C25423 _0399_ _0439_ 0.30336f
C25424 VPWR _0127_ 0.24165f
C25425 _0251_ net75 0
C25426 clkbuf_0__0461_/a_110_47# net102 0.00105f
C25427 net1 _0219_ 0.00514f
C25428 _0343_ hold78/a_391_47# 0.04336f
C25429 net64 acc0.A\[8\] 0.36024f
C25430 _0315_ _1007_/a_891_413# 0
C25431 _0366_ _1007_/a_381_47# 0.01801f
C25432 _0174_ net173 0.13616f
C25433 _0713_/a_27_47# clknet_1_0__leaf__0459_ 0.03802f
C25434 _0188_ _0156_ 0
C25435 _0369_ _0161_ 0
C25436 VPWR _0399_ 6.46201f
C25437 _0522_/a_27_297# acc0.A\[6\] 0.10918f
C25438 hold65/a_49_47# _0434_ 0.00127f
C25439 _0257_ _0440_ 0.00215f
C25440 _0722_/a_297_297# _0347_ 0.00573f
C25441 _0976_/a_76_199# _0976_/a_218_47# 0.00783f
C25442 _0800_/a_51_297# _0800_/a_240_47# 0.03076f
C25443 clkbuf_1_1__f__0461_/a_110_47# _0219_ 0.01791f
C25444 acc0.A\[29\] _0568_/a_109_297# 0.0015f
C25445 hold87/a_285_47# _0269_ 0
C25446 _0290_ net66 0.08313f
C25447 _0855_/a_384_47# _0345_ 0
C25448 _1017_/a_381_47# _0369_ 0.00168f
C25449 _1002_/a_193_47# _0352_ 0
C25450 net44 _1031_/a_1059_315# 0
C25451 _0981_/a_27_297# _1068_/a_381_47# 0
C25452 clknet_1_1__leaf__0462_ net244 0
C25453 _0183_ _0261_ 0
C25454 _0996_/a_27_47# _0277_ 0
C25455 net248 net62 0
C25456 VPWR _0545_/a_68_297# 0.16982f
C25457 net185 net186 0
C25458 acc0.A\[16\] _0347_ 0.00662f
C25459 hold97/a_49_47# clknet_0__0462_ 0
C25460 _0369_ _0158_ 0
C25461 _0179_ hold7/a_285_47# 0.03213f
C25462 _0627_/a_215_53# _0254_ 0.28737f
C25463 clknet_1_0__leaf__0459_ _0612_/a_59_75# 0
C25464 VPWR _1031_/a_27_47# 0.68479f
C25465 _0381_ _0237_ 0.34877f
C25466 clkbuf_0__0465_/a_110_47# _0986_/a_27_47# 0.01708f
C25467 net178 _0988_/a_381_47# 0.02055f
C25468 hold31/a_49_47# net74 0
C25469 _0399_ _0654_/a_27_413# 0
C25470 _0216_ net223 0
C25471 net203 _0496_/a_27_47# 0
C25472 _0290_ _0991_/a_27_47# 0
C25473 _0423_ _0991_/a_193_47# 0
C25474 _0430_ net76 0
C25475 _0343_ net163 0
C25476 _0983_/a_381_47# _0399_ 0.01691f
C25477 _0749_/a_81_21# _0460_ 0.01203f
C25478 net51 _1022_/a_891_413# 0.02079f
C25479 net205 _0173_ 0.17133f
C25480 _0345_ _0806_/a_113_297# 0.00476f
C25481 net204 clkbuf_1_0__f__0463_/a_110_47# 0
C25482 hold26/a_49_47# VPWR 0.27717f
C25483 hold42/a_285_47# A[12] 0
C25484 hold35/a_391_47# A[9] 0.00556f
C25485 _0835_/a_78_199# _0835_/a_493_297# 0
C25486 _0185_ _0219_ 0.02741f
C25487 _0399_ output62/a_27_47# 0
C25488 net8 A[1] 0.00671f
C25489 hold35/a_49_47# net182 0.00134f
C25490 _0159_ _0497_/a_68_297# 0
C25491 net143 hold70/a_391_47# 0
C25492 _1038_/a_1059_315# _0137_ 0
C25493 _1004_/a_27_47# clknet_1_0__leaf__0460_ 0.00106f
C25494 hold78/a_285_47# net60 0.03843f
C25495 hold23/a_49_47# net10 0.02269f
C25496 net160 _1037_/a_975_413# 0
C25497 _0984_/a_1059_315# _0347_ 0.02083f
C25498 _0217_ _0459_ 0.02557f
C25499 hold72/a_49_47# hold72/a_285_47# 0.22264f
C25500 hold69/a_391_47# _0462_ 0.00756f
C25501 clknet_0__0465_ _0425_ 0
C25502 hold36/a_49_47# _0172_ 0.00305f
C25503 clk input34/a_27_47# 0.00451f
C25504 hold89/a_49_47# _0468_ 0
C25505 hold5/a_391_47# _1042_/a_381_47# 0
C25506 hold65/a_285_47# net65 0.10734f
C25507 _0982_/a_891_413# _0216_ 0
C25508 hold65/a_49_47# _0989_/a_1059_315# 0.00621f
C25509 clknet_1_0__leaf__0462_ _0360_ 0
C25510 VPWR _0466_ 2.41553f
C25511 _1001_/a_193_47# control0.add 0
C25512 acc0.A\[12\] _0285_ 0.00819f
C25513 _0464_ net157 0.6757f
C25514 clkbuf_1_0__f__0457_/a_110_47# _1019_/a_27_47# 0
C25515 _0966_/a_27_47# _0483_ 0.03885f
C25516 _0516_/a_373_47# clknet_1_1__leaf__0465_ 0.0024f
C25517 _0369_ _0391_ 0.0035f
C25518 _0290_ _0350_ 0.3085f
C25519 clknet_0__0457_ _0391_ 0
C25520 hold49/a_391_47# comp0.B\[12\] 0.00773f
C25521 net85 _0306_ 0
C25522 clknet_1_1__leaf__0459_ _0417_ 0.2298f
C25523 comp0.B\[6\] _0175_ 0.09359f
C25524 _0238_ _1006_/a_193_47# 0
C25525 _0384_ _0373_ 0.15542f
C25526 net38 _0419_ 0
C25527 _0649_/a_113_47# _0281_ 0.0096f
C25528 hold22/a_49_47# hold22/a_285_47# 0.22264f
C25529 _0190_ _0990_/a_1059_315# 0
C25530 _0180_ comp0.B\[15\] 0.48509f
C25531 net61 _0449_ 0
C25532 _0261_ acc0.A\[15\] 0.09645f
C25533 _0684_/a_59_75# _1009_/a_27_47# 0
C25534 net89 control0.state\[2\] 0.00516f
C25535 _0473_ net20 0.19476f
C25536 VPWR _0808_/a_266_297# 0.00116f
C25537 _1055_/a_634_159# _0153_ 0
C25538 _0367_ clkbuf_1_0__f__0462_/a_110_47# 0.03165f
C25539 _0998_/a_1059_315# _0219_ 0
C25540 _0218_ _0779_/a_215_47# 0.04984f
C25541 hold77/a_285_47# VPWR 0.31147f
C25542 _0314_ _1025_/a_891_413# 0
C25543 net64 _0621_/a_117_297# 0.00789f
C25544 _0769_/a_81_21# _0769_/a_299_297# 0.08213f
C25545 _0136_ net7 0
C25546 _0621_/a_35_297# _0621_/a_285_297# 0.02504f
C25547 _0581_/a_373_47# _0247_ 0
C25548 _0349_ net239 0
C25549 _0462_ _0617_/a_150_297# 0
C25550 clknet_1_0__leaf__0458_ clkbuf_0__0465_/a_110_47# 0
C25551 _0575_/a_27_297# acc0.A\[23\] 0
C25552 clknet_1_0__leaf__0464_ net134 0.26801f
C25553 net200 net210 0.0017f
C25554 hold53/a_391_47# _0124_ 0
C25555 hold87/a_49_47# hold87/a_285_47# 0.22264f
C25556 hold63/a_391_47# acc0.A\[25\] 0
C25557 _0593_/a_113_47# clknet_1_0__leaf__0460_ 0
C25558 hold68/a_285_47# hold68/a_391_47# 0.41909f
C25559 _0820_/a_215_47# _0292_ 0
C25560 acc0.A\[14\] _0369_ 0.04203f
C25561 _1060_/a_561_413# _0184_ 0
C25562 hold79/a_391_47# _0978_/a_109_297# 0
C25563 _0948_/a_109_297# control0.state\[2\] 0.00188f
C25564 acc0.A\[16\] _1016_/a_891_413# 0.03344f
C25565 _0714_/a_149_47# _0342_ 0.018f
C25566 net182 A[9] 0.00148f
C25567 _0812_/a_510_47# net67 0.00121f
C25568 clknet_1_0__leaf__0463_ _1039_/a_561_413# 0
C25569 clkbuf_1_1__f__0464_/a_110_47# net20 0.00214f
C25570 _1057_/a_1017_47# clknet_1_1__leaf__0465_ 0
C25571 VPWR _1036_/a_592_47# 0
C25572 _1050_/a_193_47# _0524_/a_27_297# 0
C25573 _1050_/a_27_47# _0524_/a_109_297# 0
C25574 input7/a_75_212# net127 0.0214f
C25575 clknet_0__0457_ _0982_/a_381_47# 0
C25576 _1044_/a_466_413# _1044_/a_561_413# 0.00772f
C25577 _1044_/a_634_159# _1044_/a_975_413# 0
C25578 _0654_/a_207_413# _0808_/a_81_21# 0
C25579 _1065_/a_193_47# _0564_/a_68_297# 0.00191f
C25580 comp0.B\[13\] _0954_/a_32_297# 0.06465f
C25581 net158 _0536_/a_51_297# 0.0032f
C25582 net101 _0584_/a_373_47# 0
C25583 _1038_/a_1059_315# comp0.B\[6\] 0.12875f
C25584 _1038_/a_891_413# comp0.B\[5\] 0
C25585 _0966_/a_27_47# control0.count\[1\] 0
C25586 net236 VPWR 0.43009f
C25587 hold41/a_391_47# _1058_/a_193_47# 0.00154f
C25588 hold41/a_285_47# _1058_/a_634_159# 0
C25589 _0212_ _0211_ 0.0759f
C25590 _0815_/a_199_47# _0425_ 0.00151f
C25591 net137 acc0.A\[5\] 0
C25592 hold22/a_285_47# net169 0.00997f
C25593 VPWR _0743_/a_245_297# 0.00512f
C25594 _0183_ net47 0.00314f
C25595 _0217_ _0265_ 0.06806f
C25596 _1058_/a_27_47# _0510_/a_27_297# 0
C25597 net149 _1048_/a_891_413# 0
C25598 net18 _0541_/a_150_297# 0
C25599 _0302_ _0410_ 0
C25600 clknet_1_1__leaf_clk _1065_/a_193_47# 0.1062f
C25601 _0410_ _0795_/a_299_297# 0.00163f
C25602 acc0.A\[1\] _0350_ 0.2709f
C25603 _0999_/a_634_159# _0778_/a_68_297# 0.00106f
C25604 net36 net234 0.0401f
C25605 pp[17] _0345_ 0
C25606 _0985_/a_1059_315# _0629_/a_59_75# 0
C25607 _0381_ _1005_/a_27_47# 0
C25608 _0107_ VPWR 0.37499f
C25609 _1067_/a_891_413# net17 0
C25610 net46 _1023_/a_975_413# 0
C25611 _0216_ _1028_/a_27_47# 0
C25612 _0195_ _1028_/a_634_159# 0.01609f
C25613 hold49/a_49_47# net20 0.04027f
C25614 _1057_/a_634_159# _1057_/a_466_413# 0.23992f
C25615 _1057_/a_193_47# _1057_/a_1059_315# 0.03405f
C25616 _1057_/a_27_47# _1057_/a_891_413# 0.03224f
C25617 _0299_ VPWR 0.65944f
C25618 _0260_ _0446_ 0.07279f
C25619 _0509_/a_27_47# acc0.A\[15\] 0
C25620 clknet_1_1__leaf__0459_ _0669_/a_183_297# 0
C25621 net88 _0165_ 0
C25622 _0579_/a_109_297# clknet_1_0__leaf__0459_ 0.00181f
C25623 _0812_/a_79_21# _0288_ 0.00306f
C25624 pp[17] _0712_/a_381_47# 0
C25625 net225 _1013_/a_193_47# 0
C25626 hold81/a_285_47# _0419_ 0
C25627 VPWR _1064_/a_193_47# 0.30512f
C25628 _0854_/a_79_21# _0116_ 0
C25629 _0432_ clknet_0__0465_ 0.50903f
C25630 net8 clkbuf_0__0463_/a_110_47# 0.12206f
C25631 _0101_ _0467_ 0
C25632 _1059_/a_27_47# _1059_/a_891_413# 0.03224f
C25633 _1059_/a_193_47# _1059_/a_1059_315# 0.03405f
C25634 _1059_/a_634_159# _1059_/a_466_413# 0.23992f
C25635 VPWR _0295_ 1.06848f
C25636 _0343_ _0427_ 0
C25637 comp0.B\[2\] _1065_/a_1059_315# 0
C25638 _0712_/a_79_21# VPWR 0.17708f
C25639 _0179_ _0261_ 0.02022f
C25640 net231 _1062_/a_27_47# 0.00393f
C25641 _0858_/a_27_47# _0146_ 0
C25642 hold96/a_285_47# _0123_ 0
C25643 _0849_/a_79_21# _0082_ 0.05104f
C25644 _0849_/a_510_47# net222 0
C25645 _1015_/a_193_47# _0345_ 0
C25646 hold3/a_391_47# net91 0
C25647 clknet_1_0__leaf__0459_ _0399_ 0.43751f
C25648 clkload4/a_268_47# _0181_ 0.00137f
C25649 _1032_/a_381_47# net202 0.11466f
C25650 _0953_/a_32_297# clknet_1_1__leaf__0457_ 0.01029f
C25651 _0982_/a_891_413# net247 0
C25652 _0713_/a_27_47# _0113_ 0
C25653 _0346_ acc0.A\[13\] 0.02239f
C25654 _0330_ _0729_/a_150_297# 0
C25655 hold37/a_49_47# clknet_1_1__leaf__0464_ 0.04156f
C25656 _1032_/a_381_47# clknet_1_1__leaf__0463_ 0
C25657 _0569_/a_109_47# _0127_ 0
C25658 _0457_ clkbuf_1_1__f__0457_/a_110_47# 0
C25659 _1065_/a_634_159# clkbuf_1_1__f_clk/a_110_47# 0.00238f
C25660 net187 _0721_/a_27_47# 0
C25661 _0481_ _0978_/a_109_297# 0.01339f
C25662 _0179_ _1058_/a_1059_315# 0
C25663 comp0.B\[13\] _0540_/a_245_297# 0.00123f
C25664 _0983_/a_27_47# _0219_ 0
C25665 _0388_ _0773_/a_285_297# 0.08951f
C25666 _0386_ _0773_/a_285_47# 0
C25667 _0180_ net184 0
C25668 net45 _0306_ 0.00574f
C25669 _0783_/a_79_21# _0399_ 0.15204f
C25670 net124 net172 0.02584f
C25671 input33/a_75_212# control0.sh 0
C25672 net33 clknet_1_1__leaf_clk 0.03145f
C25673 net44 hold16/a_391_47# 0
C25674 hold46/a_285_47# _0138_ 0
C25675 _0250_ _0318_ 0
C25676 _0337_ _0705_/a_145_75# 0.00332f
C25677 net47 acc0.A\[15\] 0.04076f
C25678 _0718_/a_129_47# _0336_ 0.00115f
C25679 _0718_/a_285_47# _0220_ 0
C25680 net158 hold46/a_49_47# 0
C25681 hold86/a_49_47# _0846_/a_240_47# 0
C25682 hold86/a_285_47# _0846_/a_149_47# 0
C25683 net55 net57 0.03409f
C25684 acc0.A\[27\] _1028_/a_381_47# 0.00903f
C25685 net40 _0994_/a_27_47# 0
C25686 _0960_/a_27_47# clknet_1_0__leaf_clk 0.10678f
C25687 _0478_ _1069_/a_1059_315# 0
C25688 hold38/a_49_47# _1062_/a_193_47# 0
C25689 hold11/a_391_47# _1046_/a_193_47# 0
C25690 _0707_/a_75_199# _0723_/a_207_413# 0
C25691 _0293_ _0814_/a_181_47# 0
C25692 clknet_0__0461_ hold72/a_285_47# 0.00508f
C25693 hold17/a_285_47# _0466_ 0.05497f
C25694 hold17/a_391_47# _0488_ 0
C25695 net54 _0329_ 0
C25696 _1052_/a_634_159# _0186_ 0.01138f
C25697 hold21/a_391_47# _0180_ 0
C25698 _0836_/a_68_297# _0433_ 0.05687f
C25699 _0267_ _0444_ 0
C25700 _0352_ _1006_/a_975_413# 0.0014f
C25701 _0288_ _0347_ 0.12692f
C25702 _0399_ _0453_ 0
C25703 _0284_ _0993_/a_975_413# 0
C25704 net186 _1033_/a_634_159# 0
C25705 _0179_ _0509_/a_27_47# 0
C25706 _0225_ _0219_ 0.09651f
C25707 _0433_ net212 0
C25708 clkbuf_1_0__f__0464_/a_110_47# _1048_/a_634_159# 0
C25709 _0159_ comp0.B\[8\] 0
C25710 _0305_ _1060_/a_27_47# 0
C25711 _0217_ _0585_/a_109_297# 0.05487f
C25712 _0410_ net6 0
C25713 _0399_ _0794_/a_110_297# 0
C25714 _1014_/a_634_159# clkbuf_0__0457_/a_110_47# 0
C25715 _1056_/a_891_413# _0515_/a_81_21# 0.00142f
C25716 _1056_/a_1059_315# _0515_/a_299_297# 0
C25717 VPWR _0619_/a_68_297# 0.16615f
C25718 net58 net165 0
C25719 _0533_/a_109_297# net8 0.00625f
C25720 net34 clknet_1_0__leaf_clk 0.0508f
C25721 net168 net75 0
C25722 _0349_ _0357_ 0
C25723 _0180_ hold71/a_285_47# 0
C25724 _0182_ hold71/a_391_47# 0.00186f
C25725 _0183_ _1060_/a_1059_315# 0.00195f
C25726 clkbuf_1_1__f__0463_/a_110_47# _0473_ 0.0011f
C25727 _0555_/a_51_297# net28 0.13025f
C25728 acc0.A\[24\] _1007_/a_381_47# 0.00196f
C25729 hold71/a_285_47# net218 0.01097f
C25730 hold32/a_285_47# net179 0.01139f
C25731 comp0.B\[7\] _0206_ 0
C25732 _0123_ _1024_/a_27_47# 0
C25733 clknet_1_0__leaf__0462_ _1022_/a_27_47# 0.08536f
C25734 _0247_ _0347_ 0.08788f
C25735 pp[8] hold34/a_391_47# 0.06045f
C25736 _0616_/a_215_47# _0352_ 0.00328f
C25737 _0383_ _0373_ 0.27299f
C25738 _1031_/a_466_413# _0567_/a_27_297# 0
C25739 _0375_ hold94/a_49_47# 0
C25740 _0234_ hold94/a_391_47# 0.00265f
C25741 hold88/a_391_47# _0369_ 0.00103f
C25742 _0762_/a_79_21# _0352_ 0.1265f
C25743 _0334_ hold62/a_391_47# 0
C25744 net62 _0447_ 0
C25745 VPWR _1023_/a_592_47# 0
C25746 _0546_/a_149_47# net152 0.00734f
C25747 _0546_/a_512_297# net32 0.00106f
C25748 _1047_/a_634_159# clknet_1_1__leaf__0457_ 0.0015f
C25749 net161 _0175_ 0.00336f
C25750 _0190_ _0439_ 0
C25751 _0984_/a_193_47# _0849_/a_79_21# 0
C25752 control0.state\[0\] _0974_/a_79_199# 0
C25753 _0450_ _0447_ 0
C25754 _0607_/a_109_297# _0387_ 0
C25755 control0.state\[1\] _0880_/a_27_47# 0.02712f
C25756 _0991_/a_891_413# _0991_/a_975_413# 0.00851f
C25757 _0991_/a_27_47# net77 0.23091f
C25758 _0991_/a_381_47# _0991_/a_561_413# 0.00123f
C25759 VPWR _0190_ 0.31466f
C25760 net160 _0173_ 0.12031f
C25761 _0210_ _0213_ 0
C25762 _1067_/a_27_47# _0487_ 0
C25763 _0458_ _0195_ 0.00941f
C25764 _0355_ _0345_ 0
C25765 _0467_ net23 0.05415f
C25766 _0440_ clknet_1_1__leaf__0458_ 0.01132f
C25767 _0179_ net47 0.0234f
C25768 hold79/a_391_47# _0480_ 0
C25769 acc0.A\[12\] _0218_ 0
C25770 net78 hold70/a_285_47# 0
C25771 hold58/a_391_47# net25 0.00179f
C25772 _0794_/a_27_47# _0277_ 0.0026f
C25773 _0794_/a_326_47# _0300_ 0.00381f
C25774 _1043_/a_27_47# _0541_/a_68_297# 0
C25775 _0343_ net142 0
C25776 net158 comp0.B\[14\] 0
C25777 net216 _0369_ 0.10254f
C25778 _0814_/a_109_47# clknet_1_1__leaf__0465_ 0
C25779 _0216_ _1029_/a_381_47# 0.01716f
C25780 net97 net115 0
C25781 _0496_/a_27_47# _0176_ 0.17234f
C25782 _0286_ _0808_/a_81_21# 0.06252f
C25783 clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ 1.62961f
C25784 _0563_/a_51_297# _0171_ 0
C25785 _0799_/a_303_47# net5 0.00306f
C25786 _0714_/a_51_297# net59 0
C25787 clknet_1_0__leaf__0457_ hold73/a_285_47# 0.01557f
C25788 net26 _0175_ 0.77348f
C25789 _0982_/a_193_47# acc0.A\[0\] 0.03449f
C25790 _0080_ _1014_/a_1059_315# 0
C25791 _0982_/a_891_413# net100 0
C25792 _1004_/a_1059_315# acc0.A\[23\] 0.00865f
C25793 VPWR _1065_/a_634_159# 0.17789f
C25794 _0600_/a_103_199# _0600_/a_253_297# 0.01483f
C25795 clknet_0__0459_ _0219_ 0.10231f
C25796 hold64/a_49_47# _0391_ 0
C25797 hold64/a_285_47# net223 0
C25798 net7 _1046_/a_381_47# 0
C25799 _0159_ _1046_/a_466_413# 0
C25800 _0195_ _1016_/a_466_413# 0
C25801 net123 _1037_/a_891_413# 0
C25802 clknet_1_0__leaf__0462_ _0124_ 0.01099f
C25803 VPWR _0811_/a_299_297# 0.27668f
C25804 net50 pp[22] 0.00663f
C25805 _0399_ _0996_/a_1017_47# 0.00171f
C25806 net168 net138 0
C25807 _0725_/a_209_297# acc0.A\[29\] 0.00456f
C25808 _0995_/a_27_47# _0995_/a_634_159# 0.14145f
C25809 _0838_/a_109_297# _0465_ 0
C25810 net23 comp0.B\[0\] 0.025f
C25811 _0739_/a_297_297# _0364_ 0.00271f
C25812 _0230_ _0369_ 0
C25813 net77 _0350_ 0.10159f
C25814 net173 comp0.B\[9\] 0.10515f
C25815 _1060_/a_1059_315# acc0.A\[15\] 0.00423f
C25816 hold11/a_391_47# comp0.B\[9\] 0
C25817 _0455_ _0347_ 0
C25818 _0367_ net51 0
C25819 _0467_ net35 0.01024f
C25820 clknet_0__0461_ _0392_ 0
C25821 _1058_/a_1017_47# acc0.A\[10\] 0
C25822 hold9/a_49_47# _1027_/a_27_47# 0
C25823 net36 _0550_/a_51_297# 0
C25824 _0223_ _0350_ 0
C25825 _0218_ _0445_ 0.01508f
C25826 _0398_ _0777_/a_47_47# 0
C25827 net53 _1007_/a_466_413# 0.00177f
C25828 _1070_/a_27_47# _1069_/a_891_413# 0.00368f
C25829 _1070_/a_193_47# _1069_/a_1059_315# 0
C25830 _1070_/a_1059_315# _1069_/a_193_47# 0
C25831 _1070_/a_891_413# _1069_/a_27_47# 0.00368f
C25832 acc0.A\[6\] _0193_ 0.00138f
C25833 acc0.A\[4\] clknet_1_1__leaf__0464_ 0.00397f
C25834 hold64/a_391_47# _0982_/a_1059_315# 0
C25835 _0976_/a_218_47# _0488_ 0
C25836 _0976_/a_535_374# _0466_ 0
C25837 control0.state\[1\] _1062_/a_27_47# 0.02454f
C25838 control0.state\[0\] _1062_/a_193_47# 0.03421f
C25839 _0800_/a_512_297# _0093_ 0
C25840 _0216_ clkbuf_0__0457_/a_110_47# 0.12861f
C25841 _0789_/a_75_199# _0399_ 0
C25842 hold74/a_285_47# net221 0.00962f
C25843 output56/a_27_47# hold95/a_49_47# 0.02626f
C25844 VPWR _0322_ 0.64903f
C25845 pp[8] _0181_ 0.0013f
C25846 _0508_/a_384_47# net229 0
C25847 _1011_/a_634_159# _1011_/a_466_413# 0.23992f
C25848 _1011_/a_193_47# _1011_/a_1059_315# 0.03405f
C25849 _1011_/a_27_47# _1011_/a_891_413# 0.03224f
C25850 _1016_/a_634_159# _0369_ 0.00416f
C25851 net50 _1023_/a_27_47# 0.00194f
C25852 _0170_ _1068_/a_381_47# 0
C25853 hold10/a_49_47# _0171_ 0.00196f
C25854 A[8] _0186_ 0
C25855 net61 _0260_ 0.2359f
C25856 VPWR _0327_ 2.56844f
C25857 _0643_/a_103_199# _0446_ 0
C25858 pp[27] hold62/a_285_47# 0.00731f
C25859 _0481_ _0480_ 0.09904f
C25860 _1034_/a_634_159# net23 0
C25861 pp[9] hold34/a_285_47# 0.03148f
C25862 _0827_/a_27_47# acc0.A\[6\] 0
C25863 _0350_ _1006_/a_1059_315# 0.03198f
C25864 _0217_ net51 0.01892f
C25865 _0295_ _0283_ 0.1705f
C25866 clknet_0__0465_ _0986_/a_381_47# 0.00164f
C25867 _0714_/a_240_47# _0195_ 0.0059f
C25868 _0618_/a_79_21# _0460_ 0.00156f
C25869 VPWR hold51/a_285_47# 0.29622f
C25870 net140 A[7] 0.00792f
C25871 _0296_ _0286_ 0.03523f
C25872 hold55/a_285_47# _1067_/a_891_413# 0
C25873 _0449_ _0431_ 0
C25874 _0752_/a_27_413# hold4/a_391_47# 0
C25875 _1021_/a_27_47# hold73/a_391_47# 0
C25876 _1021_/a_193_47# hold73/a_285_47# 0
C25877 _1020_/a_891_413# VPWR 0.21839f
C25878 _0350_ _0986_/a_1059_315# 0.02339f
C25879 hold33/a_285_47# _0200_ 0
C25880 _0266_ _0345_ 0.00814f
C25881 clkbuf_1_1__f__0462_/a_110_47# net242 0
C25882 _1001_/a_634_159# _0610_/a_59_75# 0
C25883 _1031_/a_193_47# net208 0
C25884 _0971_/a_81_21# _1063_/a_381_47# 0
C25885 _0181_ _1063_/a_27_47# 0
C25886 net188 output67/a_27_47# 0.00242f
C25887 hold41/a_391_47# pp[9] 0.0012f
C25888 _0534_/a_299_297# _0198_ 0
C25889 net83 net41 0.00454f
C25890 clkbuf_0_clk/a_110_47# control0.state\[2\] 0.00948f
C25891 _0955_/a_220_297# comp0.B\[5\] 0.01011f
C25892 VPWR _0515_/a_299_297# 0.20931f
C25893 _0567_/a_109_297# _0345_ 0.00159f
C25894 hold44/a_49_47# acc0.A\[29\] 0.04602f
C25895 _0789_/a_201_297# _0277_ 0.00243f
C25896 _0789_/a_544_297# _0300_ 0.00123f
C25897 _0789_/a_315_47# _0297_ 0.00739f
C25898 _0404_ _0794_/a_326_47# 0.00128f
C25899 _0311_ _0748_/a_81_21# 0.17209f
C25900 _0523_/a_384_47# _0193_ 0
C25901 clknet_1_0__leaf__0463_ clknet_1_0__leaf__0464_ 0
C25902 _0305_ _0748_/a_384_47# 0
C25903 _0680_/a_472_297# _0294_ 0.00427f
C25904 clknet_1_1__leaf__0459_ _0799_/a_209_47# 0
C25905 _1025_/a_1017_47# acc0.A\[25\] 0.00169f
C25906 _0486_ _1063_/a_193_47# 0
C25907 hold33/a_285_47# comp0.B\[8\] 0.04446f
C25908 _0828_/a_113_297# _0989_/a_891_413# 0
C25909 net55 _1010_/a_1059_315# 0
C25910 _0183_ _0848_/a_109_297# 0
C25911 _0170_ _0961_/a_113_297# 0
C25912 hold21/a_49_47# _0152_ 0.0028f
C25913 hold75/a_285_47# _0399_ 0
C25914 net240 _1067_/a_975_413# 0
C25915 _0165_ _1067_/a_891_413# 0.00142f
C25916 net40 _0411_ 0.00123f
C25917 _0181_ _1060_/a_27_47# 0.07783f
C25918 net54 _1008_/a_975_413# 0
C25919 _0503_/a_109_297# _0465_ 0
C25920 _0183_ _0294_ 0.43492f
C25921 hold45/a_285_47# clknet_1_1__leaf__0465_ 0.00488f
C25922 B[12] input32/a_75_212# 0.00253f
C25923 _0516_/a_27_297# _0516_/a_109_47# 0.00393f
C25924 _0173_ acc0.A\[15\] 0
C25925 _1010_/a_27_47# _0352_ 0.03374f
C25926 _1010_/a_466_413# _0347_ 0.01777f
C25927 hold28/a_285_47# acc0.A\[15\] 0
C25928 _1051_/a_466_413# clknet_1_1__leaf__0464_ 0
C25929 _0531_/a_27_297# _1061_/a_1059_315# 0
C25930 clknet_1_1__leaf__0460_ _0730_/a_79_21# 0.01003f
C25931 hold63/a_49_47# net155 0
C25932 hold63/a_285_47# _0195_ 0
C25933 hold63/a_391_47# net210 0.13114f
C25934 _0800_/a_240_47# _0298_ 0
C25935 net55 _1009_/a_891_413# 0.00338f
C25936 _0800_/a_245_297# _0345_ 0
C25937 _0368_ hold90/a_391_47# 0
C25938 _1045_/a_891_413# clknet_1_1__leaf__0464_ 0.00335f
C25939 VPWR _0091_ 0.43436f
C25940 acc0.A\[14\] _0409_ 0
C25941 net141 _0153_ 0
C25942 _1036_/a_1059_315# _1036_/a_891_413# 0.31086f
C25943 _1036_/a_193_47# _1036_/a_975_413# 0
C25944 _1036_/a_466_413# _1036_/a_381_47# 0.03733f
C25945 _0401_ _0986_/a_193_47# 0
C25946 _0244_ _0388_ 0.04002f
C25947 hold97/a_49_47# hold9/a_391_47# 0
C25948 hold26/a_285_47# net180 0.0038f
C25949 control0.sh hold84/a_391_47# 0
C25950 _0994_/a_592_47# acc0.A\[13\] 0
C25951 _0248_ _0772_/a_79_21# 0
C25952 _0347_ _1009_/a_1059_315# 0
C25953 _0523_/a_299_297# _0150_ 0.00112f
C25954 clkload0/X VPWR 0.34223f
C25955 comp0.B\[7\] _0555_/a_240_47# 0
C25956 _0200_ net20 0.00385f
C25957 control0.add _0208_ 0
C25958 _0646_/a_47_47# _0297_ 0.00202f
C25959 clknet_1_0__leaf__0463_ _0553_/a_240_47# 0
C25960 _0176_ net152 0.13171f
C25961 _1041_/a_1059_315# _0204_ 0
C25962 _1041_/a_193_47# net18 0
C25963 _0458_ _1048_/a_193_47# 0
C25964 _0732_/a_80_21# _1007_/a_27_47# 0
C25965 net24 net201 0
C25966 clkbuf_1_1__f__0459_/a_110_47# _0301_ 0.03997f
C25967 _0317_ _0328_ 0.03542f
C25968 _0796_/a_510_47# acc0.A\[15\] 0.00102f
C25969 _1065_/a_891_413# _0215_ 0
C25970 output37/a_27_47# _0188_ 0
C25971 pp[0] input29/a_75_212# 0.00695f
C25972 _0529_/a_109_297# net10 0.00698f
C25973 _0236_ _0369_ 0.02447f
C25974 hold69/a_391_47# _0312_ 0.00133f
C25975 _0483_ _0981_/a_27_297# 0.11241f
C25976 _0996_/a_1059_315# _0219_ 0
C25977 hold13/a_285_47# clkbuf_1_1__f__0463_/a_110_47# 0
C25978 hold49/a_285_47# _0203_ 0
C25979 VPWR _0306_ 0.67647f
C25980 hold33/a_49_47# _1046_/a_1059_315# 0.00115f
C25981 _0985_/a_1017_47# _0465_ 0
C25982 _0181_ _1062_/a_1059_315# 0
C25983 _0163_ _1062_/a_634_159# 0
C25984 _0576_/a_27_297# VPWR 0.24823f
C25985 clknet_1_0__leaf__0462_ _1024_/a_466_413# 0.00271f
C25986 _0467_ _1063_/a_466_413# 0.01275f
C25987 _1058_/a_634_159# net4 0.0407f
C25988 _1058_/a_27_47# _0187_ 0
C25989 _0992_/a_193_47# _0282_ 0
C25990 _0596_/a_59_75# _0760_/a_47_47# 0
C25991 _0742_/a_299_297# net51 0
C25992 _0869_/a_27_47# _0242_ 0
C25993 _0415_ net39 0.0984f
C25994 _1052_/a_1059_315# _0518_/a_27_297# 0.01884f
C25995 net36 _1038_/a_1017_47# 0
C25996 output36/a_27_47# net124 0.01236f
C25997 pp[0] _1038_/a_975_413# 0
C25998 _0218_ net42 0.29404f
C25999 _0294_ acc0.A\[15\] 0.03979f
C26000 _0329_ net227 0
C26001 net224 hold77/a_391_47# 0.1316f
C26002 _1012_/a_193_47# net239 0
C26003 _0428_ _0990_/a_891_413# 0.03876f
C26004 _0663_/a_27_413# net67 0
C26005 net111 hold8/a_391_47# 0
C26006 _0195_ net114 0.00768f
C26007 _0570_/a_109_297# hold8/a_391_47# 0
C26008 _0736_/a_311_297# _0107_ 0.004f
C26009 _1057_/a_634_159# net189 0.03816f
C26010 B[13] _1042_/a_592_47# 0
C26011 pp[30] _0352_ 0
C26012 _0216_ _0534_/a_299_297# 0
C26013 _0111_ _1013_/a_1017_47# 0
C26014 _0250_ _1007_/a_27_47# 0
C26015 _0179_ hold28/a_285_47# 0.08141f
C26016 _0189_ acc0.A\[9\] 0.0094f
C26017 _0216_ hold62/a_285_47# 0
C26018 _0093_ _0995_/a_193_47# 0.22816f
C26019 _0789_/a_75_199# _0299_ 0.10228f
C26020 _0789_/a_201_297# _0298_ 0.03027f
C26021 _0626_/a_68_297# _0636_/a_59_75# 0
C26022 _1059_/a_466_413# net145 0
C26023 _0754_/a_51_297# _0754_/a_245_297# 0.01218f
C26024 _1041_/a_891_413# _1041_/a_1017_47# 0.00617f
C26025 _0693_/a_150_297# net52 0
C26026 _0528_/a_299_297# _0148_ 0.00103f
C26027 _0174_ clknet_1_1__leaf__0457_ 0.16816f
C26028 net220 _0381_ 0.00238f
C26029 _0470_ _0951_/a_109_93# 0
C26030 _0713_/a_27_47# _0345_ 0.3368f
C26031 _0510_/a_109_47# _0186_ 0.0034f
C26032 _0433_ _0989_/a_891_413# 0
C26033 _0221_ net227 0
C26034 _1055_/a_193_47# clknet_1_1__leaf__0465_ 0.04086f
C26035 _0811_/a_299_297# _0283_ 0.0648f
C26036 _0181_ _1047_/a_381_47# 0
C26037 _0710_/a_109_47# _0340_ 0.00237f
C26038 _0779_/a_297_297# _0347_ 0.00188f
C26039 _0176_ _1042_/a_466_413# 0
C26040 _0323_ clkbuf_0__0462_/a_110_47# 0.00334f
C26041 _0443_ _0986_/a_193_47# 0.00243f
C26042 _0432_ _0986_/a_27_47# 0
C26043 _0352_ _0771_/a_215_297# 0.07604f
C26044 net168 hold83/a_285_47# 0.0696f
C26045 clknet_0__0458_ _0271_ 0.00474f
C26046 _1002_/a_1059_315# _0578_/a_27_297# 0
C26047 net193 net20 0.08649f
C26048 net214 _0088_ 0
C26049 _0672_/a_79_21# _0296_ 0.05685f
C26050 _0383_ _0761_/a_113_47# 0.00973f
C26051 _0891_/a_27_47# VPWR 0.19902f
C26052 pp[16] hold98/a_285_47# 0.00387f
C26053 _0992_/a_27_47# _0281_ 0
C26054 _0369_ _0422_ 0.15874f
C26055 _0717_/a_80_21# _0723_/a_27_413# 0.0023f
C26056 clkbuf_1_0__f__0458_/a_110_47# _0458_ 0
C26057 _0536_/a_245_297# net22 0.00277f
C26058 control0.state\[0\] hold85/a_49_47# 0.00102f
C26059 input10/a_75_212# A[2] 0.00628f
C26060 A[3] input9/a_27_47# 0
C26061 _0372_ _0218_ 0
C26062 _0974_/a_222_93# _1068_/a_27_47# 0
C26063 _0974_/a_79_199# _1068_/a_193_47# 0.00129f
C26064 acc0.A\[27\] acc0.A\[28\] 0.0073f
C26065 _1054_/a_891_413# _0087_ 0
C26066 VPWR _1008_/a_561_413# 0.00355f
C26067 clkbuf_1_0__f__0463_/a_110_47# _0205_ 0
C26068 _0981_/a_109_297# clkbuf_1_0__f_clk/a_110_47# 0
C26069 _0476_ hold58/a_285_47# 0
C26070 hold11/a_285_47# net132 0.01211f
C26071 net158 _1046_/a_561_413# 0
C26072 _0335_ _0723_/a_297_47# 0
C26073 _0338_ _0723_/a_207_413# 0
C26074 _0343_ _0988_/a_27_47# 0
C26075 _0891_/a_27_47# _1015_/a_466_413# 0
C26076 _1028_/a_193_47# _1027_/a_1059_315# 0
C26077 _1028_/a_27_47# _1027_/a_891_413# 0.01107f
C26078 _1020_/a_891_413# clknet_1_0__leaf__0459_ 0.00914f
C26079 output55/a_27_47# _1011_/a_193_47# 0
C26080 comp0.B\[2\] net24 0.0215f
C26081 _0195_ _0365_ 0.00371f
C26082 net36 _0913_/a_27_47# 0
C26083 net22 _0547_/a_68_297# 0
C26084 _0179_ _0294_ 0.08417f
C26085 pp[27] _0350_ 0
C26086 net239 clknet_1_1__leaf__0461_ 0
C26087 _0180_ _0845_/a_193_297# 0
C26088 _0217_ _0178_ 0.01599f
C26089 clknet_1_0__leaf__0458_ _0180_ 0
C26090 input14/a_75_212# A[7] 0.21986f
C26091 net120 net185 0
C26092 _0341_ _1013_/a_634_159# 0
C26093 _0340_ _1013_/a_193_47# 0
C26094 net186 net119 0
C26095 _0269_ _0449_ 0.00119f
C26096 clknet_1_0__leaf__0458_ net218 0.00108f
C26097 _0478_ _0974_/a_79_199# 0
C26098 net144 _0513_/a_384_47# 0
C26099 _0469_ _0468_ 0.01923f
C26100 clknet_1_0__leaf__0463_ _0536_/a_245_297# 0
C26101 _0218_ hold40/a_49_47# 0.00403f
C26102 _0762_/a_79_21# _0237_ 0
C26103 _0369_ _0760_/a_377_297# 0.00149f
C26104 clkbuf_1_0__f__0464_/a_110_47# net134 0
C26105 _0699_/a_150_297# _0331_ 0
C26106 _0995_/a_27_47# _0345_ 0
C26107 _0222_ _0600_/a_103_199# 0
C26108 _1010_/a_193_47# hold95/a_391_47# 0
C26109 _0361_ hold90/a_49_47# 0.02791f
C26110 _0676_/a_113_47# _0218_ 0
C26111 _1030_/a_193_47# net239 0
C26112 net108 _0577_/a_27_297# 0
C26113 clknet_1_0__leaf__0462_ _0577_/a_109_47# 0.00105f
C26114 _1031_/a_27_47# _1031_/a_634_159# 0.14145f
C26115 clknet_1_0__leaf__0463_ _0547_/a_68_297# 0.02995f
C26116 hold19/a_391_47# _0181_ 0
C26117 pp[18] _0344_ 0
C26118 _0517_/a_81_21# _0186_ 0
C26119 net45 _0778_/a_68_297# 0.00216f
C26120 VPWR _0563_/a_240_47# 0.00143f
C26121 _0121_ hold96/a_285_47# 0.00186f
C26122 hold26/a_391_47# _0545_/a_68_297# 0
C26123 control0.state\[1\] _1063_/a_561_413# 0.002f
C26124 hold44/a_285_47# hold44/a_391_47# 0.41909f
C26125 _1005_/a_634_159# _1005_/a_975_413# 0
C26126 _1005_/a_466_413# _1005_/a_561_413# 0.00772f
C26127 _1067_/a_1059_315# _0352_ 0
C26128 net178 hold88/a_49_47# 0
C26129 _0534_/a_299_297# net247 0.05462f
C26130 VPWR net192 0.17002f
C26131 net32 _0139_ 0.02514f
C26132 _0984_/a_634_159# _0082_ 0.05333f
C26133 _0984_/a_891_413# net222 0.00757f
C26134 _1066_/a_193_47# _1062_/a_193_47# 0.00464f
C26135 net9 A[3] 0.00101f
C26136 _0646_/a_47_47# _0646_/a_377_297# 0.00899f
C26137 _0195_ _0408_ 0
C26138 _1013_/a_193_47# _1013_/a_381_47# 0.09799f
C26139 _1013_/a_634_159# _1013_/a_891_413# 0.03684f
C26140 _1013_/a_27_47# _1013_/a_561_413# 0.0027f
C26141 clknet_1_0__leaf__0465_ net7 0
C26142 VPWR _0527_/a_109_297# 0.19641f
C26143 _1002_/a_193_47# _1002_/a_634_159# 0.11072f
C26144 _1002_/a_27_47# _1002_/a_466_413# 0.27314f
C26145 VPWR _0346_ 4.67401f
C26146 hold64/a_285_47# clkbuf_0__0457_/a_110_47# 0.00254f
C26147 _1027_/a_27_47# _0739_/a_79_21# 0
C26148 hold26/a_49_47# hold26/a_391_47# 0.00188f
C26149 clkbuf_0__0463_/a_110_47# _0492_/a_27_47# 0.0244f
C26150 _0461_ _0526_/a_27_47# 0.00527f
C26151 _0339_ _0352_ 0
C26152 _1027_/a_193_47# _0347_ 0.00103f
C26153 _0749_/a_81_21# _0373_ 0.12206f
C26154 net205 net204 0.00139f
C26155 _0367_ _0324_ 0
C26156 _0252_ _0438_ 0.00168f
C26157 _0985_/a_975_413# _0261_ 0
C26158 _0607_/a_109_297# acc0.A\[16\] 0.0015f
C26159 _0283_ _0091_ 0
C26160 net165 _1060_/a_466_413# 0
C26161 clknet_0_clk hold84/a_49_47# 0
C26162 comp0.B\[4\] net29 0
C26163 input30/a_75_212# A[15] 0.00103f
C26164 B[7] input7/a_75_212# 0
C26165 VPWR net65 0.60101f
C26166 hold35/a_49_47# _1055_/a_27_47# 0
C26167 clknet_1_1__leaf__0459_ _0992_/a_1017_47# 0
C26168 VPWR _0989_/a_466_413# 0.25084f
C26169 hold32/a_391_47# pp[9] 0
C26170 _0108_ _0317_ 0
C26171 _0180_ _0525_/a_299_297# 0.01206f
C26172 _0174_ net19 0.01799f
C26173 _1038_/a_1059_315# _1040_/a_466_413# 0
C26174 _1038_/a_891_413# _1040_/a_634_159# 0
C26175 clknet_1_0__leaf__0459_ _0306_ 0
C26176 _0217_ _1019_/a_27_47# 0.01912f
C26177 VPWR _0992_/a_466_413# 0.24755f
C26178 _0260_ _0431_ 0.18245f
C26179 _0734_/a_47_47# _0361_ 0.3737f
C26180 _0195_ net166 0
C26181 VPWR hold94/a_49_47# 0.26209f
C26182 _0462_ _0219_ 0.05836f
C26183 _0719_/a_27_47# _0242_ 0.02986f
C26184 _0995_/a_891_413# _0995_/a_975_413# 0.00851f
C26185 _0995_/a_381_47# _0995_/a_561_413# 0.00123f
C26186 _0765_/a_79_21# _0765_/a_215_47# 0.04584f
C26187 hold65/a_49_47# _0186_ 0
C26188 _0346_ _0654_/a_27_413# 0.01832f
C26189 net10 net170 0.51377f
C26190 hold46/a_285_47# clknet_1_0__leaf__0463_ 0
C26191 VPWR _0935_/a_27_47# 0.20068f
C26192 output56/a_27_47# _1011_/a_27_47# 0
C26193 _0437_ _0829_/a_27_47# 0.05636f
C26194 VPWR _1061_/a_193_47# 0.32728f
C26195 _0820_/a_215_47# clkbuf_1_1__f__0465_/a_110_47# 0
C26196 clknet_1_1__leaf__0459_ _0668_/a_79_21# 0.00366f
C26197 _0983_/a_381_47# _0346_ 0
C26198 _0732_/a_209_297# _0460_ 0
C26199 net82 _0507_/a_109_297# 0
C26200 _0501_/a_27_47# net8 0.03684f
C26201 _0783_/a_79_21# _0306_ 0.00426f
C26202 _0369_ _0370_ 0
C26203 _1070_/a_891_413# _0489_ 0
C26204 acc0.A\[12\] net228 0
C26205 _0534_/a_81_21# _1048_/a_1059_315# 0
C26206 _1017_/a_1059_315# _0675_/a_68_297# 0
C26207 _1034_/a_634_159# _0213_ 0.00279f
C26208 _1034_/a_193_47# _0173_ 0.03466f
C26209 _1034_/a_891_413# _0561_/a_240_47# 0
C26210 _0629_/a_59_75# VPWR 0.22493f
C26211 _0183_ _0581_/a_109_297# 0.00929f
C26212 net36 _0172_ 0.05249f
C26213 _1000_/a_27_47# _0775_/a_79_21# 0
C26214 clknet_0_clk _1065_/a_381_47# 0
C26215 _0096_ _0395_ 0
C26216 _0139_ _1042_/a_1059_315# 0
C26217 net32 _1042_/a_561_413# 0.0021f
C26218 input4/a_75_212# net192 0
C26219 _1018_/a_891_413# _0459_ 0.00103f
C26220 _0251_ _0622_/a_109_47# 0
C26221 net53 _0105_ 0
C26222 _0369_ acc0.A\[8\] 0.27766f
C26223 hold86/a_285_47# acc0.A\[15\] 0.00705f
C26224 _1019_/a_1059_315# _0580_/a_27_297# 0
C26225 _0227_ net213 0.00121f
C26226 net1 net23 0
C26227 _1070_/a_466_413# clknet_1_0__leaf_clk 0
C26228 VPWR _1069_/a_1059_315# 0.39173f
C26229 net48 _0346_ 0.00919f
C26230 _0982_/a_561_413# _0183_ 0
C26231 _1034_/a_1059_315# _0475_ 0
C26232 _1034_/a_891_413# _0472_ 0
C26233 _0399_ _0345_ 0.36783f
C26234 _0343_ _0459_ 0.10111f
C26235 _0476_ _0134_ 0
C26236 _1052_/a_1059_315# _0987_/a_27_47# 0
C26237 _0762_/a_79_21# _1005_/a_27_47# 0
C26238 _1011_/a_466_413# net97 0
C26239 _0275_ net62 0.57136f
C26240 _0985_/a_466_413# _0186_ 0.01078f
C26241 net55 clkbuf_1_1__f__0460_/a_110_47# 0.21648f
C26242 net81 _0405_ 0
C26243 _0133_ _1034_/a_592_47# 0
C26244 _1055_/a_27_47# A[9] 0
C26245 _0644_/a_47_47# hold91/a_391_47# 0
C26246 net243 _0574_/a_27_297# 0
C26247 clkbuf_0__0462_/a_110_47# _0686_/a_27_53# 0
C26248 net176 acc0.A\[23\] 0.22998f
C26249 _0216_ _0350_ 0.37024f
C26250 _1006_/a_193_47# _1006_/a_891_413# 0.19489f
C26251 _1006_/a_27_47# _1006_/a_381_47# 0.06222f
C26252 _1006_/a_634_159# _1006_/a_1059_315# 0
C26253 _0182_ _0532_/a_384_47# 0
C26254 _0538_/a_149_47# VPWR 0
C26255 clkload2/Y net170 0
C26256 _0532_/a_299_297# net218 0.05953f
C26257 _0993_/a_193_47# _0807_/a_68_297# 0
C26258 _1049_/a_27_47# _0186_ 0
C26259 _0139_ net10 0.32635f
C26260 acc0.A\[1\] _1014_/a_27_47# 0
C26261 _0111_ _0216_ 0
C26262 _0305_ _0094_ 0
C26263 _0984_/a_193_47# _0984_/a_634_159# 0.11072f
C26264 _0984_/a_27_47# _0984_/a_466_413# 0.27314f
C26265 net181 input16/a_75_212# 0
C26266 net21 _1043_/a_27_47# 0
C26267 _0352_ _1026_/a_193_47# 0
C26268 _0231_ _0328_ 0.00195f
C26269 clknet_1_0__leaf__0462_ _0756_/a_285_47# 0.00289f
C26270 net39 _0347_ 0.0626f
C26271 _1031_/a_27_47# _0345_ 0
C26272 _0808_/a_81_21# _0808_/a_585_47# 0.00695f
C26273 _0808_/a_266_297# _0808_/a_266_47# 0
C26274 _1055_/a_592_47# VPWR 0
C26275 net79 _0808_/a_81_21# 0
C26276 net182 _0515_/a_299_297# 0
C26277 _0399_ hold2/a_49_47# 0
C26278 _1018_/a_381_47# clknet_1_0__leaf__0461_ 0.00338f
C26279 _0390_ _0346_ 0
C26280 hold52/a_285_47# net50 0
C26281 _0352_ _1024_/a_891_413# 0
C26282 net150 net49 0.39871f
C26283 _1003_/a_975_413# VPWR 0.00487f
C26284 _0251_ _0436_ 0.01702f
C26285 hold65/a_285_47# _0253_ 0.00193f
C26286 _0440_ _0218_ 0.00707f
C26287 net9 net154 0
C26288 _0235_ net51 0
C26289 _0955_/a_32_297# hold84/a_391_47# 0
C26290 pp[26] net113 0
C26291 _1039_/a_193_47# VPWR 0.28535f
C26292 _0231_ _0599_/a_113_47# 0.00998f
C26293 _0195_ _0632_/a_113_47# 0
C26294 net35 net1 0
C26295 _0712_/a_79_21# _1031_/a_634_159# 0
C26296 _0986_/a_193_47# _0986_/a_891_413# 0.19489f
C26297 _0986_/a_27_47# _0986_/a_381_47# 0.06222f
C26298 _0986_/a_634_159# _0986_/a_1059_315# 0
C26299 net149 _0181_ 0.66437f
C26300 net148 _0987_/a_381_47# 0.00229f
C26301 _0194_ _0987_/a_193_47# 0
C26302 _0297_ _0219_ 0
C26303 _0566_/a_27_47# control0.reset 0
C26304 _1017_/a_466_413# _0181_ 0
C26305 hold43/a_285_47# _0569_/a_27_297# 0.00327f
C26306 _1023_/a_466_413# _1023_/a_381_47# 0.03733f
C26307 _1023_/a_193_47# _1023_/a_975_413# 0
C26308 _1023_/a_1059_315# _1023_/a_891_413# 0.31086f
C26309 _0627_/a_109_93# _0271_ 0
C26310 _0221_ net208 0
C26311 B[14] net153 0
C26312 net22 net127 0.07175f
C26313 _1042_/a_634_159# _1042_/a_592_47# 0
C26314 hold59/a_285_47# hold59/a_391_47# 0.41909f
C26315 _1019_/a_193_47# control0.add 0
C26316 net54 _0696_/a_109_297# 0
C26317 _1003_/a_193_47# clknet_0_clk 0
C26318 control0.state\[0\] net17 0.03004f
C26319 _0516_/a_109_47# _0190_ 0
C26320 _1037_/a_891_413# _0209_ 0.00185f
C26321 _0425_ _0288_ 0.00325f
C26322 _1033_/a_27_47# _0181_ 0
C26323 net50 net52 0.05406f
C26324 clknet_1_1__leaf__0464_ _1044_/a_1059_315# 0.04236f
C26325 _1011_/a_1059_315# _0707_/a_75_199# 0
C26326 _1045_/a_1059_315# _0202_ 0
C26327 _1045_/a_193_47# net20 0.03582f
C26328 net9 _0465_ 0.00339f
C26329 _1017_/a_891_413# _0307_ 0
C26330 hold68/a_49_47# acc0.A\[23\] 0.31291f
C26331 _0149_ clknet_1_1__leaf__0464_ 0.00748f
C26332 hold86/a_285_47# _0179_ 0
C26333 _0412_ _0219_ 0.14894f
C26334 _0347_ _0444_ 0.0959f
C26335 clknet_0__0458_ clknet_1_0__leaf__0465_ 0.00224f
C26336 _1036_/a_381_47# net161 0.14335f
C26337 _1036_/a_466_413# comp0.B\[4\] 0
C26338 _0625_/a_145_75# _0442_ 0
C26339 _0466_ _1064_/a_466_413# 0
C26340 _0195_ _0528_/a_81_21# 0
C26341 acc0.A\[2\] net9 0
C26342 hold16/a_49_47# _1031_/a_27_47# 0.01435f
C26343 net10 _1042_/a_561_413# 0
C26344 _0498_/a_51_297# _0176_ 0
C26345 hold18/a_391_47# acc0.A\[1\] 0
C26346 hold18/a_285_47# _0182_ 0
C26347 _0230_ hold66/a_391_47# 0
C26348 _0742_/a_299_297# _0324_ 0
C26349 clknet_1_0__leaf__0463_ net127 0.15837f
C26350 _0984_/a_634_159# net145 0
C26351 _0750_/a_27_47# _0374_ 0.08788f
C26352 _1059_/a_27_47# _0506_/a_299_297# 0.02367f
C26353 net64 _0369_ 0.0308f
C26354 _0808_/a_266_297# _0345_ 0
C26355 _0621_/a_117_297# _0369_ 0
C26356 _1057_/a_1059_315# _0511_/a_81_21# 0.01733f
C26357 _0746_/a_81_21# _0462_ 0.0141f
C26358 pp[29] _1011_/a_634_159# 0
C26359 _0476_ _0554_/a_68_297# 0
C26360 _0992_/a_381_47# clknet_1_1__leaf__0465_ 0
C26361 VPWR _1040_/a_592_47# 0
C26362 _0280_ acc0.A\[10\] 0
C26363 _0997_/a_27_47# _0407_ 0.00777f
C26364 _0560_/a_68_297# _0560_/a_150_297# 0.00477f
C26365 net240 _0971_/a_299_297# 0
C26366 acc0.A\[4\] net148 0.13694f
C26367 clknet_1_0__leaf__0459_ _0346_ 0.05271f
C26368 _0423_ _0369_ 0
C26369 _0367_ _0347_ 0.00157f
C26370 _0743_/a_51_297# _0743_/a_240_47# 0.03076f
C26371 _0998_/a_193_47# _0459_ 0
C26372 hold88/a_285_47# pp[1] 0
C26373 _0483_ _0170_ 0.10706f
C26374 _0777_/a_47_47# _0308_ 0.01318f
C26375 _1002_/a_193_47# net220 0
C26376 _1002_/a_27_47# _0385_ 0
C26377 _0305_ _0393_ 0
C26378 _1054_/a_634_159# net11 0
C26379 hold85/a_285_47# _1066_/a_27_47# 0.00754f
C26380 clknet_1_0__leaf__0462_ _0122_ 0.00662f
C26381 _0467_ _0161_ 0.18576f
C26382 net144 net4 0.22699f
C26383 hold34/a_391_47# A[10] 0.02543f
C26384 pp[9] _0153_ 0.00107f
C26385 _0251_ _1054_/a_1059_315# 0
C26386 net247 _0350_ 0.19334f
C26387 _0099_ hold40/a_49_47# 0
C26388 _0391_ hold40/a_391_47# 0
C26389 _0195_ acc0.A\[1\] 0.15842f
C26390 hold19/a_49_47# _0114_ 0.31334f
C26391 _1052_/a_1059_315# _0191_ 0.00249f
C26392 net117 _0195_ 0.00856f
C26393 _0999_/a_891_413# _0218_ 0.05553f
C26394 _0856_/a_510_47# acc0.A\[1\] 0.00458f
C26395 _0346_ _0283_ 0.06328f
C26396 clknet_1_0__leaf__0464_ _1049_/a_381_47# 0.00393f
C26397 _1058_/a_891_413# acc0.A\[11\] 0
C26398 _0463_ net247 0
C26399 hold89/a_49_47# _0480_ 0
C26400 _0278_ _0403_ 0
C26401 VPWR _1035_/a_1059_315# 0.40716f
C26402 A[10] _0510_/a_27_297# 0
C26403 _1000_/a_193_47# net223 0.00149f
C26404 _1001_/a_634_159# net45 0
C26405 _0217_ _0347_ 0.11441f
C26406 net145 _0157_ 0.09303f
C26407 _0299_ _0345_ 0
C26408 _0754_/a_245_297# _0219_ 0
C26409 _0467_ _1033_/a_466_413# 0
C26410 _0260_ _0269_ 0.26228f
C26411 _0754_/a_149_47# _0377_ 0.00697f
C26412 _0272_ _0256_ 0
C26413 _0274_ _0270_ 0
C26414 _0982_/a_466_413# _0181_ 0.03502f
C26415 acc0.A\[20\] net46 0
C26416 _0343_ _0220_ 0.15502f
C26417 comp0.B\[0\] _0161_ 0.10046f
C26418 _0179_ _1053_/a_466_413# 0
C26419 _0853_/a_68_297# _0452_ 0
C26420 _0236_ _0764_/a_384_47# 0
C26421 _0992_/a_634_159# _0286_ 0
C26422 _0992_/a_466_413# _0283_ 0
C26423 clknet_0_clk _0471_ 0.0017f
C26424 _1056_/a_193_47# pp[8] 0
C26425 _0844_/a_382_297# _0350_ 0
C26426 net215 clknet_1_0__leaf__0460_ 0
C26427 _0453_ _0346_ 0.01539f
C26428 _0295_ _0345_ 0.08791f
C26429 _1055_/a_27_47# _0516_/a_27_297# 0
C26430 _1064_/a_27_47# _1064_/a_1059_315# 0.04861f
C26431 _1064_/a_193_47# _1064_/a_466_413# 0.08301f
C26432 _0643_/a_103_199# _0431_ 0.00813f
C26433 _1018_/a_27_47# net149 0
C26434 _0752_/a_300_297# _0750_/a_27_47# 0
C26435 clknet_1_1__leaf__0459_ _0786_/a_472_297# 0.00172f
C26436 net228 net42 0
C26437 _1054_/a_634_159# hold7/a_391_47# 0
C26438 _1054_/a_466_413# hold7/a_285_47# 0
C26439 _1000_/a_27_47# _0581_/a_27_297# 0
C26440 clk A[0] 0.02967f
C26441 clknet_1_0__leaf_clk _0166_ 0.03337f
C26442 net204 net160 0
C26443 _0255_ _0826_/a_27_53# 0.12354f
C26444 VPWR _0778_/a_68_297# 0.16934f
C26445 clknet_1_1__leaf__0460_ net93 0.10219f
C26446 _0712_/a_79_21# _0712_/a_381_47# 0.00247f
C26447 _0574_/a_27_297# _0366_ 0
C26448 net1 _1063_/a_466_413# 0
C26449 _1051_/a_27_47# net12 0.00863f
C26450 _1051_/a_466_413# net148 0
C26451 _0819_/a_81_21# _0399_ 0
C26452 _1033_/a_466_413# comp0.B\[0\] 0
C26453 _1053_/a_592_47# net12 0
C26454 _0348_ _0723_/a_207_413# 0
C26455 _0852_/a_35_297# acc0.A\[1\] 0.00319f
C26456 clknet_1_1__leaf_clk _0880_/a_27_47# 0
C26457 _0181_ _0094_ 0
C26458 _0568_/a_109_297# clknet_1_1__leaf__0462_ 0
C26459 _0343_ _1060_/a_381_47# 0
C26460 _0520_/a_27_297# VPWR 0.18143f
C26461 net159 _1068_/a_891_413# 0
C26462 control0.state\[0\] _0970_/a_285_47# 0.0024f
C26463 net34 _0970_/a_27_297# 0.06904f
C26464 hold19/a_391_47# clknet_1_1__leaf__0461_ 0
C26465 clknet_1_0__leaf__0458_ _0854_/a_510_47# 0
C26466 clknet_0__0465_ _0841_/a_215_47# 0.00111f
C26467 clkbuf_0__0465_/a_110_47# _0444_ 0.00148f
C26468 _0946_/a_30_53# control0.state\[2\] 0.06696f
C26469 _0118_ net87 0.02416f
C26470 _0576_/a_109_47# net50 0.00121f
C26471 _0477_ _0951_/a_368_53# 0
C26472 _0399_ net212 0.12041f
C26473 _0183_ _0458_ 0
C26474 _0737_/a_35_297# _0360_ 0.20474f
C26475 _0157_ net67 0
C26476 A[10] _0181_ 0.00963f
C26477 _0259_ _0990_/a_1059_315# 0
C26478 net45 net221 0.00317f
C26479 VPWR clkbuf_0__0464_/a_110_47# 1.2293f
C26480 _0697_/a_80_21# _0322_ 0.16715f
C26481 _0350_ _0841_/a_79_21# 0
C26482 _0216_ _0244_ 0.13471f
C26483 clknet_1_1__leaf__0460_ _0294_ 0.08918f
C26484 _0565_/a_240_47# _0173_ 0.02408f
C26485 net157 _1061_/a_561_413# 0
C26486 net56 _0322_ 0
C26487 _0989_/a_193_47# acc0.A\[6\] 0
C26488 hold1/a_285_47# acc0.A\[6\] 0
C26489 _0697_/a_80_21# _0327_ 0
C26490 _0857_/a_27_47# clknet_1_1__leaf_clk 0.19588f
C26491 hold70/a_391_47# net37 0
C26492 _0420_ hold81/a_285_47# 0.00457f
C26493 _0712_/a_79_21# hold16/a_49_47# 0
C26494 _0830_/a_79_21# _0830_/a_297_297# 0.01735f
C26495 _1056_/a_193_47# _0988_/a_891_413# 0
C26496 _0399_ _0791_/a_113_297# 0
C26497 comp0.B\[4\] comp0.B\[6\] 0
C26498 net56 _0327_ 0.01515f
C26499 _0151_ _0179_ 0.00603f
C26500 _0695_/a_217_297# _0327_ 0.00405f
C26501 input31/a_75_212# net31 0.10986f
C26502 _1037_/a_193_47# VPWR 0.32201f
C26503 _0837_/a_81_21# acc0.A\[4\] 0.00264f
C26504 _0183_ _1016_/a_466_413# 0
C26505 _0228_ _0377_ 0
C26506 comp0.B\[10\] net18 0.02911f
C26507 net175 _1047_/a_27_47# 0
C26508 _0531_/a_27_297# _1047_/a_381_47# 0
C26509 _1031_/a_891_413# _1031_/a_975_413# 0.00851f
C26510 _1031_/a_381_47# _1031_/a_561_413# 0.00123f
C26511 _0289_ _0786_/a_217_297# 0.0027f
C26512 _0287_ _0786_/a_80_21# 0.00217f
C26513 net100 _0350_ 0
C26514 _0121_ _0756_/a_47_47# 0.00847f
C26515 _1041_/a_1059_315# VPWR 0.39299f
C26516 clknet_0__0458_ net76 0.00128f
C26517 _0252_ _0829_/a_27_47# 0
C26518 net207 acc0.A\[0\] 0
C26519 _1022_/a_193_47# _1005_/a_193_47# 0
C26520 _0645_/a_285_47# acc0.A\[14\] 0.03532f
C26521 pp[15] _0995_/a_466_413# 0.00377f
C26522 _0722_/a_79_21# _0351_ 0.18838f
C26523 net145 acc0.A\[9\] 0
C26524 net17 _0565_/a_51_297# 0.12032f
C26525 _0742_/a_299_297# _0347_ 0
C26526 _0386_ _0240_ 0.00141f
C26527 _0326_ _0366_ 0
C26528 net70 _0082_ 0.00867f
C26529 clknet_1_1__leaf_clk _1062_/a_27_47# 0.33441f
C26530 _1056_/a_27_47# pp[9] 0
C26531 _1060_/a_891_413# net5 0
C26532 _1060_/a_466_413# _0185_ 0
C26533 _0158_ _0507_/a_27_297# 0
C26534 _1020_/a_27_47# _1020_/a_193_47# 0.9705f
C26535 _1002_/a_1059_315# _1002_/a_1017_47# 0
C26536 _1002_/a_193_47# net88 0.04879f
C26537 _1002_/a_27_47# _0100_ 0.09088f
C26538 _0792_/a_80_21# net42 0.0022f
C26539 _0405_ _0790_/a_35_297# 0
C26540 pp[16] output45/a_27_47# 0.00249f
C26541 _1027_/a_466_413# _0365_ 0
C26542 _1027_/a_193_47# _0106_ 0
C26543 _1021_/a_891_413# net1 0.01747f
C26544 _0984_/a_1017_47# clknet_1_0__leaf__0458_ 0.0013f
C26545 _0458_ acc0.A\[15\] 0.01097f
C26546 _0820_/a_297_297# _0820_/a_215_47# 0
C26547 _0820_/a_79_21# _0820_/a_510_47# 0.00844f
C26548 net103 net43 0
C26549 net165 _0158_ 0
C26550 hold28/a_391_47# _1049_/a_1059_315# 0.01554f
C26551 _0343_ _0642_/a_215_297# 0.00443f
C26552 hold64/a_285_47# _0350_ 0.00618f
C26553 net53 _0359_ 0.21641f
C26554 _1058_/a_27_47# clknet_1_1__leaf__0465_ 0.04336f
C26555 _0181_ _0393_ 0
C26556 acc0.A\[3\] _0262_ 0
C26557 _1038_/a_1059_315# net174 0
C26558 _1059_/a_975_413# _0369_ 0
C26559 _0182_ _1048_/a_27_47# 0.00459f
C26560 _0799_/a_209_297# _0297_ 0
C26561 _1001_/a_193_47# net46 0.00174f
C26562 pp[26] hold8/a_285_47# 0
C26563 _1041_/a_466_413# _0550_/a_51_297# 0
C26564 _1035_/a_592_47# _0175_ 0.00112f
C26565 _0292_ net47 0
C26566 _0222_ _0762_/a_79_21# 0.00452f
C26567 _0284_ net38 0.15248f
C26568 _0285_ acc0.A\[11\] 0.18195f
C26569 _0343_ net51 0.3569f
C26570 _0266_ _0634_/a_113_47# 0.00937f
C26571 _0248_ _0104_ 0
C26572 B[15] _0175_ 0
C26573 net69 _0853_/a_150_297# 0
C26574 net67 acc0.A\[9\] 0.32994f
C26575 net36 hold2/a_285_47# 0
C26576 net40 output39/a_27_47# 0
C26577 _0146_ net170 0
C26578 clknet_1_0__leaf__0463_ _1046_/a_975_413# 0
C26579 _0957_/a_32_297# control0.sh 0
C26580 _0811_/a_299_297# _0345_ 0.00379f
C26581 _0837_/a_266_47# _1051_/a_27_47# 0
C26582 _1039_/a_27_47# _0913_/a_27_47# 0
C26583 _0399_ _0394_ 0
C26584 clknet_0__0464_ net9 0
C26585 net44 _0705_/a_59_75# 0
C26586 acc0.A\[12\] net3 0
C26587 control0.state\[0\] _0165_ 0
C26588 _0570_/a_27_297# _0687_/a_59_75# 0
C26589 _1035_/a_1017_47# control0.sh 0.00115f
C26590 _0172_ _0527_/a_27_297# 0
C26591 _1000_/a_466_413# _0393_ 0.00279f
C26592 _0107_ net52 0
C26593 net23 control0.sh 0.02732f
C26594 _0413_ _0799_/a_80_21# 0.07799f
C26595 clkbuf_1_0__f__0459_/a_110_47# _0459_ 0.02713f
C26596 _0985_/a_1059_315# _0446_ 0
C26597 _0680_/a_217_297# _0238_ 0.00262f
C26598 comp0.B\[12\] _1044_/a_634_159# 0
C26599 _0449_ clkbuf_0__0458_/a_110_47# 0.00148f
C26600 _0456_ _0261_ 0
C26601 _1066_/a_193_47# net17 0
C26602 _0534_/a_81_21# clkbuf_1_1__f__0457_/a_110_47# 0
C26603 net207 _0580_/a_109_297# 0
C26604 clknet_1_1__leaf__0460_ _0690_/a_68_297# 0.00215f
C26605 _0254_ _0622_/a_193_47# 0.01172f
C26606 _0967_/a_109_93# control0.state\[2\] 0
C26607 net143 acc0.A\[10\] 0.08989f
C26608 control0.count\[1\] _1069_/a_1017_47# 0.002f
C26609 _0168_ clknet_1_0__leaf_clk 0.43158f
C26610 _0486_ _0485_ 0
C26611 control0.state\[2\] _0487_ 0.79527f
C26612 hold39/a_391_47# clknet_1_1__leaf__0463_ 0.03228f
C26613 hold79/a_285_47# _0478_ 0
C26614 pp[25] _0123_ 0
C26615 net53 net200 0.08904f
C26616 hold75/a_285_47# _0346_ 0
C26617 _1018_/a_381_47# _0218_ 0
C26618 _1030_/a_891_413# _0336_ 0.01837f
C26619 _0414_ _0994_/a_634_159# 0
C26620 _0369_ _1005_/a_891_413# 0
C26621 _1017_/a_466_413# clknet_1_1__leaf__0461_ 0
C26622 _0083_ _0186_ 0.01464f
C26623 _1000_/a_381_47# _0245_ 0.01487f
C26624 _1000_/a_1059_315# _0246_ 0
C26625 acc0.A\[14\] _0507_/a_27_297# 0.00625f
C26626 _0216_ _1006_/a_634_159# 0.01148f
C26627 _1006_/a_1059_315# net92 0
C26628 _0322_ _0345_ 0
C26629 VPWR _0974_/a_79_199# 0.31887f
C26630 _0179_ _0458_ 0.04419f
C26631 init B[3] 0.1196f
C26632 _0839_/a_109_297# _0841_/a_79_21# 0
C26633 _0570_/a_109_297# hold9/a_285_47# 0
C26634 _0570_/a_27_297# hold9/a_391_47# 0.01653f
C26635 hold10/a_285_47# _0137_ 0
C26636 net59 _0340_ 0
C26637 output59/a_27_47# _0342_ 0
C26638 _0327_ _0345_ 0
C26639 _0984_/a_1059_315# _0984_/a_1017_47# 0
C26640 _0984_/a_193_47# net70 0.00474f
C26641 _0201_ net196 0
C26642 _0172_ _1061_/a_27_47# 0.04542f
C26643 _0583_/a_27_297# net219 0
C26644 _0312_ _0219_ 0.11448f
C26645 _0643_/a_103_199# _0269_ 0.13581f
C26646 _0200_ hold6/a_285_47# 0
C26647 _0984_/a_27_47# _0506_/a_81_21# 0
C26648 acc0.A\[14\] net165 0
C26649 _0808_/a_266_47# _0091_ 0
C26650 clkload3/Y _1017_/a_193_47# 0
C26651 _0424_ _0347_ 0
C26652 acc0.A\[17\] _0218_ 0.54037f
C26653 A[4] net12 0.00212f
C26654 net178 net76 0
C26655 acc0.A\[19\] _0391_ 0.01953f
C26656 _0765_/a_297_297# _0369_ 0.00382f
C26657 net58 pp[4] 0.00832f
C26658 clknet_1_0__leaf__0465_ input15/a_75_212# 0
C26659 _0568_/a_27_297# net116 0
C26660 net213 _0352_ 0.00115f
C26661 VPWR _0988_/a_634_159# 0.17885f
C26662 _0514_/a_109_47# acc0.A\[10\] 0.00173f
C26663 _0474_ hold84/a_391_47# 0
C26664 acc0.A\[29\] _0703_/a_109_297# 0
C26665 _1015_/a_193_47# clknet_1_0__leaf__0457_ 0.00115f
C26666 _0529_/a_27_297# _0447_ 0
C26667 _0285_ hold81/a_391_47# 0
C26668 _1059_/a_193_47# _0184_ 0
C26669 hold78/a_285_47# _1031_/a_891_413# 0
C26670 _0344_ _1031_/a_193_47# 0
C26671 hold78/a_391_47# _1031_/a_1059_315# 0
C26672 net168 _1054_/a_1059_315# 0
C26673 hold6/a_49_47# _0206_ 0
C26674 VPWR _0953_/a_114_297# 0.00681f
C26675 net12 _0085_ 0
C26676 _1056_/a_466_413# _0186_ 0
C26677 clknet_1_1__leaf_clk net107 0.01475f
C26678 output59/a_27_47# _0334_ 0
C26679 _1023_/a_466_413# acc0.A\[23\] 0
C26680 hold43/a_285_47# _0127_ 0.00287f
C26681 _1023_/a_381_47# net177 0.1369f
C26682 _0277_ _0301_ 0.02014f
C26683 _0581_/a_27_297# acc0.A\[19\] 0
C26684 _0512_/a_373_47# acc0.A\[10\] 0
C26685 _0369_ _1006_/a_466_413# 0.00304f
C26686 _0465_ _0840_/a_68_297# 0.00619f
C26687 _1044_/a_27_47# net20 0.02684f
C26688 _0259_ VPWR 1.28278f
C26689 net23 net157 0
C26690 acc0.A\[27\] net97 0
C26691 _0216_ _0571_/a_109_297# 0.0505f
C26692 net155 _0571_/a_109_47# 0.00243f
C26693 _0538_/a_512_297# _0172_ 0.00116f
C26694 _0699_/a_68_297# _0318_ 0
C26695 net60 _0218_ 0
C26696 _0337_ hold62/a_285_47# 0
C26697 _0757_/a_150_297# _0378_ 0
C26698 _0380_ _0756_/a_47_47# 0.00103f
C26699 _0263_ _0842_/a_145_75# 0
C26700 net161 comp0.B\[4\] 0.00211f
C26701 _0218_ net5 0.17148f
C26702 _0724_/a_113_297# _0334_ 0.03025f
C26703 clkbuf_1_0__f__0463_/a_110_47# _0548_/a_149_47# 0
C26704 _1001_/a_634_159# VPWR 0.18383f
C26705 net45 _1017_/a_27_47# 0.01415f
C26706 net120 net119 0.24205f
C26707 net163 _1031_/a_1059_315# 0
C26708 _0477_ _0163_ 0
C26709 net70 net145 0.00329f
C26710 VPWR _1062_/a_193_47# 0.29086f
C26711 _0616_/a_292_297# _0247_ 0.00476f
C26712 _1059_/a_381_47# net229 0.02216f
C26713 _0091_ _0345_ 0.00214f
C26714 _1039_/a_27_47# _0172_ 0.01058f
C26715 VPWR hold90/a_49_47# 0.26466f
C26716 _0376_ net51 0.04173f
C26717 _1038_/a_891_413# _1037_/a_891_413# 0
C26718 net43 output41/a_27_47# 0
C26719 _0499_/a_59_75# net201 0
C26720 _0537_/a_68_297# _0473_ 0
C26721 VPWR hold8/a_391_47# 0.19167f
C26722 net167 _0488_ 0.02573f
C26723 _0762_/a_79_21# _0762_/a_297_297# 0.01735f
C26724 _0490_ _0466_ 0.08237f
C26725 _0997_/a_381_47# _0095_ 0.1145f
C26726 hold20/a_285_47# _1068_/a_1059_315# 0.00334f
C26727 _0677_/a_377_297# _0393_ 0
C26728 _0574_/a_27_297# acc0.A\[24\] 0.02206f
C26729 _0456_ net47 0
C26730 net54 clknet_0__0462_ 0
C26731 net193 hold6/a_285_47# 0
C26732 pp[8] clknet_1_1__leaf__0465_ 0.03562f
C26733 comp0.B\[4\] net26 0.35673f
C26734 net212 _0619_/a_68_297# 0
C26735 _1053_/a_466_413# hold83/a_49_47# 0
C26736 _0406_ net41 0.02761f
C26737 _0389_ clknet_1_0__leaf__0457_ 0
C26738 _1065_/a_634_159# _1065_/a_1059_315# 0
C26739 _1065_/a_27_47# _1065_/a_381_47# 0.05761f
C26740 _1065_/a_193_47# _1065_/a_891_413# 0.19226f
C26741 VPWR _0561_/a_245_297# 0.00545f
C26742 net140 net11 0.10518f
C26743 control0.count\[2\] _0489_ 0
C26744 net232 _1066_/a_891_413# 0
C26745 _0998_/a_634_159# _0218_ 0
C26746 _1036_/a_1059_315# _1035_/a_27_47# 0
C26747 _1036_/a_466_413# _1035_/a_193_47# 0.00112f
C26748 _0532_/a_81_21# _0146_ 0.11484f
C26749 net31 _0548_/a_51_297# 0.1178f
C26750 _0707_/a_201_297# _0707_/a_544_297# 0.00702f
C26751 _0707_/a_75_199# _0707_/a_208_47# 0.0159f
C26752 _1033_/a_1059_315# _0565_/a_240_47# 0
C26753 _1033_/a_891_413# _0565_/a_149_47# 0
C26754 _0209_ net27 0
C26755 hold79/a_285_47# _1070_/a_193_47# 0
C26756 hold79/a_49_47# _1070_/a_634_159# 0
C26757 _0954_/a_32_297# _1042_/a_1059_315# 0
C26758 _0954_/a_304_297# _1042_/a_193_47# 0
C26759 _1014_/a_27_47# _1014_/a_634_159# 0.14145f
C26760 _0311_ _0352_ 0.00265f
C26761 VPWR _1047_/a_466_413# 0.25465f
C26762 _0627_/a_297_297# clknet_0__0465_ 0
C26763 _0238_ _0372_ 0.62817f
C26764 _0181_ net206 0
C26765 clknet_0__0463_ comp0.B\[1\] 0
C26766 clknet_1_0__leaf__0464_ acc0.A\[3\] 0.00246f
C26767 _0995_/a_27_47# _0411_ 0
C26768 _0457_ _0566_/a_27_47# 0
C26769 VPWR net221 1.66438f
C26770 _0483_ net35 0
C26771 VPWR _1007_/a_381_47# 0.0794f
C26772 _0399_ _0989_/a_891_413# 0
C26773 _0996_/a_193_47# _0459_ 0
C26774 net180 _1040_/a_1017_47# 0
C26775 _1058_/a_975_413# VPWR 0.00464f
C26776 _0179_ _1051_/a_891_413# 0.00444f
C26777 net236 _0490_ 0
C26778 hold34/a_49_47# A[11] 0
C26779 _0080_ _0181_ 0.15583f
C26780 clknet_0__0465_ _0817_/a_266_47# 0
C26781 _0312_ _0746_/a_81_21# 0.01053f
C26782 net61 hold65/a_285_47# 0.03289f
C26783 _0734_/a_47_47# VPWR 0.40869f
C26784 hold49/a_49_47# _0537_/a_68_297# 0.00216f
C26785 _0171_ _0173_ 0.24903f
C26786 _0298_ _0301_ 0
C26787 _0278_ acc0.A\[13\] 0.08942f
C26788 _0558_/a_150_297# VPWR 0.00166f
C26789 _1055_/a_27_47# _0190_ 0.00422f
C26790 _1055_/a_634_159# net16 0.00638f
C26791 clknet_1_1__leaf__0465_ _1060_/a_27_47# 0.00241f
C26792 _1064_/a_891_413# _1064_/a_1017_47# 0.00617f
C26793 hold78/a_49_47# _0219_ 0
C26794 _0728_/a_145_75# _0219_ 0
C26795 net169 hold7/a_285_47# 0
C26796 _1018_/a_193_47# net103 0
C26797 _1000_/a_27_47# _0116_ 0
C26798 hold41/a_285_47# A[11] 0
C26799 _0837_/a_266_47# _0085_ 0
C26800 net112 _1025_/a_634_159# 0
C26801 _0296_ _0301_ 0.12554f
C26802 _0712_/a_297_297# _0344_ 0.00116f
C26803 _1002_/a_193_47# _1067_/a_891_413# 0
C26804 _0326_ acc0.A\[24\] 0
C26805 comp0.B\[14\] _0140_ 0
C26806 _0389_ _1001_/a_1059_315# 0
C26807 net1 _0161_ 0.21529f
C26808 _0959_/a_300_47# clknet_1_1__leaf_clk 0
C26809 _0728_/a_59_75# _0728_/a_145_75# 0.00658f
C26810 _0149_ net148 0
C26811 _0343_ _1017_/a_592_47# 0
C26812 net230 hold83/a_391_47# 0.13412f
C26813 _0151_ hold83/a_49_47# 0.0012f
C26814 _1025_/a_634_159# acc0.A\[24\] 0
C26815 clkbuf_0__0461_/a_110_47# _0459_ 0.01979f
C26816 _0131_ comp0.B\[0\] 0.00255f
C26817 clknet_1_0__leaf__0462_ _0753_/a_381_47# 0
C26818 _0257_ _0624_/a_145_75# 0
C26819 _0230_ _0374_ 0.04301f
C26820 _0363_ _0318_ 0.00338f
C26821 _0985_/a_1059_315# net61 0.13106f
C26822 _1013_/a_1059_315# _0339_ 0.00206f
C26823 _0349_ _0356_ 0
C26824 _0981_/a_27_297# _0981_/a_109_297# 0.17136f
C26825 _0804_/a_79_21# _0647_/a_285_47# 0
C26826 acc0.A\[12\] _0644_/a_47_47# 0
C26827 _0285_ _0281_ 0.31995f
C26828 _1017_/a_975_413# acc0.A\[17\] 0
C26829 _0195_ _0704_/a_68_297# 0
C26830 _0603_/a_68_297# _0352_ 0.00202f
C26831 net114 net156 0
C26832 hold24/a_391_47# clkbuf_1_0__f__0463_/a_110_47# 0.01292f
C26833 A[4] pp[5] 0
C26834 _0136_ _0209_ 0.12994f
C26835 _0352_ hold73/a_391_47# 0
C26836 pp[27] _0195_ 0.12618f
C26837 VPWR _0782_/a_27_47# 0.4512f
C26838 hold13/a_391_47# comp0.B\[2\] 0
C26839 _0129_ _0219_ 0
C26840 _0222_ _1022_/a_634_159# 0.01041f
C26841 _0855_/a_299_297# net149 0.05915f
C26842 _0481_ _1070_/a_27_47# 0
C26843 _0854_/a_510_47# _0455_ 0.00404f
C26844 _1037_/a_193_47# _1036_/a_27_47# 0
C26845 _1037_/a_27_47# _1036_/a_193_47# 0
C26846 _0313_ _1026_/a_466_413# 0
C26847 acc0.A\[12\] _0401_ 0
C26848 hold21/a_285_47# net12 0
C26849 _0600_/a_103_199# _0366_ 0
C26850 _0817_/a_81_21# _0423_ 0.03177f
C26851 _0346_ _0808_/a_266_47# 0.00415f
C26852 _0999_/a_193_47# _0352_ 0.02253f
C26853 _0224_ net51 0.02099f
C26854 _0255_ net154 0
C26855 hold28/a_391_47# net175 0.16343f
C26856 _0477_ _1066_/a_27_47# 0
C26857 _0498_/a_245_297# _0498_/a_240_47# 0
C26858 _0830_/a_215_47# _0087_ 0.00324f
C26859 _0841_/a_215_47# _0986_/a_27_47# 0
C26860 clknet_1_1__leaf__0460_ _1028_/a_634_159# 0
C26861 _0640_/a_215_297# _0255_ 0.16533f
C26862 _0313_ hold97/a_391_47# 0
C26863 _1015_/a_381_47# clknet_1_0__leaf__0461_ 0
C26864 clknet_1_0__leaf__0464_ net157 0.00181f
C26865 clknet_1_0__leaf__0465_ _1052_/a_1017_47# 0
C26866 _0272_ clknet_0__0465_ 0.0044f
C26867 net36 _1040_/a_193_47# 0
C26868 clknet_1_1__leaf__0459_ input5/a_75_212# 0
C26869 _0195_ _0198_ 0.04676f
C26870 _0557_/a_149_47# _0557_/a_240_47# 0.06872f
C26871 net138 net139 0.00171f
C26872 net173 net10 0
C26873 _0183_ net166 0.00108f
C26874 _0514_/a_373_47# _0181_ 0.00122f
C26875 _0216_ _1014_/a_27_47# 0
C26876 _0195_ _1014_/a_634_159# 0
C26877 output56/a_27_47# net59 0
C26878 _0684_/a_59_75# clknet_0__0460_ 0.06097f
C26879 hold11/a_391_47# net10 0
C26880 _0292_ _0294_ 0.00173f
C26881 comp0.B\[12\] _0176_ 0.10412f
C26882 _0682_/a_68_297# _0352_ 0
C26883 _0330_ _0727_/a_109_47# 0
C26884 _0329_ _0221_ 0
C26885 _0341_ net99 0
C26886 _0856_/a_79_21# _1014_/a_891_413# 0
C26887 _0439_ _0253_ 0
C26888 _1001_/a_27_47# net87 0.22161f
C26889 _0305_ net78 0
C26890 acc0.A\[27\] _1010_/a_27_47# 0
C26891 _0255_ _0465_ 0.01686f
C26892 _0260_ clkbuf_0__0458_/a_110_47# 0.08515f
C26893 _1018_/a_27_47# net206 0.02616f
C26894 VPWR _0253_ 0.61564f
C26895 _0158_ _0185_ 0.01758f
C26896 _0356_ _0701_/a_209_297# 0
C26897 _0707_/a_75_199# acc0.A\[30\] 0
C26898 _1008_/a_634_159# _1008_/a_466_413# 0.23992f
C26899 _1008_/a_193_47# _1008_/a_1059_315# 0.03405f
C26900 _1008_/a_27_47# _1008_/a_891_413# 0.03224f
C26901 _0423_ _0084_ 0
C26902 acc0.A\[20\] _0902_/a_27_47# 0.00194f
C26903 _0976_/a_439_47# clknet_1_0__leaf_clk 0
C26904 _0976_/a_505_21# control0.count\[0\] 0.24407f
C26905 hold16/a_391_47# net163 0.13094f
C26906 clknet_1_0__leaf__0463_ B[7] 0.02412f
C26907 output43/a_27_47# _0995_/a_193_47# 0
C26908 hold76/a_391_47# net211 0
C26909 _1020_/a_634_159# _1020_/a_1017_47# 0
C26910 _1020_/a_466_413# _1020_/a_592_47# 0.00553f
C26911 _0343_ _0324_ 0
C26912 _0408_ acc0.A\[15\] 0
C26913 _0250_ _0758_/a_215_47# 0
C26914 _1035_/a_1059_315# comp0.B\[3\] 0.08411f
C26915 _0195_ net83 0.03287f
C26916 net156 _0365_ 0
C26917 net23 _0955_/a_32_297# 0
C26918 _0230_ _0752_/a_300_297# 0
C26919 _0598_/a_79_21# _0376_ 0
C26920 _0770_/a_79_21# _0218_ 0
C26921 hold28/a_49_47# acc0.A\[3\] 0.04604f
C26922 _0983_/a_1017_47# net47 0
C26923 _0502_/a_27_47# control0.reset 0
C26924 hold85/a_49_47# VPWR 0.27906f
C26925 _0346_ _0345_ 1.77227f
C26926 _0746_/a_299_297# _0219_ 0
C26927 acc0.A\[27\] _1009_/a_193_47# 0
C26928 _0346_ _0814_/a_27_47# 0
C26929 clknet_0__0458_ _0986_/a_193_47# 0.00575f
C26930 _0195_ _0781_/a_68_297# 0
C26931 clknet_0__0457_ _1014_/a_193_47# 0.00562f
C26932 hold34/a_49_47# net66 0
C26933 control0.sh _0213_ 0
C26934 _0471_ _1065_/a_27_47# 0
C26935 net216 _0249_ 0
C26936 _0180_ _1048_/a_1017_47# 0
C26937 _1031_/a_891_413# hold61/a_391_47# 0
C26938 _0188_ _0512_/a_373_47# 0
C26939 _1054_/a_27_47# _0518_/a_27_297# 0.00144f
C26940 _1013_/a_891_413# net99 0
C26941 hold14/a_285_47# VPWR 0.29492f
C26942 _0314_ _0367_ 0.01624f
C26943 _0313_ _0315_ 0.42328f
C26944 _1041_/a_466_413# _0172_ 0.01427f
C26945 _1041_/a_891_413# net180 0
C26946 _1041_/a_193_47# _0137_ 0
C26947 clknet_1_1__leaf__0459_ pp[12] 0
C26948 _0266_ _0635_/a_27_47# 0.00471f
C26949 VPWR input27/a_75_212# 0.2142f
C26950 _0559_/a_512_297# _0133_ 0
C26951 pp[28] net57 0.06308f
C26952 _0988_/a_27_47# acc0.A\[6\] 0
C26953 _0992_/a_466_413# _0345_ 0
C26954 _0109_ hold80/a_285_47# 0
C26955 net166 acc0.A\[15\] 0
C26956 _0226_ clkbuf_1_0__f__0460_/a_110_47# 0
C26957 clkbuf_1_1__f__0457_/a_110_47# hold71/a_391_47# 0.00131f
C26958 hold94/a_49_47# _0345_ 0.00282f
C26959 hold21/a_49_47# A[8] 0.01398f
C26960 _0570_/a_27_297# _0352_ 0.00147f
C26961 _0991_/a_634_159# acc0.A\[15\] 0
C26962 _0441_ _1051_/a_891_413# 0
C26963 _0984_/a_27_47# _0184_ 0
C26964 clknet_0__0459_ _0796_/a_215_47# 0
C26965 _0346_ hold2/a_49_47# 0.00224f
C26966 hold63/a_391_47# net53 0
C26967 clknet_1_0__leaf__0459_ net221 0.02013f
C26968 _0982_/a_1059_315# _0855_/a_81_21# 0.00146f
C26969 net185 _0175_ 0.08764f
C26970 _0953_/a_32_297# _0913_/a_27_47# 0.01241f
C26971 _1010_/a_27_47# _0110_ 0
C26972 _0230_ _0249_ 0
C26973 hold42/a_391_47# _1058_/a_193_47# 0.00224f
C26974 net26 _0549_/a_150_297# 0
C26975 _0098_ _0393_ 0.03266f
C26976 VPWR _0535_/a_150_297# 0.00127f
C26977 _0578_/a_109_297# net150 0.01656f
C26978 _0578_/a_27_297# _0217_ 0.16909f
C26979 _1058_/a_891_413# _1057_/a_193_47# 0.00115f
C26980 _1058_/a_466_413# _1057_/a_466_413# 0.00177f
C26981 _1058_/a_193_47# _1057_/a_891_413# 0.00115f
C26982 clknet_1_1__leaf__0460_ _0371_ 0.1633f
C26983 _0788_/a_68_297# net80 0
C26984 comp0.B\[12\] net130 0
C26985 _0795_/a_81_21# hold91/a_49_47# 0
C26986 net168 hold22/a_285_47# 0.0464f
C26987 B[12] net196 0
C26988 _0576_/a_109_297# clknet_1_0__leaf__0460_ 0
C26989 _0236_ _0374_ 0.01426f
C26990 _1000_/a_891_413# _0352_ 0.03168f
C26991 _0212_ control0.sh 0.02794f
C26992 VPWR _1063_/a_975_413# 0.00418f
C26993 _0088_ _0186_ 0
C26994 _0284_ _0654_/a_297_47# 0.00124f
C26995 net213 _0237_ 0.03638f
C26996 _0383_ _0103_ 0
C26997 net45 _0245_ 0.12445f
C26998 _0195_ _0216_ 1.54561f
C26999 hold36/a_391_47# _0473_ 0
C27000 acc0.A\[14\] _0185_ 0.37412f
C27001 hold13/a_49_47# VPWR 0.27255f
C27002 VPWR _0585_/a_373_47# 0
C27003 _1014_/a_27_47# net247 0
C27004 _0216_ net92 0.00188f
C27005 _0580_/a_27_297# _0264_ 0
C27006 _0328_ _0462_ 0.04505f
C27007 VPWR _1017_/a_27_47# 0.4266f
C27008 acc0.A\[26\] _0365_ 0.00369f
C27009 _0126_ hold9/a_391_47# 0.05249f
C27010 _0267_ _0842_/a_59_75# 0.19941f
C27011 _0432_ _0444_ 0.05156f
C27012 _0443_ _0445_ 0.09431f
C27013 net219 _0615_/a_109_297# 0.00303f
C27014 net180 net147 0
C27015 net55 clkbuf_1_1__f__0462_/a_110_47# 0.0023f
C27016 _0548_/a_51_297# _0548_/a_240_47# 0.03076f
C27017 VPWR _1060_/a_975_413# 0.00489f
C27018 _1015_/a_27_47# net149 0
C27019 clkload1/a_268_47# _0346_ 0.00205f
C27020 _1043_/a_27_47# net153 0
C27021 _1056_/a_193_47# A[10] 0
C27022 hold65/a_391_47# clkbuf_1_0__f__0465_/a_110_47# 0.00138f
C27023 _0179_ _0291_ 0
C27024 hold36/a_391_47# clkbuf_1_1__f__0464_/a_110_47# 0
C27025 clknet_0_clk _1063_/a_193_47# 0
C27026 VPWR net74 0.53379f
C27027 net17 clkbuf_1_1__f_clk/a_110_47# 0.01886f
C27028 _0157_ net6 0
C27029 _0713_/a_27_47# clknet_1_0__leaf__0457_ 0
C27030 clknet_1_0__leaf__0459_ _0782_/a_27_47# 0
C27031 VPWR _1050_/a_193_47# 0.30603f
C27032 _0511_/a_299_297# _0511_/a_384_47# 0
C27033 net157 _1047_/a_592_47# 0.00315f
C27034 _0452_ _0850_/a_150_297# 0
C27035 _0305_ _0387_ 0.4562f
C27036 hold21/a_285_47# pp[5] 0
C27037 net177 acc0.A\[23\] 0
C27038 acc0.A\[14\] _0998_/a_1059_315# 0
C27039 clknet_0_clk _0460_ 0
C27040 acc0.A\[7\] _0619_/a_150_297# 0
C27041 comp0.B\[15\] _0181_ 0.00463f
C27042 hold45/a_49_47# net192 0.00157f
C27043 acc0.A\[8\] net75 0.1347f
C27044 _1010_/a_27_47# _1010_/a_193_47# 0.96639f
C27045 _0179_ _0991_/a_634_159# 0
C27046 _1016_/a_1017_47# _0181_ 0
C27047 _0116_ acc0.A\[19\] 0
C27048 _0644_/a_47_47# net42 0.37179f
C27049 _0348_ _1011_/a_1059_315# 0
C27050 _0670_/a_79_21# _0302_ 0.05038f
C27051 pp[27] _1010_/a_891_413# 0
C27052 _0183_ acc0.A\[1\] 0.02175f
C27053 _0217_ _0180_ 0
C27054 pp[30] _0110_ 0
C27055 clkbuf_0__0462_/a_110_47# clkbuf_1_0__f__0462_/a_110_47# 0.00301f
C27056 _0299_ _0411_ 0.05403f
C27057 VPWR output61/a_27_47# 0.40665f
C27058 _0457_ _1015_/a_1017_47# 0
C27059 _0319_ _0350_ 0
C27060 _0198_ _1048_/a_193_47# 0
C27061 _0143_ _0172_ 0.0219f
C27062 net36 _0853_/a_68_297# 0.00147f
C27063 _0536_/a_245_297# net157 0.00106f
C27064 VPWR _0973_/a_27_297# 0.23896f
C27065 hold96/a_49_47# _0216_ 0.05534f
C27066 _0218_ _0281_ 0.01242f
C27067 _1033_/a_1059_315# _0171_ 0
C27068 _0195_ _0852_/a_285_297# 0
C27069 _0236_ acc0.A\[19\] 0
C27070 _1002_/a_27_47# net150 0
C27071 _0746_/a_81_21# _0746_/a_299_297# 0.08213f
C27072 _0276_ _0409_ 0
C27073 hold18/a_391_47# net247 0.0134f
C27074 hold88/a_49_47# _0990_/a_27_47# 0
C27075 VPWR _0772_/a_215_47# 0
C27076 _0749_/a_81_21# _1006_/a_193_47# 0
C27077 _1020_/a_634_159# _0461_ 0.00207f
C27078 _0397_ _0347_ 0.43421f
C27079 _1018_/a_891_413# _0347_ 0.01069f
C27080 net78 _0181_ 0
C27081 _0174_ _0550_/a_51_297# 0.10216f
C27082 _0578_/a_109_297# control0.add 0.05291f
C27083 clknet_0__0465_ _0181_ 0.26504f
C27084 _1021_/a_1017_47# VPWR 0
C27085 _0369_ _0240_ 0.04873f
C27086 _0172_ _0953_/a_32_297# 0.00256f
C27087 acc0.A\[12\] hold70/a_49_47# 0
C27088 _0231_ _0758_/a_510_47# 0
C27089 _0343_ _0347_ 1.22317f
C27090 _1000_/a_466_413# _0773_/a_35_297# 0
C27091 _1009_/a_27_47# _1009_/a_466_413# 0.27314f
C27092 _1009_/a_193_47# _1009_/a_634_159# 0.12482f
C27093 _0306_ _0394_ 0.21109f
C27094 _0698_/a_113_297# acc0.A\[28\] 0
C27095 VPWR _0518_/a_109_297# 0.17811f
C27096 net36 _1061_/a_1059_315# 0
C27097 _0576_/a_27_297# _0576_/a_109_47# 0.00393f
C27098 _0645_/a_47_47# _1059_/a_27_47# 0
C27099 _0195_ net247 0.05325f
C27100 _1065_/a_27_47# control0.reset 0.00454f
C27101 _0677_/a_285_47# _0352_ 0
C27102 net36 _0207_ 0.04053f
C27103 _0982_/a_27_47# VPWR 0.67147f
C27104 clknet_0_clk _1062_/a_891_413# 0.02202f
C27105 net228 net5 0
C27106 _0967_/a_215_297# _1066_/a_381_47# 0
C27107 net213 _1005_/a_27_47# 0
C27108 _0424_ _0991_/a_1059_315# 0
C27109 net84 _0218_ 0.03145f
C27110 _1036_/a_634_159# net121 0.01565f
C27111 _1036_/a_193_47# _0133_ 0.00655f
C27112 _0343_ _0104_ 0
C27113 _0346_ net52 0.35061f
C27114 _0180_ _0142_ 0.03681f
C27115 _0186_ _0522_/a_373_47# 0.00182f
C27116 net111 _1025_/a_634_159# 0
C27117 net7 _0548_/a_51_297# 0.10126f
C27118 net202 control0.add 0
C27119 net14 acc0.A\[6\] 0
C27120 net168 net13 0.00458f
C27121 _1036_/a_381_47# B[15] 0
C27122 _0236_ _0249_ 0
C27123 _0967_/a_215_297# net1 0.10701f
C27124 _0166_ _0970_/a_27_297# 0
C27125 _0819_/a_81_21# _0346_ 0.17697f
C27126 _0992_/a_891_413# _0811_/a_299_297# 0
C27127 _0856_/a_510_47# net247 0
C27128 _0707_/a_544_297# _0339_ 0
C27129 _0218_ _0842_/a_145_75# 0.00125f
C27130 acc0.A\[1\] acc0.A\[15\] 0.34814f
C27131 comp0.B\[1\] _0565_/a_512_297# 0.00169f
C27132 _0243_ _0241_ 0.05649f
C27133 hold79/a_285_47# VPWR 0.31097f
C27134 comp0.B\[11\] _1042_/a_592_47# 0.00188f
C27135 _1014_/a_891_413# _1014_/a_975_413# 0.00851f
C27136 _1014_/a_27_47# net100 0.44062f
C27137 _1014_/a_381_47# _1014_/a_561_413# 0.00123f
C27138 _0643_/a_103_199# clkbuf_0__0458_/a_110_47# 0
C27139 _1071_/a_193_47# _1071_/a_381_47# 0.09972f
C27140 _1071_/a_634_159# _1071_/a_891_413# 0.03684f
C27141 _1071_/a_27_47# _1071_/a_561_413# 0.0027f
C27142 net152 _0142_ 0
C27143 VPWR _0145_ 0.33582f
C27144 net48 _0973_/a_27_297# 0
C27145 _1015_/a_1059_315# _0208_ 0.067f
C27146 _0333_ hold62/a_285_47# 0
C27147 VPWR pp[23] 0.1845f
C27148 B[13] input19/a_75_212# 0.00313f
C27149 input21/a_75_212# B[11] 0.04738f
C27150 hold96/a_49_47# hold96/a_391_47# 0.00188f
C27151 clknet_0__0463_ _0496_/a_27_47# 0
C27152 _0985_/a_975_413# _0458_ 0
C27153 net54 _0687_/a_59_75# 0.17945f
C27154 _1013_/a_27_47# net42 0
C27155 _0852_/a_35_297# _0852_/a_285_297# 0.02504f
C27156 _0717_/a_80_21# pp[29] 0
C27157 pp[0] B[1] 0
C27158 _0179_ _0290_ 0.38686f
C27159 _1050_/a_381_47# net9 0.00433f
C27160 _0983_/a_27_47# acc0.A\[14\] 0
C27161 _0343_ _0792_/a_209_297# 0.01241f
C27162 _0231_ _0230_ 0.26444f
C27163 _0458_ _1049_/a_891_413# 0
C27164 _0183_ _0388_ 0
C27165 hold39/a_49_47# hold39/a_285_47# 0.22264f
C27166 _1035_/a_193_47# net26 0.02379f
C27167 VPWR net17 1.12243f
C27168 _0815_/a_199_47# _0181_ 0.00128f
C27169 _0836_/a_68_297# net65 0
C27170 _0280_ _0806_/a_113_297# 0
C27171 _0178_ _0147_ 0
C27172 VPWR net238 0.39035f
C27173 _0670_/a_79_21# net6 0.12166f
C27174 net141 net16 0
C27175 _0216_ net90 0.03425f
C27176 net65 net212 0.32538f
C27177 _0087_ _0989_/a_27_47# 0.09207f
C27178 net212 _0989_/a_466_413# 0
C27179 _0437_ _0989_/a_634_159# 0.00356f
C27180 _0179_ _0528_/a_81_21# 0.0074f
C27181 hold98/a_49_47# pp[14] 0.03072f
C27182 net40 output41/a_27_47# 0.00586f
C27183 hold98/a_391_47# net41 0
C27184 _0346_ _0791_/a_113_297# 0
C27185 VPWR _0446_ 1.82396f
C27186 _1015_/a_466_413# net17 0
C27187 VPWR input2/a_75_212# 0.22544f
C27188 _0081_ _0852_/a_285_297# 0
C27189 _1026_/a_592_47# acc0.A\[25\] 0.00121f
C27190 _0295_ _0809_/a_299_297# 0.0989f
C27191 net36 _1039_/a_1059_315# 0.08648f
C27192 A[11] net4 0.0257f
C27193 _0195_ _1048_/a_466_413# 0
C27194 _0390_ _0772_/a_215_47# 0
C27195 _1002_/a_27_47# control0.add 0
C27196 net88 _1067_/a_1059_315# 0.00176f
C27197 _1012_/a_466_413# _0352_ 0.01197f
C27198 _1012_/a_381_47# _0347_ 0.00913f
C27199 net54 hold9/a_391_47# 0.01999f
C27200 _0819_/a_384_47# _0427_ 0
C27201 _0819_/a_299_297# _0428_ 0.04426f
C27202 clknet_1_0__leaf__0460_ hold94/a_285_47# 0.00181f
C27203 acc0.A\[25\] net110 0
C27204 _0343_ _1016_/a_891_413# 0.0046f
C27205 _1033_/a_27_47# _0215_ 0.00602f
C27206 net194 VPWR 0.6136f
C27207 output40/a_27_47# pp[13] 0.16123f
C27208 net180 _0473_ 0.00539f
C27209 clknet_1_0__leaf__0459_ _1017_/a_27_47# 0.02637f
C27210 net193 _0537_/a_68_297# 0
C27211 _0216_ _1010_/a_891_413# 0
C27212 acc0.A\[31\] _0341_ 0.33917f
C27213 _0981_/a_109_297# _0170_ 0.00469f
C27214 net48 pp[23] 0
C27215 pp[20] net51 0
C27216 _1052_/a_891_413# _0180_ 0.00179f
C27217 hold54/a_49_47# comp0.B\[0\] 0
C27218 _0521_/a_299_297# VPWR 0.20337f
C27219 _0320_ _1008_/a_27_47# 0
C27220 _0963_/a_285_47# control0.count\[1\] 0.002f
C27221 comp0.B\[3\] _1062_/a_193_47# 0
C27222 _0179_ acc0.A\[1\] 0
C27223 _0500_/a_27_47# _0199_ 0.02418f
C27224 hold20/a_285_47# control0.count\[3\] 0.00612f
C27225 _0998_/a_193_47# _0347_ 0
C27226 _0533_/a_109_47# _0181_ 0
C27227 _0399_ clknet_1_0__leaf__0457_ 0
C27228 _0232_ _0315_ 0
C27229 _0424_ _0425_ 0.17085f
C27230 _0181_ hold71/a_285_47# 0
C27231 _0387_ _0181_ 0.04934f
C27232 hold23/a_391_47# _0197_ 0.03389f
C27233 clknet_1_1__leaf__0463_ net231 0.0026f
C27234 _1030_/a_27_47# hold62/a_49_47# 0.01435f
C27235 _0361_ _0326_ 0
C27236 input28/a_75_212# B[5] 0.18905f
C27237 _0498_/a_149_47# _0159_ 0.00123f
C27238 _0084_ _0986_/a_466_413# 0.01443f
C27239 _0445_ _0986_/a_891_413# 0
C27240 clknet_1_1__leaf__0460_ net114 0
C27241 _0254_ _0255_ 0.15306f
C27242 acc0.A\[21\] VPWR 1.37458f
C27243 hold97/a_49_47# acc0.A\[27\] 0
C27244 hold96/a_285_47# _1024_/a_27_47# 0
C27245 hold96/a_49_47# _1024_/a_193_47# 0
C27246 _0592_/a_150_297# _0756_/a_47_47# 0
C27247 _1053_/a_193_47# net9 0
C27248 _1038_/a_891_413# _0136_ 0.02507f
C27249 net172 _0553_/a_240_47# 0
C27250 _0311_ _0392_ 0
C27251 _0257_ _0826_/a_27_53# 0
C27252 net150 _1005_/a_592_47# 0
C27253 _0120_ _1005_/a_1059_315# 0
C27254 net190 _1028_/a_1017_47# 0.00183f
C27255 _0452_ net149 0
C27256 _0404_ _0787_/a_80_21# 0
C27257 _0195_ net100 0
C27258 clknet_1_0__leaf__0465_ A[6] 0.11739f
C27259 clknet_1_1__leaf__0462_ _1008_/a_193_47# 0.00384f
C27260 hold42/a_391_47# pp[9] 0
C27261 _0715_/a_27_47# _0819_/a_299_297# 0
C27262 _0955_/a_32_297# _0213_ 0.00517f
C27263 _1032_/a_27_47# _0565_/a_240_47# 0
C27264 _1032_/a_1059_315# _0565_/a_51_297# 0
C27265 _0573_/a_27_47# _0216_ 0.00446f
C27266 _0449_ _0447_ 0.38872f
C27267 VPWR _1046_/a_634_159# 0.17654f
C27268 acc0.A\[31\] _1013_/a_891_413# 0.00233f
C27269 net162 _1013_/a_466_413# 0
C27270 _0736_/a_56_297# clknet_0__0462_ 0
C27271 _1022_/a_27_47# _1022_/a_891_413# 0.03224f
C27272 _1022_/a_193_47# _1022_/a_1059_315# 0.03405f
C27273 _1022_/a_634_159# _1022_/a_466_413# 0.23992f
C27274 _1003_/a_592_47# clknet_1_0__leaf__0460_ 0.00107f
C27275 _0686_/a_219_297# _0318_ 0.14862f
C27276 _1021_/a_891_413# _0462_ 0
C27277 _1052_/a_27_47# _0525_/a_299_297# 0
C27278 _1052_/a_193_47# _0525_/a_81_21# 0
C27279 _1059_/a_592_47# acc0.A\[15\] 0
C27280 hold58/a_49_47# net28 0
C27281 _1008_/a_1059_315# _0318_ 0
C27282 _0272_ _0986_/a_27_47# 0.00232f
C27283 net98 _0352_ 0
C27284 clknet_1_0__leaf__0461_ acc0.A\[18\] 0.57648f
C27285 _0957_/a_32_297# _0474_ 0.1707f
C27286 _1018_/a_975_413# _0116_ 0.0013f
C27287 net104 net219 0
C27288 _0957_/a_220_297# comp0.B\[6\] 0.00169f
C27289 hold38/a_285_47# clknet_1_1__leaf__0463_ 0.01036f
C27290 _0338_ acc0.A\[30\] 0.08935f
C27291 _1055_/a_1059_315# _1055_/a_891_413# 0.31086f
C27292 _1055_/a_193_47# _1055_/a_975_413# 0
C27293 _1055_/a_466_413# _1055_/a_381_47# 0.03733f
C27294 _1008_/a_466_413# net94 0
C27295 clknet_0__0459_ acc0.A\[14\] 0.30991f
C27296 _0466_ control0.count\[0\] 0.39142f
C27297 _0278_ VPWR 0.62411f
C27298 hold74/a_285_47# clknet_0__0461_ 0
C27299 hold24/a_49_47# hold24/a_391_47# 0.00188f
C27300 _1020_/a_592_47# _0118_ 0.00188f
C27301 net53 _1025_/a_1017_47# 0
C27302 net121 comp0.B\[5\] 0
C27303 _0559_/a_512_297# _0208_ 0
C27304 _0771_/a_215_297# _0771_/a_298_297# 0.07178f
C27305 hold14/a_285_47# _1036_/a_27_47# 0.00329f
C27306 hold14/a_49_47# _1036_/a_193_47# 0
C27307 net89 hold12/a_49_47# 0.05946f
C27308 _1003_/a_27_47# _1003_/a_561_413# 0.0027f
C27309 _1003_/a_634_159# _1003_/a_891_413# 0.03684f
C27310 _1003_/a_193_47# _1003_/a_381_47# 0.09503f
C27311 hold97/a_391_47# _0321_ 0
C27312 hold97/a_49_47# _0364_ 0.00695f
C27313 net23 _0474_ 0
C27314 clkbuf_1_0__f__0464_/a_110_47# acc0.A\[3\] 0.00242f
C27315 _0855_/a_299_297# _1019_/a_891_413# 0
C27316 VPWR _0245_ 0.95438f
C27317 _1001_/a_1059_315# _0399_ 0
C27318 hold64/a_285_47# _0195_ 0
C27319 _0466_ _0974_/a_544_297# 0.00394f
C27320 VPWR _0970_/a_285_47# 0
C27321 clknet_0__0463_ _0180_ 0.01465f
C27322 _0212_ _0955_/a_32_297# 0
C27323 net185 _0955_/a_114_297# 0.00123f
C27324 hold81/a_391_47# net228 0.13562f
C27325 hold55/a_391_47# _0584_/a_27_297# 0
C27326 _0165_ clkbuf_1_1__f_clk/a_110_47# 0.01655f
C27327 acc0.A\[21\] net48 0.68045f
C27328 net224 clknet_0__0462_ 0
C27329 _0556_/a_68_297# B[5] 0
C27330 VPWR _0747_/a_297_297# 0.01117f
C27331 _1054_/a_634_159# net15 0.01015f
C27332 _1054_/a_27_47# _0191_ 0.00557f
C27333 _0525_/a_81_21# net12 0.02063f
C27334 clknet_1_1__leaf__0460_ _0365_ 0.03218f
C27335 _1032_/a_1017_47# comp0.B\[0\] 0
C27336 _0997_/a_381_47# _0219_ 0
C27337 _0764_/a_81_21# _0384_ 0.0041f
C27338 _0465_ _0843_/a_68_297# 0.00535f
C27339 _0216_ _0779_/a_510_47# 0
C27340 _1004_/a_466_413# _0347_ 0
C27341 _1004_/a_27_47# _0352_ 0.14888f
C27342 net230 net9 0
C27343 output55/a_27_47# _0332_ 0
C27344 net8 clknet_1_1__leaf__0457_ 0.00104f
C27345 clknet_1_1__leaf__0461_ _0405_ 0
C27346 net77 acc0.A\[15\] 0
C27347 _0174_ _0913_/a_27_47# 0.04193f
C27348 _0440_ acc0.A\[5\] 0.22075f
C27349 A[10] clknet_1_1__leaf__0465_ 0
C27350 _0362_ clkbuf_0__0462_/a_110_47# 0
C27351 _1054_/a_634_159# _1053_/a_1059_315# 0.0057f
C27352 _1054_/a_193_47# _1053_/a_891_413# 0.00399f
C27353 VPWR hold9/a_285_47# 0.27418f
C27354 _0799_/a_209_297# _0799_/a_209_47# 0
C27355 _0799_/a_80_21# _0799_/a_303_47# 0.01146f
C27356 _0088_ net62 0.00318f
C27357 pp[27] hold15/a_49_47# 0
C27358 input22/a_75_212# net10 0.00257f
C27359 _0598_/a_297_47# VPWR 0.00356f
C27360 VPWR _0987_/a_193_47# 0.3401f
C27361 _0256_ _0636_/a_59_75# 0.00248f
C27362 net144 _1057_/a_1059_315# 0.00915f
C27363 _1058_/a_466_413# net189 0.0173f
C27364 _0219_ _0668_/a_79_21# 0
C27365 hold64/a_49_47# clknet_0__0457_ 0
C27366 _0516_/a_109_297# _0186_ 0.05677f
C27367 clknet_1_0__leaf__0459_ net238 0
C27368 _0664_/a_79_21# _0296_ 0.13654f
C27369 _0333_ _0350_ 0
C27370 _0347_ hold81/a_285_47# 0
C27371 _0985_/a_1059_315# _0269_ 0
C27372 _1000_/a_193_47# _0244_ 0.00395f
C27373 _1000_/a_27_47# _0386_ 0.00143f
C27374 _1000_/a_891_413# _0769_/a_299_297# 0
C27375 VPWR _1029_/a_193_47# 0.36889f
C27376 _0367_ _0360_ 0.02448f
C27377 _0315_ _0321_ 0
C27378 _0128_ _0220_ 0
C27379 hold59/a_49_47# clknet_1_0__leaf__0461_ 0.00456f
C27380 _0982_/a_27_47# _0453_ 0
C27381 _0982_/a_466_413# _0452_ 0
C27382 clkbuf_0__0460_/a_110_47# _0315_ 0.00658f
C27383 hold61/a_49_47# hold61/a_285_47# 0.22264f
C27384 clknet_1_0__leaf_clk _1064_/a_891_413# 0
C27385 _1048_/a_27_47# _1048_/a_1059_315# 0.04875f
C27386 _1048_/a_193_47# _1048_/a_466_413# 0.07482f
C27387 _0117_ _0264_ 0
C27388 _1015_/a_891_413# _0178_ 0
C27389 _0399_ _0850_/a_68_297# 0
C27390 _0548_/a_51_297# _0202_ 0
C27391 _0357_ _0353_ 0
C27392 VPWR B[2] 0.47644f
C27393 clknet_1_1__leaf__0465_ _0508_/a_299_297# 0.0021f
C27394 _0232_ _0742_/a_81_21# 0
C27395 net99 acc0.A\[30\] 0
C27396 _0622_/a_193_47# _0086_ 0
C27397 _0563_/a_149_47# _0214_ 0.00154f
C27398 _0548_/a_512_297# _0138_ 0
C27399 _0555_/a_512_297# VPWR 0.00744f
C27400 _0506_/a_384_47# net229 0.01004f
C27401 _0312_ _1007_/a_193_47# 0
C27402 hold11/a_49_47# hold11/a_285_47# 0.22264f
C27403 VPWR _1033_/a_975_413# 0.00464f
C27404 net129 _0543_/a_68_297# 0
C27405 clknet_1_0__leaf__0465_ _1049_/a_975_413# 0
C27406 hold59/a_285_47# net47 0.00426f
C27407 _0389_ _0246_ 0
C27408 _0535_/a_68_297# _0172_ 0.00158f
C27409 hold55/a_285_47# VPWR 0.29093f
C27410 acc0.A\[7\] _0434_ 0
C27411 _0470_ clknet_0_clk 0
C27412 _0783_/a_510_47# _0218_ 0
C27413 net61 VPWR 1.28809f
C27414 _0598_/a_297_47# net48 0.00381f
C27415 _0494_/a_27_47# _0173_ 0.21005f
C27416 _0183_ _0854_/a_297_297# 0
C27417 net192 _0156_ 0.04997f
C27418 _0642_/a_215_297# acc0.A\[6\] 0
C27419 _0546_/a_51_297# _0204_ 0
C27420 _0205_ _0544_/a_51_297# 0
C27421 hold76/a_49_47# hold76/a_285_47# 0.22264f
C27422 _0151_ _1054_/a_466_413# 0
C27423 net211 clknet_1_0__leaf__0461_ 0.00975f
C27424 hold57/a_285_47# hold57/a_391_47# 0.41909f
C27425 _0349_ _0722_/a_297_297# 0.00274f
C27426 _1010_/a_466_413# _1010_/a_592_47# 0.00553f
C27427 _1010_/a_634_159# _1010_/a_1017_47# 0
C27428 _0179_ net77 0
C27429 clknet_1_0__leaf__0462_ _1004_/a_592_47# 0
C27430 hold55/a_391_47# _1015_/a_634_159# 0
C27431 hold55/a_49_47# _1015_/a_1059_315# 0.0037f
C27432 _1056_/a_1059_315# _0514_/a_27_297# 0
C27433 clkbuf_1_0__f__0460_/a_110_47# _0350_ 0.02858f
C27434 _0978_/a_27_297# _0978_/a_373_47# 0.01338f
C27435 _1040_/a_466_413# _1040_/a_381_47# 0.03733f
C27436 _1040_/a_193_47# _1040_/a_975_413# 0
C27437 _1040_/a_1059_315# _1040_/a_891_413# 0.31086f
C27438 _0795_/a_299_297# _0795_/a_384_47# 0
C27439 _0453_ _0446_ 0
C27440 _0305_ acc0.A\[16\] 0.3755f
C27441 _0230_ _0225_ 0.147f
C27442 _0146_ _1048_/a_592_47# 0.00164f
C27443 hold19/a_285_47# _0399_ 0
C27444 _0250_ _0350_ 0.44805f
C27445 _0216_ _1027_/a_466_413# 0.03044f
C27446 _0195_ _1027_/a_891_413# 0
C27447 VPWR _0165_ 0.45218f
C27448 _0279_ _0801_/a_113_47# 0
C27449 _0259_ _0345_ 0.00338f
C27450 _1002_/a_975_413# _0183_ 0
C27451 _0328_ _0312_ 0.13763f
C27452 VPWR _1019_/a_634_159# 0.17531f
C27453 _0303_ net228 0
C27454 net96 _1009_/a_27_47# 0
C27455 net39 output40/a_27_47# 0
C27456 net213 _0222_ 0
C27457 net1 _0760_/a_377_297# 0
C27458 clknet_1_0__leaf__0462_ output48/a_27_47# 0
C27459 acc0.A\[14\] _0996_/a_1059_315# 0.01288f
C27460 _0537_/a_150_297# _1045_/a_27_47# 0
C27461 _0537_/a_68_297# _1045_/a_193_47# 0
C27462 _1067_/a_1059_315# _1067_/a_891_413# 0.31086f
C27463 _1067_/a_193_47# _1067_/a_975_413# 0
C27464 _1067_/a_466_413# _1067_/a_381_47# 0.03733f
C27465 control0.state\[0\] _0468_ 0.34326f
C27466 net9 _0987_/a_381_47# 0.00987f
C27467 _0174_ _0172_ 0.31863f
C27468 _0821_/a_113_47# net65 0
C27469 _1001_/a_634_159# _0345_ 0.00845f
C27470 _0137_ comp0.B\[10\] 0
C27471 _0179_ _0656_/a_59_75# 0
C27472 _0462_ _0614_/a_183_297# 0
C27473 _1071_/a_27_47# _0169_ 0.11082f
C27474 _0346_ _0992_/a_891_413# 0
C27475 _1050_/a_27_47# _0172_ 0
C27476 _1072_/a_891_413# _1071_/a_1059_315# 0
C27477 _0985_/a_466_413# _0529_/a_27_297# 0
C27478 _0985_/a_634_159# _0529_/a_109_297# 0
C27479 _0487_ _0175_ 0
C27480 hold90/a_49_47# _0345_ 0
C27481 _0149_ hold83/a_391_47# 0
C27482 _1004_/a_193_47# _0757_/a_150_297# 0
C27483 _0120_ _0592_/a_68_297# 0
C27484 _1009_/a_1059_315# _1009_/a_1017_47# 0
C27485 control0.state\[1\] _1002_/a_27_47# 0
C27486 net65 _0989_/a_891_413# 0.03803f
C27487 _0717_/a_80_21# _0717_/a_209_297# 0.06257f
C27488 _0252_ _0989_/a_634_159# 0.03106f
C27489 _0989_/a_634_159# _0989_/a_381_47# 0
C27490 clknet_1_0__leaf__0462_ hold29/a_285_47# 0.01481f
C27491 clknet_1_0__leaf__0459_ _0245_ 0.00353f
C27492 net228 _0281_ 0
C27493 _0228_ _0460_ 0
C27494 _0544_/a_51_297# _1042_/a_193_47# 0.00155f
C27495 _0248_ _0616_/a_292_297# 0
C27496 _0181_ _0986_/a_27_47# 0.00103f
C27497 net101 _0457_ 0.21217f
C27498 _0372_ _0616_/a_78_199# 0
C27499 _0717_/a_303_47# _0335_ 0.00165f
C27500 clkbuf_1_1__f__0465_/a_110_47# _0294_ 0
C27501 _0967_/a_215_297# control0.sh 0
C27502 _0476_ _1066_/a_1017_47# 0
C27503 _0992_/a_634_159# _0992_/a_381_47# 0
C27504 net24 _0563_/a_240_47# 0.05778f
C27505 _0695_/a_80_21# clknet_0__0462_ 0
C27506 _0648_/a_27_297# _0399_ 0.00439f
C27507 clkbuf_1_0__f__0457_/a_110_47# _0749_/a_299_297# 0
C27508 _0606_/a_465_297# VPWR 0
C27509 VPWR _1045_/a_27_47# 0.6336f
C27510 VPWR _1053_/a_561_413# 0.00292f
C27511 net54 _0739_/a_215_47# 0.00662f
C27512 clkbuf_1_0__f__0458_/a_110_47# _0841_/a_79_21# 0
C27513 net226 control0.count\[1\] 0.04311f
C27514 hold10/a_391_47# control0.reset 0
C27515 _1014_/a_561_413# acc0.A\[0\] 0
C27516 _0959_/a_217_297# comp0.B\[6\] 0
C27517 hold94/a_49_47# hold94/a_391_47# 0.00188f
C27518 net71 _0186_ 0.14614f
C27519 _0996_/a_561_413# _0094_ 0
C27520 net54 _0352_ 0.30837f
C27521 _0261_ _0219_ 0.00563f
C27522 _0573_/a_27_47# net100 0
C27523 hold10/a_285_47# _0465_ 0.01309f
C27524 hold76/a_391_47# _0461_ 0.00867f
C27525 _0935_/a_27_47# _1061_/a_466_413# 0.00102f
C27526 hold10/a_391_47# _1061_/a_891_413# 0.00107f
C27527 _0983_/a_891_413# net219 0.00166f
C27528 _0983_/a_27_47# _0116_ 0
C27529 _1061_/a_27_47# _1061_/a_1059_315# 0.04885f
C27530 _1061_/a_193_47# _1061_/a_466_413# 0.08301f
C27531 _0476_ comp0.B\[2\] 0.03009f
C27532 acc0.A\[4\] net9 0.19251f
C27533 _0688_/a_109_297# _0320_ 0.01197f
C27534 _0429_ _0087_ 0
C27535 _0626_/a_68_297# _0258_ 0.10609f
C27536 _0216_ _1026_/a_381_47# 0
C27537 _1007_/a_634_159# _0219_ 0
C27538 _1054_/a_27_47# input11/a_75_212# 0
C27539 clknet_1_1__leaf__0459_ pp[14] 0
C27540 _0319_ _0737_/a_285_297# 0
C27541 _0689_/a_150_297# _0321_ 0.00199f
C27542 _1065_/a_193_47# _1063_/a_27_47# 0
C27543 _0817_/a_266_47# _0288_ 0
C27544 acc0.A\[16\] _0675_/a_150_297# 0
C27545 _0648_/a_109_297# _0277_ 0
C27546 clknet_1_1__leaf__0458_ _0826_/a_27_53# 0.00645f
C27547 _0190_ _0988_/a_1059_315# 0
C27548 acc0.A\[10\] net37 0.29834f
C27549 _0504_/a_27_47# _0458_ 0
C27550 _0113_ net17 0
C27551 net199 _0574_/a_27_297# 0.06686f
C27552 clkbuf_0__0459_/a_110_47# hold82/a_285_47# 0
C27553 clkbuf_1_0__f__0459_/a_110_47# _1016_/a_891_413# 0
C27554 hold2/a_391_47# _1047_/a_193_47# 0
C27555 _0387_ clknet_1_1__leaf__0461_ 0.00141f
C27556 _1020_/a_975_413# acc0.A\[20\] 0
C27557 _0217_ _1014_/a_1059_315# 0.07424f
C27558 _0559_/a_51_297# net25 0
C27559 acc0.A\[27\] _0685_/a_150_297# 0
C27560 _0787_/a_80_21# _0419_ 0.08178f
C27561 _1042_/a_891_413# net195 0
C27562 _1042_/a_1059_315# net19 0
C27563 _0977_/a_75_212# _1069_/a_634_159# 0
C27564 _0260_ _0447_ 0.06067f
C27565 _1065_/a_634_159# clknet_1_0__leaf__0457_ 0
C27566 _0803_/a_68_297# _0218_ 0.18433f
C27567 _0182_ _0530_/a_299_297# 0
C27568 _0197_ hold71/a_391_47# 0
C27569 _0530_/a_81_21# net218 0
C27570 net119 _0175_ 0
C27571 _0404_ _0402_ 0
C27572 clkbuf_0__0463_/a_110_47# net201 0
C27573 _0539_/a_68_297# _0539_/a_150_297# 0.00477f
C27574 _0984_/a_975_413# acc0.A\[15\] 0
C27575 clknet_1_0__leaf__0458_ _0181_ 0.0018f
C27576 net76 _0990_/a_27_47# 0.22704f
C27577 _1069_/a_193_47# _1069_/a_592_47# 0.00135f
C27578 _1069_/a_466_413# _1069_/a_561_413# 0.00772f
C27579 _1069_/a_634_159# _1069_/a_975_413# 0
C27580 VPWR _1028_/a_381_47# 0.07326f
C27581 net44 hold62/a_49_47# 0
C27582 _0469_ _0163_ 0
C27583 VPWR _0812_/a_215_47# 0.0021f
C27584 _0718_/a_377_297# pp[30] 0
C27585 B[13] net18 0
C27586 _0243_ net219 0
C27587 VPWR _0514_/a_27_297# 0.26401f
C27588 clknet_0__0465_ _0990_/a_193_47# 0.0021f
C27589 _1059_/a_634_159# acc0.A\[13\] 0.00117f
C27590 hold69/a_285_47# _0359_ 0
C27591 pp[9] net16 0.01634f
C27592 net10 net19 0.02976f
C27593 pp[16] hold78/a_49_47# 0
C27594 _0954_/a_114_297# comp0.B\[12\] 0.01222f
C27595 _0131_ control0.sh 0
C27596 _0225_ _0236_ 0.04856f
C27597 _0200_ net180 0
C27598 _1041_/a_1059_315# _1040_/a_27_47# 0.00227f
C27599 _1041_/a_193_47# _1040_/a_466_413# 0
C27600 _1041_/a_466_413# _1040_/a_193_47# 0
C27601 _1031_/a_1059_315# _0220_ 0.04046f
C27602 _1031_/a_466_413# _0336_ 0
C27603 B[8] B[14] 0.18164f
C27604 hold66/a_391_47# _0369_ 0.04262f
C27605 net213 _0762_/a_297_297# 0
C27606 hold66/a_49_47# _0383_ 0
C27607 net69 _0451_ 0
C27608 _0399_ _1017_/a_634_159# 0
C27609 hold85/a_391_47# _0466_ 0
C27610 pp[8] _0515_/a_81_21# 0
C27611 net3 acc0.A\[11\] 0.00698f
C27612 net124 net153 0
C27613 _0782_/a_27_47# _0345_ 0
C27614 _1030_/a_1059_315# net209 0
C27615 _1027_/a_27_47# _1026_/a_27_47# 0.00315f
C27616 net205 net186 0
C27617 _0386_ acc0.A\[19\] 0
C27618 _0596_/a_59_75# _0183_ 0.00326f
C27619 VPWR _0512_/a_109_297# 0.17647f
C27620 _1039_/a_27_47# _0207_ 0
C27621 _1018_/a_466_413# clknet_0__0461_ 0.00129f
C27622 _1018_/a_381_47# clkbuf_1_0__f__0461_/a_110_47# 0
C27623 _0804_/a_79_21# _0399_ 0.10858f
C27624 _0176_ _0544_/a_240_47# 0
C27625 _0349_ output56/a_27_47# 0.04354f
C27626 _0624_/a_145_75# _0218_ 0
C27627 net180 comp0.B\[8\] 0.11245f
C27628 _1002_/a_1059_315# _0181_ 0
C27629 _0218_ acc0.A\[18\] 0.21786f
C27630 _0480_ _0978_/a_109_47# 0
C27631 _0416_ _0286_ 0
C27632 _0217_ _1022_/a_27_47# 0
C27633 _1034_/a_891_413# _0176_ 0
C27634 clknet_1_1__leaf__0462_ _0318_ 0.00683f
C27635 acc0.A\[16\] _0181_ 0.56878f
C27636 _0231_ _0380_ 0.0033f
C27637 _0323_ _0460_ 0
C27638 hold75/a_49_47# _0450_ 0.02395f
C27639 hold75/a_285_47# _0446_ 0
C27640 _0462_ _0391_ 0
C27641 _0198_ acc0.A\[15\] 0
C27642 _0474_ _0213_ 0.00167f
C27643 _0275_ acc0.A\[9\] 0.05236f
C27644 _1022_/a_634_159# net151 0.00368f
C27645 VPWR net132 0.51255f
C27646 _0645_/a_285_47# _0276_ 0
C27647 clknet_1_1__leaf__0463_ _0565_/a_245_297# 0
C27648 _1065_/a_27_47# _1062_/a_891_413# 0
C27649 net87 _1019_/a_27_47# 0.00879f
C27650 clknet_1_0__leaf__0459_ _1019_/a_634_159# 0.00867f
C27651 _0348_ acc0.A\[30\] 0
C27652 _0992_/a_1059_315# _0421_ 0
C27653 _1018_/a_193_47# _0264_ 0
C27654 net47 _0219_ 0.02476f
C27655 net199 _1025_/a_634_159# 0
C27656 _0994_/a_1059_315# _0994_/a_891_413# 0.31086f
C27657 _0994_/a_193_47# _0994_/a_975_413# 0
C27658 _0994_/a_466_413# _0994_/a_381_47# 0.03733f
C27659 _1020_/a_891_413# clknet_1_0__leaf__0457_ 0.0011f
C27660 _0259_ _0819_/a_81_21# 0.00214f
C27661 _0275_ _0986_/a_592_47# 0
C27662 hold12/a_285_47# _0460_ 0.00167f
C27663 _0779_/a_79_21# _0396_ 0.17954f
C27664 _0287_ net217 0
C27665 VPWR hold5/a_391_47# 0.18329f
C27666 _0289_ _0422_ 0.03352f
C27667 clkbuf_0__0462_/a_110_47# _0324_ 0.17882f
C27668 _1055_/a_381_47# net179 0.13615f
C27669 VPWR _0739_/a_297_297# 0.01248f
C27670 _1023_/a_27_47# pp[23] 0
C27671 _1023_/a_634_159# net51 0.00281f
C27672 _0337_ _0195_ 0
C27673 _0305_ _0288_ 0
C27674 hold22/a_391_47# _1053_/a_193_47# 0
C27675 _1003_/a_891_413# net89 0
C27676 _1003_/a_1059_315# _0101_ 0.06877f
C27677 net36 _1047_/a_381_47# 0.01269f
C27678 _0954_/a_220_297# _0202_ 0.00132f
C27679 _0648_/a_109_297# _0298_ 0
C27680 net36 _0472_ 0.01926f
C27681 hold33/a_285_47# _0540_/a_51_297# 0
C27682 _0647_/a_47_47# net80 0
C27683 _0459_ _0611_/a_68_297# 0.01048f
C27684 _0372_ _0384_ 0.09139f
C27685 clknet_0__0463_ _0498_/a_51_297# 0
C27686 _0207_ _1040_/a_975_413# 0
C27687 _0183_ _0216_ 0.05954f
C27688 _1039_/a_27_47# _1039_/a_1059_315# 0.04718f
C27689 _1039_/a_193_47# _1039_/a_466_413# 0.07482f
C27690 clkbuf_0__0461_/a_110_47# _0347_ 0.03249f
C27691 _0257_ _0640_/a_215_297# 0.16052f
C27692 hold33/a_49_47# net173 0
C27693 _0197_ _0529_/a_373_47# 0
C27694 _1020_/a_466_413# _0457_ 0.00255f
C27695 net46 _0757_/a_68_297# 0.00467f
C27696 _0212_ _0474_ 0
C27697 _0343_ _0425_ 0
C27698 comp0.B\[13\] _0172_ 0.00539f
C27699 _0279_ _0672_/a_79_21# 0
C27700 net193 net180 0.00181f
C27701 comp0.B\[2\] clkbuf_0__0463_/a_110_47# 0
C27702 net140 net15 0
C27703 _0985_/a_634_159# net170 0
C27704 _0087_ clknet_1_1__leaf__0458_ 0.00242f
C27705 _0346_ _0809_/a_299_297# 0.00363f
C27706 _0257_ _0989_/a_975_413# 0
C27707 _0172_ _1046_/a_193_47# 0.03506f
C27708 _0498_/a_245_297# clknet_1_1__leaf__0457_ 0.00245f
C27709 _1049_/a_27_47# _0196_ 0
C27710 _0987_/a_27_47# _0523_/a_299_297# 0
C27711 _1026_/a_27_47# _1026_/a_466_413# 0.27314f
C27712 _1026_/a_193_47# _1026_/a_634_159# 0.12729f
C27713 net33 _1062_/a_1059_315# 0
C27714 _0646_/a_47_47# input5/a_75_212# 0.0012f
C27715 _0985_/a_193_47# clknet_1_0__leaf__0458_ 0.00674f
C27716 _1021_/a_27_47# clknet_1_0__leaf__0460_ 0.05234f
C27717 acc0.A\[31\] acc0.A\[30\] 0
C27718 net23 _1065_/a_592_47# 0.00247f
C27719 net140 _1053_/a_1059_315# 0.00242f
C27720 net169 _1053_/a_466_413# 0
C27721 clknet_1_1__leaf__0459_ _0408_ 0
C27722 _0714_/a_51_297# _0567_/a_27_297# 0
C27723 net220 hold73/a_391_47# 0.15379f
C27724 _0982_/a_634_159# _0399_ 0
C27725 _0385_ hold73/a_285_47# 0.04193f
C27726 _0222_ _0618_/a_510_47# 0.00248f
C27727 _0257_ _0465_ 0.00818f
C27728 clknet_1_0__leaf__0461_ _0611_/a_150_297# 0
C27729 clknet_0_clk _0485_ 0
C27730 _0179_ _0198_ 0.04456f
C27731 VPWR _0792_/a_303_47# 0
C27732 _0217_ _1067_/a_634_159# 0
C27733 _0183_ _1067_/a_27_47# 0
C27734 _1024_/a_634_159# _1024_/a_592_47# 0
C27735 _0726_/a_51_297# acc0.A\[28\] 0
C27736 net45 hold72/a_49_47# 0.01262f
C27737 net227 _0723_/a_27_413# 0
C27738 _0355_ _0723_/a_207_413# 0
C27739 VPWR _0431_ 0.62575f
C27740 _0426_ _0423_ 0
C27741 _0718_/a_377_297# _0339_ 0
C27742 B[9] _1042_/a_381_47# 0
C27743 _1021_/a_891_413# _1020_/a_193_47# 0
C27744 _0452_ net206 0
C27745 _0375_ _0600_/a_103_199# 0
C27746 _0234_ _0600_/a_337_297# 0
C27747 _1036_/a_27_47# B[2] 0
C27748 net61 _0835_/a_493_297# 0
C27749 hold97/a_49_47# hold97/a_285_47# 0.22264f
C27750 output43/a_27_47# _0997_/a_27_47# 0
C27751 _0574_/a_27_297# VPWR 0.21513f
C27752 _0514_/a_373_47# clknet_1_1__leaf__0465_ 0.00238f
C27753 VPWR _0659_/a_68_297# 0.18319f
C27754 _0786_/a_80_21# _0992_/a_27_47# 0
C27755 _0644_/a_285_47# acc0.A\[13\] 0.04434f
C27756 _0182_ _1049_/a_1059_315# 0
C27757 _0180_ _1049_/a_466_413# 0
C27758 comp0.B\[2\] _1032_/a_381_47# 0
C27759 _0601_/a_150_297# net51 0
C27760 _0540_/a_51_297# net20 0.12239f
C27761 _0540_/a_149_47# _0202_ 0.00154f
C27762 _0080_ _0452_ 0.00219f
C27763 _0953_/a_32_297# _1040_/a_193_47# 0
C27764 clk _1064_/a_381_47# 0.00226f
C27765 _0949_/a_145_75# net1 0.00293f
C27766 control0.add _0771_/a_27_413# 0
C27767 _1048_/a_891_413# _1048_/a_1017_47# 0.00617f
C27768 _1048_/a_634_159# net134 0
C27769 _0712_/a_561_47# _0220_ 0
C27770 _1034_/a_592_47# clknet_1_1__leaf__0463_ 0
C27771 net126 _0550_/a_51_297# 0
C27772 net63 acc0.A\[6\] 0.02889f
C27773 _0096_ _0410_ 0
C27774 VPWR _0956_/a_304_297# 0.00424f
C27775 _0731_/a_299_297# _0250_ 0.08937f
C27776 _1068_/a_193_47# _0468_ 0.23469f
C27777 VPWR _1016_/a_561_413# 0.00213f
C27778 net211 _0218_ 0
C27779 _0343_ _1013_/a_193_47# 0.00762f
C27780 _1035_/a_1059_315# net24 0
C27781 _0339_ _0097_ 0
C27782 _1032_/a_1059_315# clkbuf_1_1__f_clk/a_110_47# 0
C27783 _0243_ _0352_ 0.84108f
C27784 _1016_/a_891_413# clkbuf_0__0461_/a_110_47# 0
C27785 _1015_/a_27_47# comp0.B\[15\] 0
C27786 _0200_ _0545_/a_150_297# 0
C27787 _0341_ _0708_/a_68_297# 0.01708f
C27788 _0710_/a_109_297# net60 0
C27789 _1060_/a_1059_315# _0219_ 0
C27790 input33/a_75_212# input17/a_75_212# 0.01223f
C27791 _0172_ _0987_/a_27_47# 0
C27792 _0804_/a_215_47# _0404_ 0.00219f
C27793 _0478_ _0468_ 0
C27794 _0343_ _0432_ 0
C27795 _0137_ _0177_ 0
C27796 _0539_/a_68_297# net21 0.02349f
C27797 clkbuf_1_0__f__0457_/a_110_47# hold73/a_49_47# 0
C27798 net152 net198 0.05918f
C27799 _0490_ _0974_/a_79_199# 0
C27800 _0607_/a_27_297# acc0.A\[17\] 0.10569f
C27801 _0151_ net169 0
C27802 clknet_0__0465_ _0438_ 0.0015f
C27803 _0643_/a_103_199# _0447_ 0
C27804 comp0.B\[1\] _1015_/a_891_413# 0.0038f
C27805 input19/a_75_212# net128 0
C27806 pp[30] net162 0.00517f
C27807 _0183_ net247 0.45606f
C27808 _1051_/a_634_159# _0522_/a_27_297# 0
C27809 _0206_ _0545_/a_68_297# 0.00521f
C27810 hold16/a_285_47# _0336_ 0.0653f
C27811 clkbuf_1_0__f__0460_/a_110_47# _1006_/a_634_159# 0.00144f
C27812 hold69/a_391_47# _0371_ 0.00576f
C27813 _1056_/a_1059_315# _0189_ 0.02769f
C27814 hold55/a_285_47# _0113_ 0.00207f
C27815 hold69/a_49_47# _0104_ 0
C27816 hold6/a_49_47# _0139_ 0.31254f
C27817 _1040_/a_381_47# net174 0.12469f
C27818 hold26/a_285_47# _0200_ 0.00302f
C27819 _0195_ _0319_ 0
C27820 hold18/a_49_47# _0181_ 0
C27821 _0622_/a_109_47# acc0.A\[8\] 0
C27822 clknet_1_0__leaf__0465_ _1054_/a_381_47# 0
C27823 _0480_ net164 0.09293f
C27824 _0292_ _0291_ 0.30064f
C27825 _0249_ _1006_/a_466_413# 0
C27826 _0250_ _1006_/a_634_159# 0
C27827 _0273_ _0827_/a_109_297# 0
C27828 net154 net11 0.03951f
C27829 _1072_/a_634_159# _1072_/a_592_47# 0
C27830 _0216_ net156 0.07676f
C27831 VPWR _0757_/a_150_297# 0.00135f
C27832 _0891_/a_27_47# clknet_1_0__leaf__0457_ 0.22437f
C27833 clknet_1_1__leaf__0460_ _0223_ 0
C27834 _0841_/a_215_47# _0444_ 0.07179f
C27835 _0188_ net37 0.02277f
C27836 _0316_ clkbuf_0__0462_/a_110_47# 0.00217f
C27837 _0172_ comp0.B\[9\] 0.61429f
C27838 VPWR net105 0.48036f
C27839 hold39/a_285_47# clkbuf_1_1__f__0463_/a_110_47# 0
C27840 _0146_ clknet_1_1__leaf__0457_ 0.00412f
C27841 _0640_/a_215_297# _0640_/a_392_297# 0.00419f
C27842 _0640_/a_109_53# _0640_/a_297_297# 0
C27843 VPWR _0326_ 0.74742f
C27844 _1013_/a_27_47# net60 0.00389f
C27845 _0854_/a_79_21# net165 0
C27846 VPWR _1025_/a_634_159# 0.18294f
C27847 hold49/a_285_47# hold51/a_285_47# 0.00214f
C27848 _0772_/a_215_47# _0345_ 0.0094f
C27849 _0422_ _0418_ 0
C27850 clknet_1_1__leaf__0457_ _0492_/a_27_47# 0.01147f
C27851 net105 _1015_/a_466_413# 0
C27852 net214 _0186_ 0
C27853 _0538_/a_51_297# clknet_0__0464_ 0.00283f
C27854 _1012_/a_634_159# _0722_/a_79_21# 0
C27855 VPWR hold95/a_391_47# 0.18882f
C27856 _0592_/a_150_297# _0374_ 0
C27857 clknet_1_1__leaf__0460_ _1006_/a_1059_315# 0.00294f
C27858 _0217_ _1024_/a_466_413# 0.00165f
C27859 _0288_ _0181_ 0
C27860 _0179_ clknet_1_1__leaf__0464_ 0
C27861 _1004_/a_381_47# _0380_ 0
C27862 _0717_/a_209_47# _0348_ 0
C27863 hold75/a_285_47# net61 0
C27864 _0997_/a_634_159# _0997_/a_592_47# 0
C27865 _0640_/a_392_297# _0465_ 0
C27866 _1037_/a_193_47# net24 0
C27867 clknet_1_1__leaf__0459_ _0290_ 0
C27868 _0329_ clknet_0__0462_ 0
C27869 net216 _0462_ 0.00479f
C27870 _0204_ _1042_/a_891_413# 0.00349f
C27871 net198 _1042_/a_466_413# 0.01212f
C27872 net18 _1042_/a_634_159# 0.00683f
C27873 _0568_/a_27_297# hold95/a_49_47# 0
C27874 _0517_/a_81_21# acc0.A\[9\] 0
C27875 VPWR _1051_/a_592_47# 0
C27876 _0349_ _1010_/a_466_413# 0.00553f
C27877 net247 acc0.A\[15\] 0.57364f
C27878 _0356_ _0354_ 0.00119f
C27879 hold7/a_391_47# net154 0.13426f
C27880 _0280_ _0399_ 0.0348f
C27881 net190 acc0.A\[25\] 0
C27882 _0402_ _0419_ 0.36982f
C27883 _0959_/a_217_297# hold84/a_285_47# 0.00196f
C27884 _0959_/a_80_21# hold84/a_391_47# 0
C27885 _0783_/a_215_47# _0347_ 0.05298f
C27886 clknet_0__0458_ _0445_ 0.01284f
C27887 _0982_/a_27_47# _0345_ 0.00142f
C27888 net106 _0584_/a_27_297# 0
C27889 _1045_/a_1059_315# net196 0
C27890 _0793_/a_512_297# _0408_ 0
C27891 _0340_ clknet_1_1__leaf__0461_ 0
C27892 net45 clknet_0__0461_ 0.14048f
C27893 _0606_/a_215_297# _0754_/a_51_297# 0
C27894 _1027_/a_634_159# _1027_/a_381_47# 0
C27895 net185 comp0.B\[4\] 0.18553f
C27896 _0741_/a_109_297# _0367_ 0.01216f
C27897 _0253_ net212 0
C27898 _0181_ _0247_ 0
C27899 net193 hold26/a_285_47# 0.00143f
C27900 _0996_/a_891_413# net41 0.0044f
C27901 VPWR _1032_/a_1059_315# 0.40053f
C27902 comp0.B\[3\] B[2] 0
C27903 _1061_/a_891_413# _1061_/a_1017_47# 0.00617f
C27904 clknet_1_0__leaf__0465_ _0522_/a_27_297# 0.01034f
C27905 _1061_/a_634_159# net147 0
C27906 _0305_ _1009_/a_1059_315# 0
C27907 net51 _0377_ 0.00114f
C27908 net36 net149 0.11259f
C27909 _0798_/a_199_47# _0297_ 0
C27910 _0482_ _0976_/a_505_21# 0
C27911 _0555_/a_51_297# comp0.B\[5\] 0.12337f
C27912 net66 _0990_/a_1017_47# 0.00213f
C27913 acc0.A\[8\] _0990_/a_592_47# 0.00112f
C27914 _0225_ _0380_ 0
C27915 clknet_0__0457_ hold40/a_391_47# 0.03025f
C27916 hold10/a_49_47# clknet_1_0__leaf__0464_ 0.00189f
C27917 _0216_ acc0.A\[26\] 0.11148f
C27918 net93 _0219_ 0.00189f
C27919 _0982_/a_27_47# hold2/a_49_47# 0.00693f
C27920 _0340_ _1030_/a_193_47# 0
C27921 _0346_ clknet_1_0__leaf__0457_ 0.05263f
C27922 _0960_/a_27_47# _1071_/a_193_47# 0.0013f
C27923 _1035_/a_466_413# _1035_/a_561_413# 0.00772f
C27924 _1035_/a_634_159# _1035_/a_975_413# 0
C27925 _0399_ net235 0.06141f
C27926 acc0.A\[27\] _0570_/a_27_297# 0
C27927 _0571_/a_27_297# net190 0
C27928 _1035_/a_193_47# B[15] 0
C27929 net238 _0345_ 0.00232f
C27930 _0470_ _1065_/a_27_47# 0
C27931 _1053_/a_193_47# A[7] 0
C27932 comp0.B\[15\] _0215_ 0
C27933 _1000_/a_27_47# _0240_ 0
C27934 _1000_/a_466_413# _0247_ 0.01125f
C27935 _0243_ net207 0
C27936 _0183_ net100 0
C27937 _1000_/a_27_47# _0369_ 0
C27938 hold7/a_49_47# hold7/a_285_47# 0.22264f
C27939 _0977_/a_75_212# clknet_1_0__leaf_clk 0.04266f
C27940 _0412_ _0798_/a_199_47# 0.00179f
C27941 _0413_ _0798_/a_113_297# 0.00157f
C27942 net162 _0339_ 0.06586f
C27943 _0464_ _0144_ 0.00159f
C27944 _0289_ _0423_ 0.38263f
C27945 _0292_ _0290_ 0.4857f
C27946 _1013_/a_381_47# clknet_1_1__leaf__0461_ 0
C27947 net33 B[4] 0.00126f
C27948 _0446_ _0345_ 0.12235f
C27949 _1048_/a_466_413# acc0.A\[15\] 0
C27950 _0727_/a_193_47# acc0.A\[29\] 0
C27951 VPWR _0269_ 1.32583f
C27952 net134 _0138_ 0
C27953 _1010_/a_1059_315# _0701_/a_80_21# 0.00111f
C27954 _0718_/a_47_47# _0718_/a_377_297# 0.00899f
C27955 _0252_ _0988_/a_193_47# 0
C27956 VPWR _0546_/a_51_297# 0.47108f
C27957 _1054_/a_1059_315# acc0.A\[8\] 0.09464f
C27958 acc0.A\[16\] clknet_1_1__leaf__0461_ 0.64828f
C27959 _0569_/a_27_297# net191 0.00593f
C27960 _0569_/a_109_297# net115 0
C27961 acc0.A\[29\] _1029_/a_381_47# 0
C27962 _0294_ _0219_ 0.0255f
C27963 _1011_/a_634_159# _0726_/a_51_297# 0
C27964 net78 clknet_1_1__leaf__0465_ 0.01712f
C27965 _1069_/a_561_413# _0167_ 0
C27966 _1069_/a_975_413# clknet_1_0__leaf_clk 0
C27967 _1069_/a_1059_315# control0.count\[0\] 0.15941f
C27968 _1016_/a_27_47# net102 0.22366f
C27969 clknet_0__0465_ clknet_1_1__leaf__0465_ 0.00429f
C27970 VPWR acc0.A\[28\] 1.08066f
C27971 _1033_/a_27_47# _1065_/a_193_47# 0
C27972 _0455_ _0181_ 0.0636f
C27973 net64 _0436_ 0
C27974 _0179_ net247 0.09757f
C27975 net145 acc0.A\[13\] 0
C27976 VPWR _0189_ 0.34251f
C27977 _0233_ _0223_ 0.07635f
C27978 hold33/a_285_47# hold33/a_391_47# 0.41909f
C27979 VPWR net209 0.39107f
C27980 _1041_/a_193_47# net174 0
C27981 hold25/a_391_47# clknet_1_0__leaf__0463_ 0.03253f
C27982 _0835_/a_215_47# clkbuf_1_0__f__0465_/a_110_47# 0
C27983 _0399_ net103 0
C27984 acc0.A\[27\] hold50/a_49_47# 0.32015f
C27985 net125 _1061_/a_634_159# 0.01029f
C27986 output42/a_27_47# _0218_ 0.01295f
C27987 clknet_1_1__leaf__0458_ net154 0.13831f
C27988 _0488_ _0484_ 0.12651f
C27989 hold64/a_285_47# _0183_ 0.01786f
C27990 _0577_/a_373_47# net150 0
C27991 _0577_/a_27_297# _0183_ 0.24301f
C27992 _0577_/a_109_297# acc0.A\[22\] 0.0199f
C27993 _0577_/a_109_47# _0217_ 0.00145f
C27994 _0640_/a_215_297# clknet_1_1__leaf__0458_ 0.01169f
C27995 _0149_ net9 0
C27996 _0750_/a_109_47# _0219_ 0
C27997 _0181_ _0505_/a_109_297# 0.04565f
C27998 hold15/a_49_47# hold15/a_391_47# 0.00188f
C27999 net183 net21 0.17229f
C28000 _0173_ hold84/a_391_47# 0
C28001 VPWR _0381_ 0.76579f
C28002 net106 _1015_/a_634_159# 0
C28003 _0524_/a_109_297# net12 0.01154f
C28004 _0673_/a_337_297# net228 0
C28005 pp[25] net155 0
C28006 _1065_/a_634_159# _0160_ 0
C28007 hold75/a_49_47# _0637_/a_56_297# 0.00184f
C28008 clknet_1_0__leaf__0459_ net105 0.03687f
C28009 _0241_ clknet_1_0__leaf__0460_ 0
C28010 _0465_ clknet_1_1__leaf__0458_ 0.0488f
C28011 comp0.B\[12\] _0542_/a_51_297# 0
C28012 comp0.B\[11\] _0542_/a_245_297# 0
C28013 _0995_/a_27_47# output41/a_27_47# 0
C28014 _0800_/a_51_297# _0405_ 0.00247f
C28015 _0550_/a_240_47# B[7] 0
C28016 _0982_/a_466_413# net36 0.02627f
C28017 _0520_/a_27_297# _0520_/a_109_47# 0.00393f
C28018 VPWR hold72/a_49_47# 0.26998f
C28019 net211 _0099_ 0.10961f
C28020 net45 _1013_/a_466_413# 0.00962f
C28021 hold24/a_285_47# clknet_1_0__leaf__0463_ 0
C28022 _1018_/a_27_47# _0247_ 0
C28023 _0780_/a_117_297# _0240_ 0
C28024 _0238_ _0617_/a_68_297# 0.17742f
C28025 _0179_ _1048_/a_466_413# 0.01456f
C28026 _0461_ clknet_1_0__leaf__0461_ 0.05669f
C28027 _0260_ _0275_ 0.04878f
C28028 net203 _0215_ 0
C28029 net109 net51 0.06446f
C28030 _1043_/a_193_47# _1042_/a_27_47# 0.00755f
C28031 _1043_/a_27_47# _1042_/a_193_47# 0.00755f
C28032 net45 _0607_/a_373_47# 0
C28033 _1055_/a_27_47# net74 0
C28034 _0769_/a_81_21# VPWR 0.20254f
C28035 clknet_1_0__leaf__0463_ input7/a_75_212# 0.01292f
C28036 _1019_/a_1059_315# _0399_ 0
C28037 _0278_ _0345_ 0
C28038 _0993_/a_634_159# _0993_/a_592_47# 0
C28039 _0816_/a_150_297# acc0.A\[9\] 0
C28040 hold87/a_49_47# VPWR 0.28399f
C28041 _1039_/a_891_413# _1039_/a_1017_47# 0.00617f
C28042 _0186_ _0434_ 0.0219f
C28043 _1039_/a_634_159# net125 0
C28044 _0182_ net175 0.13641f
C28045 _0236_ _0462_ 0.04388f
C28046 _0257_ _0254_ 0.06729f
C28047 _0118_ _0457_ 0.00751f
C28048 _0280_ _0295_ 0
C28049 net59 _0999_/a_1059_315# 0
C28050 _0218_ _0611_/a_150_297# 0
C28051 _1038_/a_1059_315# _0463_ 0
C28052 _0973_/a_109_297# clknet_1_0__leaf__0460_ 0
C28053 _0580_/a_27_297# _0580_/a_373_47# 0.01338f
C28054 _0673_/a_253_297# _0347_ 0.00128f
C28055 net204 _0494_/a_27_47# 0
C28056 A[12] net3 0.67758f
C28057 _0310_ net43 0
C28058 pp[27] clknet_1_1__leaf__0460_ 0
C28059 _0850_/a_68_297# _0346_ 0.00567f
C28060 net48 _0381_ 0.18145f
C28061 _0465_ _0263_ 0.02094f
C28062 clknet_1_1__leaf__0463_ _0564_/a_68_297# 0.06849f
C28063 _1026_/a_193_47# net112 0.016f
C28064 _1026_/a_1059_315# _1026_/a_1017_47# 0
C28065 _1059_/a_634_159# VPWR 0.18201f
C28066 _0985_/a_466_413# _0449_ 0
C28067 net107 hold93/a_285_47# 0.00224f
C28068 _0465_ _1047_/a_27_47# 0.0147f
C28069 _0286_ net246 0
C28070 _0172_ clkbuf_1_0__f__0465_/a_110_47# 0
C28071 _0999_/a_27_47# _0779_/a_79_21# 0.00214f
C28072 _0697_/a_472_297# _0324_ 0.0044f
C28073 net179 clknet_1_1__leaf__0458_ 0
C28074 _0172_ hold5/a_285_47# 0
C28075 _0472_ _1061_/a_27_47# 0.01309f
C28076 net225 _0567_/a_27_297# 0.0054f
C28077 net58 _0261_ 0.56362f
C28078 acc0.A\[2\] _0263_ 0.06811f
C28079 _0181_ _1009_/a_1059_315# 0
C28080 _0718_/a_129_47# _0348_ 0.00213f
C28081 comp0.B\[7\] clknet_1_1__leaf__0457_ 0
C28082 _0331_ _0324_ 0
C28083 _1024_/a_891_413# acc0.A\[24\] 0.00378f
C28084 _0455_ _1018_/a_27_47# 0
C28085 _0454_ _1018_/a_193_47# 0
C28086 clknet_1_1__leaf__0463_ clknet_1_1__leaf_clk 0.05962f
C28087 _0290_ _0655_/a_215_53# 0
C28088 _0294_ _0746_/a_81_21# 0.00975f
C28089 output54/a_27_47# _0571_/a_27_297# 0.01849f
C28090 hold30/a_285_47# net50 0.00127f
C28091 net66 input16/a_75_212# 0
C28092 hold36/a_391_47# _1044_/a_27_47# 0
C28093 clkbuf_0__0465_/a_110_47# acc0.A\[6\] 0
C28094 _0527_/a_109_47# _0186_ 0.00153f
C28095 clknet_1_1__leaf__0464_ _0141_ 0.0104f
C28096 _0195_ _0333_ 0.13662f
C28097 _0343_ _0360_ 0
C28098 _0642_/a_27_413# _0087_ 0
C28099 _0662_/a_299_297# _0662_/a_384_47# 0
C28100 hold36/a_49_47# net184 0.00439f
C28101 hold36/a_285_47# net131 0.00145f
C28102 _0255_ acc0.A\[4\] 0.02621f
C28103 _0174_ _1040_/a_193_47# 0.0354f
C28104 control0.state\[0\] _0978_/a_109_297# 0
C28105 _1037_/a_27_47# _1037_/a_1059_315# 0.04875f
C28106 _1037_/a_193_47# _1037_/a_466_413# 0.07482f
C28107 pp[16] _0997_/a_381_47# 0
C28108 _0402_ _0992_/a_193_47# 0
C28109 _0180_ _0147_ 0.02206f
C28110 acc0.A\[22\] _0756_/a_129_47# 0
C28111 hold4/a_285_47# hold4/a_391_47# 0.41909f
C28112 _0147_ net218 0.00472f
C28113 comp0.B\[10\] _1040_/a_466_413# 0
C28114 _0369_ _0507_/a_27_297# 0.01093f
C28115 acc0.A\[7\] _0186_ 0.09268f
C28116 hold48/a_391_47# net20 0
C28117 clknet_1_0__leaf__0462_ _0743_/a_51_297# 0.00171f
C28118 _0186_ _0989_/a_1059_315# 0
C28119 _0785_/a_81_21# _0401_ 0.13496f
C28120 _0785_/a_299_297# _0290_ 0
C28121 _1029_/a_193_47# _0345_ 0
C28122 hold48/a_285_47# hold48/a_391_47# 0.41909f
C28123 _0501_/a_27_47# net201 0
C28124 control0.state\[1\] _1067_/a_466_413# 0
C28125 net126 _0172_ 0.00234f
C28126 _0102_ net50 0.00238f
C28127 _0562_/a_68_297# _0171_ 0.00145f
C28128 _1041_/a_193_47# _1041_/a_592_47# 0
C28129 _1041_/a_466_413# _1041_/a_561_413# 0.00772f
C28130 _1041_/a_634_159# _1041_/a_975_413# 0
C28131 _0228_ _0373_ 0
C28132 VPWR _0991_/a_381_47# 0.07725f
C28133 _0504_/a_27_47# acc0.A\[1\] 0.05497f
C28134 input25/a_75_212# net26 0.00103f
C28135 _1054_/a_193_47# _0180_ 0.01991f
C28136 _0243_ _0769_/a_299_297# 0.03297f
C28137 _0390_ _0769_/a_81_21# 0
C28138 net31 net18 0
C28139 output56/a_27_47# _1030_/a_193_47# 0
C28140 VPWR _0600_/a_103_199# 0.42723f
C28141 _1057_/a_27_47# net2 0
C28142 hold42/a_285_47# A[11] 0
C28143 _0176_ _1043_/a_1059_315# 0.00117f
C28144 _0337_ hold15/a_49_47# 0
C28145 net58 _0509_/a_27_47# 0
C28146 _0456_ acc0.A\[1\] 0.06297f
C28147 _1039_/a_27_47# _0472_ 0.02801f
C28148 _1039_/a_634_159# _0473_ 0.00861f
C28149 _0625_/a_59_75# _0989_/a_27_47# 0.00126f
C28150 _0467_ _1072_/a_27_47# 0
C28151 _0465_ clknet_1_0__leaf__0461_ 0.00211f
C28152 _0569_/a_109_47# acc0.A\[28\] 0.00275f
C28153 pp[9] net142 0
C28154 _1051_/a_634_159# _0193_ 0
C28155 net61 _0345_ 0
C28156 hold86/a_285_47# _0219_ 0.0604f
C28157 clkbuf_1_0__f__0460_/a_110_47# net92 0
C28158 clkbuf_1_1__f_clk/a_110_47# _0468_ 0
C28159 net139 net13 0.08682f
C28160 _0369_ acc0.A\[19\] 0.55178f
C28161 acc0.A\[29\] hold62/a_285_47# 0
C28162 _0593_/a_113_47# _0222_ 0
C28163 clknet_0__0457_ acc0.A\[19\] 0.00158f
C28164 _0461_ _0585_/a_27_297# 0
C28165 hold97/a_391_47# _0738_/a_68_297# 0.00107f
C28166 VPWR _1011_/a_634_159# 0.18059f
C28167 _0234_ _0762_/a_215_47# 0.00235f
C28168 _0251_ _0831_/a_285_47# 0.00313f
C28169 _0250_ net92 0
C28170 VPWR clknet_0__0461_ 2.03873f
C28171 pp[2] _0827_/a_27_47# 0
C28172 _0963_/a_35_297# _1069_/a_466_413# 0.0019f
C28173 hold65/a_285_47# net248 0.00176f
C28174 _0453_ _0269_ 0
C28175 _1030_/a_27_47# net57 0
C28176 net215 _0352_ 0
C28177 A[10] _0515_/a_81_21# 0.05736f
C28178 _1019_/a_634_159# _0345_ 0.02136f
C28179 _0985_/a_27_47# _0846_/a_512_297# 0
C28180 _0361_ _1009_/a_193_47# 0
C28181 output67/a_27_47# _1058_/a_27_47# 0.00104f
C28182 net58 net47 0
C28183 clknet_1_0__leaf__0459_ hold72/a_49_47# 0.00619f
C28184 net105 _0113_ 0
C28185 _1012_/a_466_413# _0110_ 0.00473f
C28186 _1012_/a_891_413# _0351_ 0.00119f
C28187 clknet_1_1__leaf__0460_ _0216_ 0.00677f
C28188 acc0.A\[22\] net110 0
C28189 _0217_ _0122_ 0.072f
C28190 _0413_ net41 0
C28191 _1051_/a_193_47# _0150_ 0
C28192 _0190_ net235 0
C28193 _0218_ _0799_/a_80_21# 0.02122f
C28194 net155 net197 0
C28195 _0578_/a_109_47# VPWR 0
C28196 _0644_/a_285_47# VPWR 0.00144f
C28197 net101 _0130_ 0
C28198 _0227_ clknet_1_0__leaf__0460_ 0.15618f
C28199 net135 net10 0.02261f
C28200 _0369_ _0249_ 0.02814f
C28201 _0579_/a_109_47# _0352_ 0
C28202 VPWR _1044_/a_1017_47# 0
C28203 _0146_ _1049_/a_634_159# 0.00368f
C28204 _0198_ _1049_/a_891_413# 0
C28205 _0239_ net43 0.02782f
C28206 _0684_/a_59_75# _0322_ 0.04665f
C28207 _0262_ _0261_ 0.22982f
C28208 hold35/a_391_47# _0189_ 0.00231f
C28209 comp0.B\[11\] input19/a_75_212# 0.01169f
C28210 _0661_/a_277_297# acc0.A\[9\] 0
C28211 _0661_/a_109_297# _0288_ 0
C28212 _0292_ _0656_/a_59_75# 0
C28213 _0096_ _0352_ 0.04236f
C28214 _0243_ _0392_ 0.00344f
C28215 _0316_ _0331_ 0
C28216 _0684_/a_59_75# _0327_ 0
C28217 _0095_ _0408_ 0
C28218 _1001_/a_1017_47# _0461_ 0
C28219 _0643_/a_337_297# _0272_ 0.00838f
C28220 _0643_/a_103_199# _0275_ 0.14175f
C28221 _0643_/a_253_297# _0274_ 0.00109f
C28222 _1027_/a_891_413# net156 0
C28223 _0606_/a_297_297# _0377_ 0
C28224 _0606_/a_215_297# _0219_ 0.00659f
C28225 _0606_/a_109_53# net241 0.00132f
C28226 _0606_/a_465_297# _0345_ 0
C28227 pp[17] _0341_ 0
C28228 net61 clkload1/a_268_47# 0.00152f
C28229 clknet_1_0__leaf__0463_ _0138_ 0.08824f
C28230 _1030_/a_891_413# _0707_/a_75_199# 0
C28231 _1030_/a_1059_315# _0707_/a_201_297# 0
C28232 net1 _1014_/a_193_47# 0
C28233 clknet_1_0__leaf__0463_ _0211_ 0.00268f
C28234 net239 hold92/a_391_47# 0.13065f
C28235 VPWR _0082_ 0.5138f
C28236 _0957_/a_32_297# _0957_/a_114_297# 0.01439f
C28237 _0293_ _0986_/a_193_47# 0
C28238 net101 _1019_/a_381_47# 0
C28239 clkbuf_1_1__f__0460_/a_110_47# _0701_/a_80_21# 0.00295f
C28240 clknet_1_0__leaf__0465_ _0193_ 0.01437f
C28241 _0749_/a_299_297# _0248_ 0.06189f
C28242 _0749_/a_81_21# _0372_ 0.00164f
C28243 _0331_ _0347_ 0.07364f
C28244 _0636_/a_145_75# net170 0
C28245 _0462_ _0370_ 0.03971f
C28246 clknet_1_0__leaf__0462_ _1023_/a_975_413# 0
C28247 _0482_ _0466_ 0
C28248 net64 pp[4] 0.00425f
C28249 net133 _0465_ 0.04621f
C28250 _0582_/a_27_297# _0582_/a_373_47# 0.01338f
C28251 _0131_ _0474_ 0
C28252 clkload2/Y net135 0.00467f
C28253 net202 _1015_/a_1059_315# 0
C28254 _0478_ _1071_/a_466_413# 0
C28255 _1007_/a_193_47# _1007_/a_634_159# 0.11072f
C28256 _1052_/a_634_159# _1052_/a_466_413# 0.23992f
C28257 _1052_/a_193_47# _1052_/a_1059_315# 0.03405f
C28258 _1052_/a_27_47# _1052_/a_891_413# 0.03224f
C28259 _1007_/a_27_47# _1007_/a_466_413# 0.27314f
C28260 _0125_ net190 0.01028f
C28261 acc0.A\[27\] _0126_ 0.02704f
C28262 _0343_ net59 0
C28263 hold87/a_391_47# _0266_ 0.01645f
C28264 hold87/a_49_47# _0453_ 0
C28265 _1012_/a_634_159# acc0.A\[30\] 0
C28266 net186 _1034_/a_193_47# 0.20023f
C28267 _1015_/a_1059_315# clknet_1_1__leaf__0463_ 0
C28268 hold39/a_391_47# _1034_/a_381_47# 0.00119f
C28269 _0330_ _1010_/a_1059_315# 0
C28270 _0973_/a_27_297# hold93/a_49_47# 0.00966f
C28271 _1058_/a_27_47# _1058_/a_561_413# 0.0027f
C28272 _1058_/a_634_159# _1058_/a_891_413# 0.03684f
C28273 _1058_/a_193_47# _1058_/a_381_47# 0.09503f
C28274 VPWR _0702_/a_113_47# 0
C28275 _0098_ _0247_ 0
C28276 hold14/a_285_47# net24 0
C28277 hold14/a_391_47# B[1] 0.00139f
C28278 control0.state\[0\] _0480_ 0
C28279 _0312_ net216 0
C28280 _1051_/a_975_413# _0172_ 0
C28281 _0110_ net98 0.0018f
C28282 VPWR _0468_ 1.03719f
C28283 _0353_ _0723_/a_297_47# 0
C28284 _0212_ _1035_/a_27_47# 0
C28285 net185 _1035_/a_193_47# 0.00271f
C28286 _1050_/a_466_413# _0527_/a_109_297# 0
C28287 _0585_/a_27_297# _0465_ 0.00119f
C28288 _0680_/a_80_21# _0305_ 0.17204f
C28289 hold12/a_49_47# _0487_ 0.0163f
C28290 _0262_ _0509_/a_27_47# 0
C28291 _0718_/a_285_47# _0349_ 0.04779f
C28292 _0127_ net191 0.23754f
C28293 net97 _0726_/a_51_297# 0.00776f
C28294 _1011_/a_891_413# _0354_ 0
C28295 _1011_/a_466_413# net227 0
C28296 _1011_/a_1059_315# _0355_ 0.01331f
C28297 _1011_/a_27_47# _0109_ 0.09888f
C28298 VPWR _1013_/a_466_413# 0.25188f
C28299 net182 _0189_ 0.02246f
C28300 _1002_/a_193_47# VPWR 0.29753f
C28301 net236 _0482_ 0.00967f
C28302 _0983_/a_27_47# _0854_/a_79_21# 0.00574f
C28303 _0126_ _0364_ 0
C28304 _0538_/a_51_297# comp0.B\[14\] 0.09123f
C28305 _0831_/a_117_297# clknet_1_1__leaf__0458_ 0.00101f
C28306 clknet_1_0__leaf__0462_ output52/a_27_47# 0.00141f
C28307 _0812_/a_215_47# _0345_ 0
C28308 _0179_ net148 0.16139f
C28309 _0869_/a_27_47# _0459_ 0.11122f
C28310 net125 net147 0.08115f
C28311 net149 hold60/a_391_47# 0
C28312 _0398_ _1016_/a_1017_47# 0
C28313 _0476_ _0466_ 0
C28314 _0183_ _0120_ 0.0315f
C28315 comp0.B\[10\] _1061_/a_381_47# 0
C28316 _1027_/a_891_413# acc0.A\[26\] 0
C28317 _0174_ _0207_ 0.29153f
C28318 _0254_ clknet_1_1__leaf__0458_ 0.15729f
C28319 net58 _0988_/a_592_47# 0
C28320 hold13/a_49_47# net24 0
C28321 _0277_ _0405_ 0
C28322 _0300_ _0400_ 0
C28323 _0379_ net110 0.0032f
C28324 _0786_/a_217_297# _0786_/a_472_297# 0.00517f
C28325 _0786_/a_80_21# _0786_/a_300_47# 0.00997f
C28326 _1038_/a_381_47# _0176_ 0.00229f
C28327 _0233_ _0216_ 0
C28328 hold70/a_49_47# _0281_ 0
C28329 _0165_ _1065_/a_1059_315# 0.00125f
C28330 _0214_ _0208_ 0.04324f
C28331 _0550_/a_51_297# net8 0
C28332 _0461_ _0218_ 0.1749f
C28333 _0575_/a_109_297# _0216_ 0.02083f
C28334 _0974_/a_79_199# _0974_/a_544_297# 0.00594f
C28335 _0530_/a_299_297# _1048_/a_1059_315# 0
C28336 _0257_ _0625_/a_59_75# 0.11066f
C28337 net205 _1034_/a_466_413# 0
C28338 _0996_/a_381_47# clkbuf_0__0459_/a_110_47# 0
C28339 hold11/a_285_47# _1049_/a_27_47# 0
C28340 _0984_/a_193_47# VPWR 0.30925f
C28341 _0985_/a_466_413# _0260_ 0
C28342 net36 net206 0.03072f
C28343 clknet_1_0__leaf__0459_ clknet_0__0461_ 0.14053f
C28344 _0994_/a_466_413# _0218_ 0.00853f
C28345 _0550_/a_51_297# net32 0
C28346 net59 _1012_/a_381_47# 0
C28347 output66/a_27_47# pp[9] 0.02881f
C28348 net61 _0836_/a_68_297# 0
C28349 hold100/a_285_47# _0346_ 0
C28350 _0948_/a_109_297# clk 0
C28351 net17 hold93/a_49_47# 0.01533f
C28352 hold13/a_285_47# _1039_/a_634_159# 0
C28353 net211 _1019_/a_1017_47# 0
C28354 net111 _1026_/a_193_47# 0.00255f
C28355 _0995_/a_381_47# pp[14] 0
C28356 pp[27] output44/a_27_47# 0.00194f
C28357 net46 _0232_ 0
C28358 hold44/a_285_47# net114 0
C28359 _0520_/a_109_297# _0186_ 0.01244f
C28360 hold57/a_285_47# _0552_/a_68_297# 0
C28361 _0080_ net36 0.15569f
C28362 _1002_/a_193_47# net48 0
C28363 VPWR _1042_/a_891_413# 0.18134f
C28364 _1056_/a_466_413# acc0.A\[9\] 0.00172f
C28365 net61 net212 0.00821f
C28366 _0982_/a_634_159# _0346_ 0.01188f
C28367 acc0.A\[29\] _0350_ 0.00193f
C28368 clknet_0__0459_ _0276_ 0
C28369 _0518_/a_27_297# _0252_ 0.00231f
C28370 _0518_/a_373_47# net65 0
C28371 _0783_/a_79_21# clknet_0__0461_ 0
C28372 pp[26] _0572_/a_109_297# 0
C28373 VPWR _0763_/a_109_47# 0
C28374 net22 net134 0
C28375 _0395_ _0352_ 0.05396f
C28376 clknet_0__0460_ _1009_/a_466_413# 0
C28377 _1030_/a_634_159# acc0.A\[30\] 0.02347f
C28378 _0642_/a_298_297# _0252_ 0.05917f
C28379 _0273_ _0989_/a_27_47# 0
C28380 net150 hold73/a_285_47# 0
C28381 _0217_ hold73/a_49_47# 0
C28382 _0682_/a_68_297# _0366_ 0.05948f
C28383 hold89/a_285_47# _0466_ 0.04724f
C28384 hold89/a_391_47# _0488_ 0
C28385 _0231_ _0369_ 0
C28386 hold3/a_49_47# _0219_ 0.01687f
C28387 pp[27] _1030_/a_975_413# 0
C28388 _0988_/a_634_159# _0988_/a_1059_315# 0
C28389 _0988_/a_27_47# _0988_/a_381_47# 0.06222f
C28390 _0988_/a_193_47# _0988_/a_891_413# 0.19489f
C28391 clkbuf_1_1__f__0465_/a_110_47# _0291_ 0.08723f
C28392 _1039_/a_1059_315# _0174_ 0.0033f
C28393 VPWR _0560_/a_68_297# 0.15935f
C28394 _0984_/a_193_47# _0983_/a_381_47# 0
C28395 pp[18] _1013_/a_1059_315# 0
C28396 _0368_ _0315_ 0.07089f
C28397 _0279_ _0301_ 0
C28398 _0730_/a_510_47# _0357_ 0.0017f
C28399 _0699_/a_68_297# _0350_ 0.01064f
C28400 _0730_/a_79_21# _0108_ 0.06184f
C28401 _0730_/a_215_47# _0358_ 0.00557f
C28402 hold64/a_49_47# acc0.A\[19\] 0.33857f
C28403 _1041_/a_27_47# _0547_/a_68_297# 0.00109f
C28404 net1 _0369_ 0.24009f
C28405 _0580_/a_373_47# _0117_ 0
C28406 _0228_ _0761_/a_113_47# 0
C28407 _0343_ _0335_ 0
C28408 hold20/a_49_47# _0170_ 0
C28409 net10 _1043_/a_975_413# 0
C28410 clknet_0__0457_ net1 0.00605f
C28411 VPWR clkbuf_0__0458_/a_110_47# 1.26345f
C28412 clknet_1_0__leaf__0458_ clknet_1_1__leaf__0465_ 0.00144f
C28413 hold28/a_391_47# _0465_ 0
C28414 _0478_ _0978_/a_109_297# 0.00465f
C28415 _0629_/a_59_75# hold100/a_285_47# 0
C28416 _0695_/a_217_297# _0326_ 0.00262f
C28417 clkbuf_1_1__f__0461_/a_110_47# _0240_ 0
C28418 _0162_ _1064_/a_561_413# 0
C28419 _0485_ _1064_/a_1017_47# 0
C28420 _0207_ _0208_ 0
C28421 _0559_/a_512_297# clknet_1_1__leaf__0463_ 0
C28422 _0371_ _0219_ 0.00176f
C28423 net145 VPWR 0.37595f
C28424 _0982_/a_634_159# _0629_/a_59_75# 0
C28425 _0083_ _0449_ 0.00131f
C28426 _1001_/a_634_159# clknet_1_0__leaf__0457_ 0.01301f
C28427 acc0.A\[2\] hold28/a_391_47# 0
C28428 _0225_ _0592_/a_150_297# 0
C28429 input18/a_75_212# net18 0.10862f
C28430 _0999_/a_193_47# _0097_ 0.27001f
C28431 _0999_/a_466_413# _0396_ 0.00109f
C28432 _0880_/a_27_47# _1062_/a_1059_315# 0
C28433 clknet_1_0__leaf__0457_ _1062_/a_193_47# 0
C28434 _0473_ net147 0.04955f
C28435 _0356_ _0353_ 0.00268f
C28436 _0343_ net81 0.05719f
C28437 _0817_/a_266_47# _0424_ 0.09559f
C28438 clknet_1_1__leaf__0460_ _1009_/a_975_413# 0
C28439 _1035_/a_634_159# net27 0.00755f
C28440 net56 hold95/a_391_47# 0.06999f
C28441 clkbuf_1_1__f__0459_/a_110_47# hold91/a_285_47# 0
C28442 _0316_ _1008_/a_27_47# 0
C28443 clknet_1_1__leaf__0459_ net83 0.18775f
C28444 net46 _0616_/a_493_297# 0
C28445 input23/a_75_212# input27/a_75_212# 0
C28446 net195 net20 0.043f
C28447 A[14] output40/a_27_47# 0
C28448 _0266_ _0264_ 0.78922f
C28449 net15 _0087_ 0
C28450 _0191_ _0437_ 0
C28451 output54/a_27_47# _0125_ 0.03244f
C28452 net54 acc0.A\[27\] 0.12777f
C28453 hold48/a_285_47# net195 0.00984f
C28454 hold36/a_49_47# net130 0
C28455 _1038_/a_1059_315# clkbuf_1_0__f__0463_/a_110_47# 0
C28456 acc0.A\[20\] _0586_/a_27_47# 0.02166f
C28457 _0302_ acc0.A\[13\] 0.02719f
C28458 net236 hold89/a_285_47# 0.01127f
C28459 _0279_ _0994_/a_193_47# 0
C28460 _0278_ _0994_/a_27_47# 0
C28461 _0404_ _0400_ 0
C28462 _0298_ _0405_ 0.01546f
C28463 _0792_/a_303_47# _0345_ 0
C28464 _0347_ _1008_/a_27_47# 0.03756f
C28465 _0458_ _0219_ 0.0063f
C28466 _1037_/a_891_413# _1037_/a_1017_47# 0.00617f
C28467 _1037_/a_193_47# _0135_ 0.57068f
C28468 _0345_ _0431_ 0
C28469 acc0.A\[16\] clknet_1_1__leaf__0465_ 0
C28470 _0997_/a_1059_315# _0218_ 0.01211f
C28471 hold38/a_49_47# clkbuf_1_1__f__0463_/a_110_47# 0
C28472 _0195_ _0998_/a_891_413# 0.03343f
C28473 comp0.B\[10\] net174 0.12423f
C28474 _0369_ _0185_ 0
C28475 net231 _0951_/a_296_53# 0
C28476 _0164_ _0951_/a_209_311# 0
C28477 _0465_ _0848_/a_27_47# 0.00105f
C28478 pp[30] _1030_/a_1059_315# 0.01856f
C28479 net59 _1030_/a_381_47# 0
C28480 _0633_/a_109_297# _0265_ 0.0124f
C28481 VPWR _1005_/a_1017_47# 0
C28482 _0218_ _0465_ 0.03034f
C28483 _0680_/a_80_21# _0181_ 0
C28484 acc0.A\[15\] _0406_ 0.00954f
C28485 _0285_ _0786_/a_80_21# 0
C28486 hold89/a_391_47# _1064_/a_27_47# 0
C28487 VPWR _0152_ 0.21396f
C28488 VPWR net67 2.34487f
C28489 _0255_ _0350_ 0
C28490 _1039_/a_1059_315# _0208_ 0.00747f
C28491 _0985_/a_193_47# _0448_ 0
C28492 _0985_/a_1059_315# _0447_ 0.01177f
C28493 net54 _0364_ 0.26629f
C28494 _0959_/a_80_21# net23 0.09277f
C28495 _0121_ _1023_/a_891_413# 0
C28496 pp[12] _0994_/a_1059_315# 0.00814f
C28497 _1001_/a_193_47# _1001_/a_891_413# 0.19658f
C28498 _1001_/a_27_47# _1001_/a_381_47# 0.06222f
C28499 _1001_/a_634_159# _1001_/a_1059_315# 0
C28500 _0705_/a_59_75# hold80/a_285_47# 0
C28501 _0217_ _0181_ 0.2093f
C28502 _0607_/a_373_47# clknet_1_0__leaf__0459_ 0
C28503 hold76/a_391_47# net223 0.13415f
C28504 hold76/a_285_47# _0391_ 0
C28505 _1062_/a_27_47# _1062_/a_1059_315# 0.04875f
C28506 _1062_/a_193_47# _1062_/a_466_413# 0.07874f
C28507 net125 _0473_ 0
C28508 _0608_/a_27_47# acc0.A\[17\] 0.07406f
C28509 _1020_/a_27_47# _1032_/a_27_47# 0.07618f
C28510 _0670_/a_215_47# clkbuf_1_1__f__0459_/a_110_47# 0
C28511 _0341_ _0567_/a_109_297# 0.00482f
C28512 _0340_ _0567_/a_27_297# 0.05317f
C28513 clknet_1_0__leaf__0458_ _0452_ 0.00186f
C28514 _1011_/a_27_47# _0725_/a_80_21# 0
C28515 _0472_ _0953_/a_32_297# 0.37369f
C28516 _0473_ _0953_/a_220_297# 0
C28517 hold38/a_391_47# _0951_/a_209_311# 0
C28518 net44 net57 0
C28519 hold90/a_49_47# hold90/a_391_47# 0.00188f
C28520 _1003_/a_27_47# net49 0.00377f
C28521 _0575_/a_109_297# _1024_/a_193_47# 0
C28522 _0575_/a_27_297# _1024_/a_634_159# 0
C28523 clkbuf_1_1__f__0465_/a_110_47# _0290_ 0.04525f
C28524 net79 net246 0
C28525 _0183_ _0307_ 0
C28526 _1049_/a_891_413# _1048_/a_466_413# 0.00157f
C28527 _0227_ hold94/a_285_47# 0.06423f
C28528 net133 clknet_0__0464_ 0
C28529 _0758_/a_215_47# acc0.A\[23\] 0.0047f
C28530 _0461_ _0112_ 0
C28531 VPWR net97 0.40619f
C28532 _0572_/a_109_47# VPWR 0.00104f
C28533 VPWR _1006_/a_975_413# 0.00483f
C28534 _0459_ _1060_/a_193_47# 0
C28535 _0248_ hold73/a_49_47# 0
C28536 _0280_ _0346_ 0.04888f
C28537 _0309_ net43 0.0017f
C28538 _0284_ _0787_/a_80_21# 0.13135f
C28539 _0285_ _0787_/a_209_297# 0.06987f
C28540 hold43/a_285_47# _1029_/a_193_47# 0
C28541 hold43/a_391_47# _1029_/a_27_47# 0
C28542 _0963_/a_35_297# _0167_ 0
C28543 _0481_ _1069_/a_891_413# 0
C28544 _0963_/a_117_297# clknet_1_0__leaf_clk 0.00494f
C28545 net56 acc0.A\[28\] 0.41959f
C28546 _0363_ _0350_ 0.20255f
C28547 _0195_ _1030_/a_1017_47# 0
C28548 net35 net159 0.03425f
C28549 _0327_ _0723_/a_207_413# 0
C28550 net48 _1005_/a_1017_47# 0
C28551 _0336_ net239 0.00193f
C28552 VPWR _0986_/a_975_413# 0.00484f
C28553 clknet_1_1__leaf__0464_ _1043_/a_27_47# 0.10068f
C28554 _1039_/a_634_159# comp0.B\[8\] 0
C28555 _0714_/a_240_47# _0219_ 0.05978f
C28556 net105 _0345_ 0.09614f
C28557 _0343_ _0797_/a_207_413# 0.01774f
C28558 _0742_/a_81_21# _0368_ 0.17557f
C28559 acc0.A\[13\] net6 0.07119f
C28560 _0386_ _0462_ 0
C28561 _0186_ _0988_/a_466_413# 0
C28562 hold34/a_49_47# _0179_ 0
C28563 _0371_ _0746_/a_81_21# 0.11432f
C28564 _1004_/a_891_413# _0216_ 0
C28565 _0224_ _1022_/a_27_47# 0
C28566 _0221_ _0723_/a_27_413# 0
C28567 _0561_/a_51_297# _0561_/a_240_47# 0.03076f
C28568 VPWR _0616_/a_215_47# 0.01055f
C28569 _0216_ _0171_ 0.00189f
C28570 _1072_/a_27_47# _1068_/a_381_47# 0
C28571 _1072_/a_634_159# _1068_/a_1059_315# 0
C28572 _1072_/a_466_413# _1068_/a_466_413# 0
C28573 _1072_/a_193_47# _1068_/a_891_413# 0
C28574 _0476_ _1065_/a_634_159# 0
C28575 VPWR _0762_/a_79_21# 0.45205f
C28576 _0180_ acc0.A\[6\] 0.61402f
C28577 _0662_/a_299_297# _0294_ 0.00113f
C28578 _0662_/a_81_21# _0218_ 0
C28579 net105 hold2/a_49_47# 0
C28580 clkbuf_1_0__f__0461_/a_110_47# acc0.A\[18\] 0.15754f
C28581 _0346_ _0270_ 0
C28582 hold41/a_285_47# _0179_ 0.06479f
C28583 hold30/a_49_47# clknet_1_0__leaf__0460_ 0.00122f
C28584 _0957_/a_32_297# _0173_ 0.00823f
C28585 clknet_0__0464_ comp0.B\[10\] 0
C28586 _1036_/a_193_47# clknet_1_1__leaf__0463_ 0.06466f
C28587 VPWR _0707_/a_201_297# 0.19636f
C28588 _0330_ clkbuf_1_1__f__0460_/a_110_47# 0
C28589 _0478_ _0480_ 0.28622f
C28590 _1003_/a_1017_47# acc0.A\[21\] 0
C28591 _0343_ _0741_/a_109_297# 0
C28592 _0461_ _0099_ 0.00501f
C28593 _1035_/a_891_413# _0132_ 0
C28594 _0133_ _0561_/a_240_47# 0.0432f
C28595 _0248_ _0618_/a_297_297# 0
C28596 _1041_/a_27_47# net127 0.22867f
C28597 _0437_ clkbuf_1_0__f__0465_/a_110_47# 0
C28598 _1047_/a_634_159# _1047_/a_381_47# 0
C28599 net23 _0173_ 0
C28600 _1030_/a_1059_315# _0339_ 0
C28601 _1030_/a_891_413# _0338_ 0
C28602 comp0.B\[8\] _1040_/a_1017_47# 0
C28603 hold1/a_391_47# _0987_/a_1059_315# 0
C28604 hold1/a_285_47# _0987_/a_891_413# 0.00358f
C28605 _0957_/a_304_297# _0475_ 0.00218f
C28606 _0432_ acc0.A\[6\] 0
C28607 _0131_ _0563_/a_51_297# 0.13072f
C28608 _0664_/a_382_297# _0284_ 0.01494f
C28609 _0664_/a_297_47# _0285_ 0.00711f
C28610 clknet_1_0__leaf__0460_ _0352_ 0.07908f
C28611 _0133_ _0472_ 0
C28612 output56/a_27_47# _0354_ 0.0014f
C28613 _0195_ _0526_/a_27_47# 0.35678f
C28614 _0582_/a_373_47# _0115_ 0
C28615 net58 _0833_/a_297_297# 0
C28616 net36 comp0.B\[15\] 0.05829f
C28617 hold52/a_49_47# _0574_/a_109_297# 0.00197f
C28618 hold52/a_285_47# _0574_/a_27_297# 0
C28619 comp0.B\[5\] _0496_/a_27_47# 0.00338f
C28620 acc0.A\[7\] input12/a_75_212# 0
C28621 net234 _1014_/a_891_413# 0
C28622 _0797_/a_27_413# net5 0
C28623 _0217_ _1018_/a_27_47# 0.02544f
C28624 _0178_ control0.reset 0.00514f
C28625 _0570_/a_27_297# _0689_/a_68_297# 0
C28626 _0359_ _0318_ 0
C28627 _1007_/a_193_47# net93 0.0041f
C28628 _1007_/a_1059_315# _1007_/a_1017_47# 0
C28629 _1007_/a_27_47# _0105_ 0.09169f
C28630 _0464_ _0528_/a_81_21# 0
C28631 net243 _1004_/a_27_47# 0.00786f
C28632 _0177_ _0465_ 0.00248f
C28633 _0622_/a_109_47# _0369_ 0
C28634 clkbuf_1_1__f__0464_/a_110_47# _0473_ 0
C28635 _0837_/a_266_297# _0440_ 0.01473f
C28636 _0837_/a_81_21# _0441_ 0.21702f
C28637 _1058_/a_891_413# net144 0
C28638 _0195_ net9 0.00568f
C28639 hold39/a_391_47# comp0.B\[2\] 0
C28640 _0165_ hold93/a_49_47# 0.02865f
C28641 _0172_ _1044_/a_592_47# 0.00178f
C28642 hold69/a_391_47# _1006_/a_1059_315# 0.01554f
C28643 _0289_ _0369_ 0.05526f
C28644 _1020_/a_381_47# _0352_ 0
C28645 net197 _1027_/a_1059_315# 0.0011f
C28646 net190 _1027_/a_634_159# 0
C28647 net48 _0762_/a_79_21# 0.01152f
C28648 VPWR _0498_/a_512_297# 0.00738f
C28649 _0625_/a_59_75# clknet_1_1__leaf__0458_ 0.01172f
C28650 _0629_/a_59_75# _0858_/a_27_47# 0
C28651 _0223_ _0617_/a_150_297# 0
C28652 hold74/a_49_47# hold74/a_285_47# 0.22264f
C28653 _0557_/a_149_47# VPWR 0.00182f
C28654 _0219_ pp[14] 0
C28655 _0705_/a_59_75# _0220_ 0.10146f
C28656 _0734_/a_47_47# _0734_/a_129_47# 0.00369f
C28657 _1050_/a_381_47# net11 0.01376f
C28658 _0112_ _0465_ 0
C28659 _1003_/a_891_413# _0487_ 0
C28660 control0.state\[0\] _0951_/a_368_53# 0
C28661 control0.state\[1\] _0951_/a_296_53# 0
C28662 comp0.B\[12\] net198 0
C28663 comp0.B\[11\] net18 0.02363f
C28664 _0971_/a_81_21# _0181_ 0.06167f
C28665 clkbuf_0_clk/a_110_47# clk 0.31322f
C28666 _0574_/a_27_297# net52 0.00183f
C28667 _0225_ _0369_ 0
C28668 net45 _0339_ 0.06713f
C28669 _0294_ _0582_/a_109_297# 0
C28670 _0269_ _0345_ 0.63218f
C28671 net245 net6 0
C28672 _1061_/a_1059_315# comp0.B\[9\] 0
C28673 _0819_/a_81_21# _0659_/a_68_297# 0.00128f
C28674 _0459_ _0796_/a_79_21# 0
C28675 clkbuf_0_clk/a_110_47# _1063_/a_891_413# 0
C28676 net61 _0989_/a_891_413# 0.01209f
C28677 hold59/a_49_47# clkbuf_1_0__f__0461_/a_110_47# 0.00111f
C28678 acc0.A\[4\] hold1/a_49_47# 0
C28679 _0402_ _0420_ 0.07416f
C28680 clknet_0__0462_ hold90/a_285_47# 0.00108f
C28681 acc0.A\[28\] _0345_ 0.08291f
C28682 hold75/a_285_47# _0082_ 0
C28683 _0983_/a_193_47# _0081_ 0.25723f
C28684 _0286_ hold70/a_391_47# 0
C28685 _0288_ clknet_1_1__leaf__0465_ 0.01108f
C28686 _0983_/a_1059_315# _0454_ 0
C28687 _0983_/a_466_413# _0455_ 0
C28688 _0429_ pp[3] 0
C28689 _0312_ _0370_ 0.14819f
C28690 _0369_ _0436_ 0.00246f
C28691 _1059_/a_891_413# _0277_ 0
C28692 _0319_ acc0.A\[26\] 0.0134f
C28693 _0328_ net93 0.00113f
C28694 _1063_/a_193_47# _1063_/a_381_47# 0.09503f
C28695 _1063_/a_634_159# _1063_/a_891_413# 0.03684f
C28696 _1063_/a_27_47# _1063_/a_561_413# 0.00163f
C28697 acc0.A\[9\] _0088_ 0.0389f
C28698 net247 _0171_ 0
C28699 hold86/a_391_47# _0465_ 0.00646f
C28700 _0345_ net209 0.1207f
C28701 _0179_ _0513_/a_384_47# 0
C28702 hold19/a_285_47# net221 0
C28703 _1037_/a_1059_315# _0208_ 0.00268f
C28704 clknet_1_0__leaf__0463_ net22 0.06275f
C28705 clkbuf_1_1__f__0464_/a_110_47# _0186_ 0.00329f
C28706 _0115_ clknet_1_0__leaf__0461_ 0
C28707 _1063_/a_975_413# clknet_1_0__leaf__0457_ 0
C28708 net67 _0283_ 0.0347f
C28709 _0462_ _1006_/a_466_413# 0.00231f
C28710 hold86/a_285_47# net58 0.0974f
C28711 hold86/a_391_47# acc0.A\[2\] 0
C28712 _0172_ net8 0.05507f
C28713 _1039_/a_381_47# _0177_ 0
C28714 net125 _0497_/a_68_297# 0.07633f
C28715 _0183_ _0507_/a_109_297# 0.01712f
C28716 _0343_ _0790_/a_35_297# 0.01847f
C28717 _1028_/a_27_47# clknet_1_1__leaf__0462_ 0.05381f
C28718 _0172_ net32 0.304f
C28719 net46 _0771_/a_27_413# 0
C28720 hold74/a_391_47# net43 0
C28721 _0642_/a_215_297# _0831_/a_35_297# 0
C28722 _0820_/a_510_47# net66 0
C28723 net211 clkbuf_1_0__f__0461_/a_110_47# 0
C28724 _0221_ net115 0
C28725 pp[17] acc0.A\[30\] 0.00869f
C28726 _0663_/a_207_413# _0295_ 0.07343f
C28727 _0424_ _0181_ 0.00223f
C28728 _1011_/a_561_413# acc0.A\[29\] 0
C28729 _0570_/a_27_297# net112 0
C28730 _1004_/a_466_413# _1024_/a_466_413# 0
C28731 _1004_/a_27_47# _1024_/a_381_47# 0
C28732 VPWR _1010_/a_27_47# 0.72711f
C28733 net188 acc0.A\[10\] 0
C28734 _0369_ _0990_/a_592_47# 0
C28735 _0429_ _0273_ 0.05101f
C28736 _0576_/a_109_297# _0352_ 0
C28737 A[14] _0797_/a_207_413# 0
C28738 _0587_/a_27_47# _0339_ 0.00956f
C28739 _1060_/a_193_47# _1060_/a_381_47# 0.09503f
C28740 _1060_/a_634_159# _1060_/a_891_413# 0.03684f
C28741 _1060_/a_27_47# _1060_/a_561_413# 0.0027f
C28742 net18 _0202_ 0
C28743 net68 _0346_ 0
C28744 _1051_/a_193_47# _0527_/a_27_297# 0
C28745 _0513_/a_81_21# _0513_/a_384_47# 0.00138f
C28746 _0733_/a_222_93# _0319_ 0.14032f
C28747 _1028_/a_634_159# net94 0
C28748 _0432_ _0624_/a_59_75# 0
C28749 clkbuf_0__0457_/a_110_47# hold60/a_49_47# 0.02088f
C28750 _1051_/a_27_47# _0346_ 0
C28751 _0216_ _0456_ 0
C28752 _1070_/a_193_47# _0480_ 0
C28753 _1070_/a_27_47# net164 0
C28754 _0191_ _0252_ 0.03477f
C28755 clknet_0__0459_ _0369_ 0.20221f
C28756 net126 _1040_/a_193_47# 0.01325f
C28757 _1053_/a_193_47# net11 0.01046f
C28758 hold38/a_49_47# _0163_ 0.01096f
C28759 acc0.A\[12\] _0153_ 0
C28760 _0143_ _1050_/a_1059_315# 0.0301f
C28761 _0326_ net52 0.0034f
C28762 _1039_/a_891_413# _0555_/a_51_297# 0
C28763 output58/a_27_47# _0252_ 0
C28764 net203 _1065_/a_193_47# 0
C28765 _0988_/a_1059_315# net74 0
C28766 _0553_/a_245_297# _0174_ 0.00131f
C28767 _1067_/a_466_413# clknet_1_1__leaf_clk 0
C28768 pp[29] net227 0.03162f
C28769 _0787_/a_209_297# _0218_ 0.00179f
C28770 _0968_/a_193_297# net34 0
C28771 _0331_ _1011_/a_27_47# 0
C28772 _0984_/a_891_413# net69 0
C28773 VPWR _1009_/a_193_47# 0.29834f
C28774 _1053_/a_975_413# acc0.A\[7\] 0
C28775 _0315_ clknet_0__0460_ 0.06566f
C28776 _0857_/a_27_47# _1033_/a_27_47# 0
C28777 _1041_/a_1059_315# _0206_ 0.02358f
C28778 _1041_/a_891_413# comp0.B\[8\] 0
C28779 _0399_ _0264_ 0.01318f
C28780 _0982_/a_975_413# _0465_ 0
C28781 _0234_ net150 0
C28782 _0583_/a_27_297# _0583_/a_109_297# 0.17136f
C28783 VPWR _1014_/a_381_47# 0.06974f
C28784 _1071_/a_466_413# VPWR 0.25314f
C28785 _0203_ net19 0.0336f
C28786 net248 VPWR 0.52041f
C28787 clknet_1_0__leaf__0457_ _0772_/a_215_47# 0.00578f
C28788 _0984_/a_27_47# hold75/a_391_47# 0
C28789 _0984_/a_193_47# hold75/a_285_47# 0
C28790 hold39/a_49_47# VPWR 0.28254f
C28791 hold28/a_285_47# clknet_1_0__leaf__0464_ 0.00267f
C28792 acc0.A\[15\] _0507_/a_109_297# 0.00203f
C28793 net89 net240 0
C28794 net82 _1060_/a_891_413# 0
C28795 _0172_ _1042_/a_1059_315# 0
C28796 acc0.A\[27\] _0569_/a_109_297# 0
C28797 net55 _0318_ 0.03574f
C28798 hold59/a_285_47# acc0.A\[1\] 0
C28799 _1021_/a_975_413# _0460_ 0
C28800 net121 net27 0
C28801 _1021_/a_1017_47# clknet_1_0__leaf__0457_ 0
C28802 _0479_ _0978_/a_27_297# 0.00513f
C28803 acc0.A\[15\] hold82/a_49_47# 0.00334f
C28804 _0603_/a_68_297# _0603_/a_150_297# 0.00477f
C28805 net36 hold71/a_285_47# 0
C28806 _0080_ hold60/a_391_47# 0
C28807 hold20/a_49_47# net35 0.02799f
C28808 clkbuf_0__0462_/a_110_47# _0360_ 0.01302f
C28809 _0254_ _0218_ 0
C28810 _0258_ _0256_ 0.02242f
C28811 _0183_ net118 0
C28812 _0992_/a_466_413# net143 0
C28813 clkbuf_0__0464_/a_110_47# _1046_/a_1059_315# 0.01107f
C28814 clkbuf_1_1__f__0463_/a_110_47# _0565_/a_51_297# 0
C28815 _0309_ _0677_/a_129_47# 0
C28816 _0678_/a_68_297# acc0.A\[17\] 0
C28817 hold35/a_285_47# acc0.A\[9\] 0.01789f
C28818 _0285_ net144 0
C28819 _0217_ clknet_1_1__leaf__0461_ 0.00861f
C28820 hold79/a_285_47# control0.count\[0\] 0.00393f
C28821 _1008_/a_634_159# _0365_ 0
C28822 _1008_/a_27_47# _0106_ 0.10409f
C28823 _0313_ _0697_/a_217_297# 0.02013f
C28824 clknet_1_1__leaf__0465_ _0505_/a_109_297# 0
C28825 _0408_ _0219_ 0.04328f
C28826 _0258_ _0987_/a_1059_315# 0
C28827 _0780_/a_35_297# _0307_ 0
C28828 pp[30] VPWR 0.62281f
C28829 _0718_/a_47_47# _1030_/a_1059_315# 0
C28830 _0172_ net10 0.11306f
C28831 net175 _1048_/a_1059_315# 0.03305f
C28832 net9 _1048_/a_193_47# 0.01928f
C28833 hold25/a_391_47# _1038_/a_466_413# 0
C28834 hold25/a_49_47# _1038_/a_891_413# 0
C28835 _0517_/a_384_47# acc0.A\[10\] 0
C28836 _0958_/a_27_47# _1062_/a_634_159# 0
C28837 _0538_/a_51_297# _1045_/a_891_413# 0
C28838 _0538_/a_240_47# _1045_/a_193_47# 0
C28839 net44 _0779_/a_215_47# 0
C28840 net3 _0511_/a_81_21# 0
C28841 comp0.B\[8\] net147 0
C28842 net149 _1047_/a_634_159# 0.00736f
C28843 clkload4/Y _1017_/a_891_413# 0
C28844 hold13/a_285_47# _0473_ 0.02492f
C28845 VPWR _1022_/a_634_159# 0.18536f
C28846 pp[15] _0405_ 0
C28847 net59 _0568_/a_27_297# 0
C28848 _0504_/a_27_47# net247 0.05739f
C28849 _0284_ _0402_ 0.21611f
C28850 _0155_ acc0.A\[10\] 0.00177f
C28851 _0553_/a_240_47# _0173_ 0
C28852 _0553_/a_245_297# _0208_ 0
C28853 clknet_1_1__leaf__0459_ _0993_/a_193_47# 0.00106f
C28854 _0999_/a_27_47# _0999_/a_466_413# 0.27314f
C28855 _0999_/a_193_47# _0999_/a_634_159# 0.11897f
C28856 _0993_/a_466_413# net38 0
C28857 clknet_0__0457_ net157 0
C28858 _0460_ net51 0.00102f
C28859 _0820_/a_297_297# _0290_ 0.00202f
C28860 _0820_/a_79_21# _0401_ 0
C28861 _0992_/a_27_47# net217 0
C28862 VPWR _0771_/a_215_297# 0.18567f
C28863 _1017_/a_634_159# net221 0
C28864 net166 _0219_ 0
C28865 _0341_ _1031_/a_27_47# 0
C28866 clknet_1_0__leaf__0465_ _0989_/a_193_47# 0
C28867 clknet_1_0__leaf__0465_ hold1/a_285_47# 0.02069f
C28868 _0456_ net247 0
C28869 net120 _1034_/a_193_47# 0.00519f
C28870 hold58/a_391_47# VPWR 0.1895f
C28871 _1035_/a_891_413# net25 0.00283f
C28872 hold86/a_49_47# _0261_ 0
C28873 hold86/a_285_47# _0262_ 0
C28874 _0174_ _0472_ 0.04469f
C28875 net17 clknet_1_0__leaf__0457_ 0.21411f
C28876 _1062_/a_891_413# _1062_/a_1017_47# 0.00617f
C28877 _1062_/a_193_47# _0160_ 0.24062f
C28878 input23/a_75_212# B[2] 0.04721f
C28879 B[15] input25/a_75_212# 0
C28880 clknet_1_1__leaf__0465_ _0506_/a_299_297# 0.00121f
C28881 _1011_/a_891_413# _0353_ 0
C28882 net39 _0647_/a_129_47# 0.00343f
C28883 acc0.A\[12\] _0647_/a_377_297# 0.00203f
C28884 _0600_/a_103_199# _0345_ 0
C28885 net56 _0702_/a_113_47# 0
C28886 _1021_/a_634_159# _1021_/a_592_47# 0
C28887 _1033_/a_1059_315# net23 0
C28888 net199 _1024_/a_891_413# 0.00212f
C28889 _0257_ acc0.A\[4\] 0.00269f
C28890 _0454_ _0266_ 0
C28891 _0455_ _0452_ 0.00197f
C28892 _0467_ comp0.B\[0\] 0.16326f
C28893 _1017_/a_1059_315# _0459_ 0.00674f
C28894 _0147_ _1048_/a_891_413# 0
C28895 _1049_/a_381_47# net134 0.01806f
C28896 acc0.A\[16\] _0398_ 0.00116f
C28897 _0179_ hold82/a_49_47# 0
C28898 _0476_ _0563_/a_240_47# 0
C28899 hold14/a_285_47# _0135_ 0.00217f
C28900 _0273_ clknet_1_1__leaf__0458_ 0
C28901 _0744_/a_27_47# _0992_/a_27_47# 0
C28902 clknet_1_0__leaf__0462_ net113 0
C28903 control0.state\[0\] _0163_ 0.17657f
C28904 _0843_/a_68_297# _0350_ 0.02521f
C28905 net69 hold18/a_285_47# 0
C28906 _0996_/a_27_47# _0795_/a_81_21# 0
C28907 _0733_/a_222_93# _0733_/a_448_47# 0.00596f
C28908 _1056_/a_27_47# acc0.A\[12\] 0
C28909 _0139_ _0545_/a_68_297# 0
C28910 acc0.A\[12\] _0671_/a_113_297# 0.00396f
C28911 _0963_/a_285_297# clk 0
C28912 hold65/a_391_47# _0274_ 0
C28913 _0682_/a_68_297# _0682_/a_150_297# 0.00477f
C28914 net62 _0988_/a_466_413# 0.004f
C28915 _0181_ _0583_/a_373_47# 0
C28916 _0556_/a_150_297# VPWR 0.00126f
C28917 _0252_ clkbuf_1_0__f__0465_/a_110_47# 0
C28918 hold11/a_49_47# VPWR 0.2817f
C28919 net48 _1022_/a_634_159# 0
C28920 net54 _1026_/a_634_159# 0
C28921 _1031_/a_466_413# _1013_/a_634_159# 0
C28922 _1031_/a_193_47# _1013_/a_1059_315# 0
C28923 net125 comp0.B\[8\] 0
C28924 _0216_ _0568_/a_109_47# 0.00111f
C28925 _0372_ _0242_ 0
C28926 net132 _1061_/a_466_413# 0
C28927 _1046_/a_466_413# net147 0
C28928 hold57/a_285_47# VPWR 0.27372f
C28929 _0953_/a_220_297# comp0.B\[8\] 0.01292f
C28930 _0953_/a_114_297# _0206_ 0
C28931 _0817_/a_81_21# _0426_ 0.11199f
C28932 VPWR _0302_ 0.70728f
C28933 VPWR _0978_/a_109_297# 0.19671f
C28934 _1034_/a_891_413# clknet_0__0463_ 0.00179f
C28935 VPWR _0795_/a_299_297# 0.28749f
C28936 _0742_/a_81_21# clknet_0__0460_ 0
C28937 hold97/a_285_47# net54 0.02372f
C28938 hold19/a_49_47# _1017_/a_193_47# 0
C28939 hold19/a_285_47# _1017_/a_27_47# 0
C28940 hold85/a_49_47# hold85/a_391_47# 0.00188f
C28941 _0780_/a_35_297# _0780_/a_285_297# 0.02504f
C28942 clknet_1_0__leaf__0465_ _0538_/a_245_297# 0
C28943 hold78/a_285_47# _0111_ 0.00236f
C28944 net106 clknet_1_0__leaf__0460_ 0
C28945 _1055_/a_27_47# _0189_ 0
C28946 _0352_ hold94/a_285_47# 0
C28947 _0561_/a_240_47# _0208_ 0.05745f
C28948 _0213_ _0173_ 0.54217f
C28949 _0561_/a_512_297# _0132_ 0.00138f
C28950 VPWR _1067_/a_1059_315# 0.41466f
C28951 _1050_/a_634_159# _0186_ 0.00931f
C28952 acc0.A\[14\] _0261_ 0.27402f
C28953 hold28/a_49_47# hold28/a_285_47# 0.22264f
C28954 net17 _1062_/a_466_413# 0
C28955 hold99/a_49_47# net38 0.34052f
C28956 _1033_/a_634_159# clknet_1_0__leaf__0461_ 0
C28957 _0717_/a_80_21# VPWR 0.1832f
C28958 _0228_ _1005_/a_466_413# 0.00311f
C28959 _0635_/a_27_47# _0446_ 0.04236f
C28960 VPWR B[10] 0.29663f
C28961 acc0.A\[21\] clknet_1_0__leaf__0457_ 0.00274f
C28962 _1019_/a_27_47# _0869_/a_27_47# 0
C28963 _0359_ _1007_/a_27_47# 0
C28964 _0237_ clknet_1_0__leaf__0460_ 0.0226f
C28965 _1020_/a_381_47# net106 0
C28966 _0179_ net4 0.09085f
C28967 _0472_ _0208_ 0.00887f
C28968 _0346_ _0085_ 0.01665f
C28969 VPWR _0339_ 0.83715f
C28970 _0243_ _0771_/a_298_297# 0.05314f
C28971 _0390_ _0771_/a_215_297# 0.00651f
C28972 _0348_ _1030_/a_891_413# 0
C28973 _0229_ acc0.A\[20\] 0
C28974 net215 _0222_ 0
C28975 _0746_/a_299_297# _0370_ 0.09703f
C28976 _0458_ _0640_/a_109_53# 0
C28977 comp0.B\[15\] _0563_/a_149_47# 0
C28978 net47 _0158_ 0
C28979 _1047_/a_891_413# _0145_ 0.00251f
C28980 net45 _0790_/a_285_297# 0
C28981 _1000_/a_27_47# acc0.A\[19\] 0
C28982 _1003_/a_891_413# _0760_/a_47_47# 0
C28983 _0305_ _0397_ 0.0074f
C28984 net83 _0095_ 0.08279f
C28985 clknet_1_0__leaf_clk _0485_ 0.00458f
C28986 _0212_ _0173_ 0.21245f
C28987 clknet_1_1__leaf__0460_ _0319_ 0.02028f
C28988 hold46/a_49_47# comp0.B\[10\] 0
C28989 _0082_ _0345_ 0
C28990 _0343_ _0305_ 0.03993f
C28991 _0343_ _0349_ 0
C28992 _0546_/a_51_297# _1040_/a_27_47# 0
C28993 _0456_ net100 0
C28994 net188 _0188_ 0.65041f
C28995 _0953_/a_32_297# _1046_/a_891_413# 0
C28996 _0183_ _1018_/a_592_47# 0
C28997 _0567_/a_109_297# acc0.A\[30\] 0.00152f
C28998 clknet_1_0__leaf__0461_ net223 0
C28999 _0369_ pp[4] 0
C29000 clkbuf_1_1__f__0462_/a_110_47# _0701_/a_80_21# 0.00791f
C29001 _0513_/a_81_21# net4 0.02249f
C29002 _0200_ _0473_ 0.23569f
C29003 _0305_ net95 0.00343f
C29004 output44/a_27_47# hold15/a_391_47# 0
C29005 _0101_ hold3/a_49_47# 0.0036f
C29006 _0518_/a_109_47# _0186_ 0.00371f
C29007 _0712_/a_79_21# _0341_ 0
C29008 _0994_/a_193_47# net246 0
C29009 net36 _0176_ 0.13937f
C29010 net224 acc0.A\[27\] 0
C29011 VPWR _0159_ 0.33867f
C29012 _0387_ _0308_ 0.44167f
C29013 _0544_/a_51_297# _0544_/a_512_297# 0.0116f
C29014 net58 _0458_ 0.00797f
C29015 _0956_/a_114_297# control0.reset 0.00171f
C29016 _0375_ net213 0
C29017 _0473_ comp0.B\[8\] 0.0338f
C29018 acc0.A\[4\] net11 0.01794f
C29019 _1034_/a_27_47# _1034_/a_1059_315# 0.04875f
C29020 _1034_/a_193_47# _1034_/a_466_413# 0.08301f
C29021 _0536_/a_51_297# _0536_/a_149_47# 0.02487f
C29022 _0796_/a_215_47# _0796_/a_510_47# 0.00529f
C29023 _1021_/a_193_47# acc0.A\[21\] 0
C29024 net168 _1053_/a_466_413# 0
C29025 net14 _1053_/a_27_47# 0
C29026 acc0.A\[1\] _0219_ 0
C29027 net205 _0175_ 0.06209f
C29028 VPWR net6 3.2056f
C29029 _0218_ _0115_ 0
C29030 _0430_ _0826_/a_27_53# 0.00665f
C29031 comp0.B\[1\] control0.reset 0.012f
C29032 _1057_/a_592_47# net67 0
C29033 _0982_/a_891_413# clknet_1_0__leaf__0461_ 0
C29034 net117 _0219_ 0.03467f
C29035 _0350_ acc0.A\[23\] 0.61408f
C29036 _0850_/a_68_297# _0446_ 0
C29037 _0217_ _0855_/a_299_297# 0.0092f
C29038 net86 _0372_ 0
C29039 _0516_/a_109_297# acc0.A\[9\] 0.00807f
C29040 hold36/a_285_47# _0954_/a_32_297# 0
C29041 control0.state\[0\] _1066_/a_27_47# 0.0028f
C29042 _0570_/a_27_297# _0570_/a_109_297# 0.17136f
C29043 acc0.A\[12\] _0802_/a_59_75# 0
C29044 net39 _0802_/a_145_75# 0
C29045 clkbuf_0__0464_/a_110_47# _1045_/a_634_159# 0
C29046 clkbuf_0__0463_/a_110_47# _0563_/a_240_47# 0
C29047 _0963_/a_35_297# hold79/a_49_47# 0
C29048 _0598_/a_79_21# _0460_ 0
C29049 _1063_/a_1059_315# _0161_ 0.06159f
C29050 _0225_ _0756_/a_47_47# 0.07209f
C29051 net235 _0988_/a_634_159# 0
C29052 _0746_/a_384_47# _0350_ 0.00127f
C29053 VPWR _0447_ 0.50148f
C29054 _0965_/a_47_47# _0169_ 0
C29055 control0.state\[0\] _1068_/a_27_47# 0
C29056 VPWR _1026_/a_193_47# 0.30959f
C29057 _0854_/a_215_47# acc0.A\[18\] 0
C29058 hold68/a_285_47# _0216_ 0
C29059 control0.count\[3\] _1072_/a_634_159# 0.01605f
C29060 _0483_ _1072_/a_27_47# 0
C29061 _0666_/a_113_47# VPWR 0
C29062 hold88/a_285_47# clknet_1_1__leaf__0458_ 0.01604f
C29063 _0712_/a_79_21# _1013_/a_891_413# 0
C29064 _0712_/a_297_297# _1013_/a_1059_315# 0
C29065 net78 _0992_/a_634_159# 0
C29066 _0547_/a_68_297# _0547_/a_150_297# 0.00477f
C29067 acc0.A\[14\] net47 0.02482f
C29068 _0793_/a_51_297# _0790_/a_35_297# 0.00163f
C29069 net159 _0161_ 0
C29070 VPWR _1024_/a_891_413# 0.19738f
C29071 _0959_/a_472_297# _0470_ 0.00397f
C29072 _0399_ hold91/a_49_47# 0.03102f
C29073 hold13/a_49_47# hold13/a_391_47# 0.00188f
C29074 output42/a_27_47# _1013_/a_27_47# 0
C29075 net203 _0563_/a_149_47# 0.00896f
C29076 _0585_/a_109_47# net149 0
C29077 _0172_ _0498_/a_245_297# 0
C29078 _0517_/a_81_21# _0517_/a_299_297# 0.08213f
C29079 hold97/a_49_47# VPWR 0.32069f
C29080 net62 _0186_ 0.02453f
C29081 _0956_/a_304_297# net24 0
C29082 VPWR _1048_/a_561_413# 0.00338f
C29083 comp0.B\[14\] comp0.B\[10\] 0
C29084 clknet_1_0__leaf__0460_ _1005_/a_27_47# 0.00361f
C29085 acc0.A\[4\] hold7/a_391_47# 0.00192f
C29086 net234 _0580_/a_27_297# 0.01107f
C29087 _0731_/a_384_47# _0312_ 0
C29088 hold85/a_49_47# _0160_ 0.0015f
C29089 _1017_/a_27_47# _1017_/a_634_159# 0.13601f
C29090 output45/a_27_47# pp[31] 0.02112f
C29091 _1058_/a_27_47# _0512_/a_27_297# 0
C29092 net193 _0473_ 0.00204f
C29093 _0461_ _0721_/a_27_47# 0.20427f
C29094 _0753_/a_79_21# _0752_/a_27_413# 0
C29095 _0601_/a_68_297# _0232_ 0
C29096 pp[27] _0725_/a_209_47# 0
C29097 _0211_ control0.sh 0.01734f
C29098 _0428_ clknet_0__0465_ 0.50379f
C29099 clknet_1_1__leaf__0462_ hold62/a_285_47# 0
C29100 _0472_ _1046_/a_193_47# 0
C29101 _0473_ _1046_/a_466_413# 0.00297f
C29102 _0984_/a_193_47# _0345_ 0
C29103 _0457_ _0178_ 0
C29104 _0343_ _0675_/a_150_297# 0
C29105 _0195_ acc0.A\[29\] 0.62379f
C29106 _0086_ clknet_1_1__leaf__0458_ 0.15873f
C29107 net46 _0580_/a_27_297# 0
C29108 hold101/a_285_47# _0255_ 0
C29109 _0660_/a_113_47# clknet_0__0465_ 0
C29110 net194 hold49/a_285_47# 0
C29111 _1004_/a_1059_315# net110 0.00113f
C29112 _1004_/a_27_47# acc0.A\[24\] 0
C29113 _1000_/a_634_159# _1000_/a_592_47# 0
C29114 _0600_/a_253_297# clknet_1_0__leaf__0460_ 0
C29115 _1060_/a_891_413# net146 0
C29116 _1060_/a_1059_315# _0158_ 0
C29117 _0188_ _0155_ 0.12868f
C29118 _0993_/a_634_159# _0281_ 0
C29119 _1051_/a_381_47# net154 0
C29120 net114 net94 0
C29121 _0256_ net72 0
C29122 control0.count\[1\] _0979_/a_109_47# 0
C29123 hold43/a_285_47# acc0.A\[28\] 0.08268f
C29124 VPWR _0480_ 0.82363f
C29125 _0346_ _0815_/a_113_297# 0.03285f
C29126 _0671_/a_113_297# net42 0.048f
C29127 _0459_ _0508_/a_384_47# 0
C29128 _0305_ _0998_/a_193_47# 0
C29129 _0192_ net14 0.00299f
C29130 _0151_ net168 0.02467f
C29131 _0462_ _0240_ 0.00278f
C29132 _1072_/a_27_47# control0.count\[1\] 0
C29133 _1072_/a_891_413# VPWR 0.17766f
C29134 hold55/a_285_47# clknet_1_0__leaf__0457_ 0.00585f
C29135 _0251_ clkbuf_1_1__f__0458_/a_110_47# 0.00384f
C29136 clkbuf_0__0463_/a_110_47# _0935_/a_27_47# 0
C29137 _0277_ hold91/a_285_47# 0
C29138 clkbuf_0__0463_/a_110_47# _1061_/a_193_47# 0
C29139 _0462_ _0369_ 0.03913f
C29140 _0786_/a_80_21# net228 0.0184f
C29141 clkbuf_1_1__f__0463_/a_110_47# _0493_/a_27_47# 0
C29142 _0554_/a_150_297# VPWR 0.00129f
C29143 clknet_0__0458_ _0842_/a_145_75# 0
C29144 acc0.A\[17\] _0675_/a_68_297# 0.06934f
C29145 hold56/a_391_47# control0.reset 0.00436f
C29146 _0350_ hold60/a_49_47# 0
C29147 _0625_/a_59_75# _0218_ 0.00249f
C29148 _0684_/a_59_75# _0734_/a_47_47# 0.00108f
C29149 _0399_ _0986_/a_1017_47# 0
C29150 comp0.B\[10\] _0543_/a_68_297# 0.00801f
C29151 _0763_/a_109_47# _0345_ 0
C29152 _0289_ _0817_/a_81_21# 0.00106f
C29153 net240 _1063_/a_634_159# 0
C29154 net56 net97 0
C29155 _0346_ _0849_/a_297_297# 0
C29156 _0457_ _1033_/a_381_47# 0
C29157 _0736_/a_56_297# _1009_/a_634_159# 0
C29158 _0343_ _0618_/a_297_297# 0.00441f
C29159 clkbuf_1_0__f__0457_/a_110_47# _0579_/a_27_297# 0
C29160 _0283_ _0302_ 0.0014f
C29161 _0583_/a_109_297# _0114_ 0.00277f
C29162 clknet_1_0__leaf__0458_ net36 0.00247f
C29163 VPWR acc0.A\[0\] 0.59363f
C29164 _0165_ clknet_1_0__leaf__0457_ 0.04973f
C29165 _0750_/a_27_47# _0750_/a_109_47# 0.00517f
C29166 _1072_/a_193_47# clkbuf_1_0__f_clk/a_110_47# 0.0011f
C29167 _1050_/a_27_47# _1050_/a_1059_315# 0.04875f
C29168 _1050_/a_193_47# _1050_/a_466_413# 0.08015f
C29169 _0476_ _1035_/a_1059_315# 0
C29170 _1019_/a_634_159# clknet_1_0__leaf__0457_ 0
C29171 _0557_/a_245_297# comp0.B\[5\] 0
C29172 _0985_/a_1017_47# _0179_ 0.0016f
C29173 hold50/a_49_47# hold50/a_285_47# 0.22264f
C29174 clkbuf_0__0458_/a_110_47# _0345_ 0.02853f
C29175 _0432_ _0826_/a_219_297# 0
C29176 hold85/a_391_47# net17 0.05325f
C29177 net224 _1010_/a_193_47# 0
C29178 _0294_ _0775_/a_79_21# 0.00628f
C29179 _0221_ _1011_/a_466_413# 0.03689f
C29180 hold21/a_49_47# acc0.A\[7\] 0.33279f
C29181 _0715_/a_27_47# clknet_0__0465_ 0
C29182 clknet_1_1__leaf__0460_ _0780_/a_285_297# 0
C29183 clknet_1_1__leaf__0463_ _1065_/a_891_413# 0.00558f
C29184 _0397_ _0181_ 0
C29185 net58 clkbuf_1_1__f__0458_/a_110_47# 0.01864f
C29186 _0838_/a_109_297# _0441_ 0
C29187 _0179_ _1049_/a_561_413# 0.00156f
C29188 _1051_/a_1059_315# hold7/a_285_47# 0
C29189 _0464_ _0198_ 0
C29190 _0337_ output44/a_27_47# 0
C29191 _0181_ _1049_/a_466_413# 0
C29192 _0778_/a_150_297# _0352_ 0
C29193 net54 _0689_/a_68_297# 0
C29194 _0999_/a_466_413# _1012_/a_634_159# 0
C29195 _0999_/a_634_159# _1012_/a_466_413# 0
C29196 _0499_/a_145_75# _0208_ 0
C29197 _0343_ _0181_ 0.23929f
C29198 B[4] B[0] 0
C29199 _0458_ _0262_ 0.0079f
C29200 net157 _0138_ 0
C29201 _0161_ _0173_ 0
C29202 _0718_/a_47_47# VPWR 0.31945f
C29203 _0997_/a_561_413# net41 0.00197f
C29204 _0997_/a_891_413# pp[14] 0
C29205 _0998_/a_27_47# net43 0.01389f
C29206 clknet_0__0464_ _1046_/a_1017_47# 0
C29207 _0324_ _0460_ 0.01343f
C29208 _1054_/a_193_47# _1052_/a_27_47# 0
C29209 _1054_/a_27_47# _1052_/a_193_47# 0.00785f
C29210 acc0.A\[4\] clknet_1_1__leaf__0458_ 0.07937f
C29211 hold74/a_285_47# clkload3/Y 0
C29212 net94 _0365_ 0.09508f
C29213 _0302_ _0794_/a_110_297# 0
C29214 hold33/a_285_47# VPWR 0.26788f
C29215 clknet_1_1__leaf__0459_ _0788_/a_68_297# 0.01346f
C29216 net224 _1009_/a_634_159# 0
C29217 _0249_ _0374_ 0.00425f
C29218 _0795_/a_81_21# _0794_/a_27_47# 0
C29219 net149 _0208_ 0
C29220 net95 _0181_ 0.02077f
C29221 acc0.A\[5\] _0087_ 0
C29222 _1039_/a_193_47# clkbuf_0__0463_/a_110_47# 0.00207f
C29223 _0538_/a_149_47# _1044_/a_193_47# 0
C29224 _0538_/a_240_47# _1044_/a_27_47# 0
C29225 comp0.B\[11\] _1043_/a_1017_47# 0
C29226 hold25/a_391_47# net172 0.1316f
C29227 acc0.A\[14\] _1060_/a_1059_315# 0.09726f
C29228 clknet_1_0__leaf__0464_ _0144_ 0.01329f
C29229 _0477_ _1062_/a_634_159# 0
C29230 hold65/a_49_47# hold65/a_285_47# 0.22264f
C29231 pp[28] _0725_/a_209_297# 0.00117f
C29232 hold46/a_285_47# hold46/a_391_47# 0.41909f
C29233 _1000_/a_466_413# _1018_/a_891_413# 0
C29234 _1000_/a_891_413# _1018_/a_466_413# 0
C29235 output56/a_27_47# _0353_ 0
C29236 net25 _0561_/a_512_297# 0
C29237 control0.state\[2\] _1068_/a_891_413# 0.00378f
C29238 _0486_ _1068_/a_1059_315# 0.05237f
C29239 hold27/a_285_47# net174 0.00926f
C29240 _0143_ _1045_/a_466_413# 0
C29241 hold58/a_391_47# _1036_/a_27_47# 0
C29242 hold58/a_285_47# _1036_/a_193_47# 0
C29243 _0606_/a_297_297# _0460_ 0
C29244 _0973_/a_27_297# _0973_/a_109_47# 0.00393f
C29245 net175 clkbuf_1_1__f__0457_/a_110_47# 0
C29246 _0946_/a_30_53# clk 0.0061f
C29247 _0172_ _0492_/a_27_47# 0.15496f
C29248 _0343_ _1000_/a_466_413# 0.00817f
C29249 _1033_/a_466_413# _0173_ 0
C29250 _1033_/a_27_47# _0208_ 0
C29251 _0328_ _0371_ 0
C29252 _0217_ _1015_/a_27_47# 0
C29253 _0268_ _0465_ 0.03015f
C29254 _0999_/a_193_47# net85 0.00539f
C29255 _0999_/a_1059_315# _0999_/a_1017_47# 0
C29256 _0454_ _0399_ 0.24858f
C29257 net17 _1063_/a_1017_47# 0.0018f
C29258 _0339_ _0567_/a_373_47# 0
C29259 _1001_/a_381_47# _1019_/a_27_47# 0.00111f
C29260 _1001_/a_193_47# _1019_/a_891_413# 0
C29261 _1001_/a_634_159# _1019_/a_1059_315# 0.00319f
C29262 _0487_ clknet_1_0__leaf__0461_ 0
C29263 _0472_ comp0.B\[9\] 0.00894f
C29264 net103 net221 0.02208f
C29265 clknet_1_0__leaf__0459_ net6 0
C29266 VPWR _0993_/a_891_413# 0.204f
C29267 _1001_/a_1017_47# net223 0
C29268 _1054_/a_27_47# net12 0
C29269 _1054_/a_466_413# net148 0
C29270 net204 _0957_/a_32_297# 0
C29271 net77 _0219_ 0
C29272 net67 _0345_ 0.05015f
C29273 _0663_/a_207_413# _0346_ 0.03807f
C29274 hold68/a_391_47# _1024_/a_27_47# 0
C29275 _0814_/a_27_47# net67 0
C29276 _0298_ hold91/a_285_47# 0
C29277 clknet_1_0__leaf__0462_ _1007_/a_891_413# 0.00653f
C29278 _1041_/a_381_47# hold5/a_391_47# 0
C29279 _0697_/a_217_297# _0321_ 0
C29280 VPWR _0580_/a_109_297# 0.17641f
C29281 _0983_/a_193_47# _0183_ 0
C29282 _0983_/a_466_413# _0217_ 0
C29283 hold88/a_391_47# net47 0.00876f
C29284 _0775_/a_79_21# _0775_/a_297_297# 0.01735f
C29285 _0186_ _0987_/a_634_159# 0
C29286 hold74/a_49_47# net45 0.00353f
C29287 _1043_/a_193_47# _0542_/a_149_47# 0
C29288 _1043_/a_27_47# _0542_/a_240_47# 0
C29289 _0556_/a_68_297# _1036_/a_193_47# 0
C29290 _0223_ _0219_ 0.03003f
C29291 _0642_/a_27_413# pp[3] 0
C29292 B[9] _0204_ 0
C29293 hold24/a_285_47# net172 0
C29294 _1001_/a_193_47# net206 0
C29295 net185 input25/a_75_212# 0
C29296 acc0.A\[3\] net134 0
C29297 hold34/a_285_47# acc0.A\[11\] 0
C29298 _1016_/a_27_47# _0459_ 0.00213f
C29299 _0648_/a_27_297# _0278_ 0.18564f
C29300 clknet_1_1__leaf__0459_ _0406_ 0
C29301 _0999_/a_1059_315# clknet_1_1__leaf__0461_ 0
C29302 pp[8] _0512_/a_27_297# 0.00116f
C29303 net14 A[5] 0
C29304 VPWR net20 0.45073f
C29305 hold17/a_49_47# net164 0
C29306 hold17/a_285_47# _0480_ 0
C29307 control0.count\[2\] _0979_/a_373_47# 0
C29308 _0547_/a_68_297# net153 0
C29309 _0996_/a_1059_315# _0409_ 0
C29310 _1017_/a_891_413# _0218_ 0
C29311 hold48/a_285_47# VPWR 0.35795f
C29312 _0258_ clknet_0__0465_ 0.04034f
C29313 _0237_ hold94/a_285_47# 0
C29314 VPWR _0790_/a_285_297# 0.26109f
C29315 _0249_ acc0.A\[19\] 0
C29316 _0691_/a_150_297# clknet_0__0460_ 0
C29317 net97 _0345_ 0.18874f
C29318 _1002_/a_634_159# clknet_1_0__leaf__0460_ 0
C29319 _0294_ _0158_ 0.01884f
C29320 _1006_/a_1059_315# _0219_ 0
C29321 hold41/a_391_47# acc0.A\[11\] 0.04239f
C29322 clknet_1_1__leaf__0460_ _0333_ 0
C29323 _0467_ net1 0.02987f
C29324 net160 _0175_ 0.11162f
C29325 hold83/a_49_47# hold83/a_391_47# 0.00188f
C29326 _0985_/a_27_47# _0985_/a_561_413# 0.0027f
C29327 _0985_/a_634_159# _0985_/a_891_413# 0.03684f
C29328 _0985_/a_193_47# _0985_/a_381_47# 0.09799f
C29329 _0304_ acc0.A\[9\] 0
C29330 _0183_ _0526_/a_27_47# 0
C29331 hold39/a_49_47# comp0.B\[3\] 0
C29332 _0217_ hold29/a_285_47# 0
C29333 acc0.A\[22\] hold29/a_49_47# 0.28964f
C29334 hold38/a_285_47# comp0.B\[2\] 0
C29335 _0325_ _1007_/a_27_47# 0
C29336 _0973_/a_109_47# net17 0
C29337 _0464_ clknet_1_1__leaf__0464_ 0.01887f
C29338 _0998_/a_193_47# _0181_ 0
C29339 _1018_/a_634_159# _1018_/a_466_413# 0.23992f
C29340 _1018_/a_193_47# _1018_/a_1059_315# 0.03405f
C29341 _1018_/a_27_47# _1018_/a_891_413# 0.03089f
C29342 _0794_/a_110_297# net6 0.0014f
C29343 net235 _0253_ 0.00366f
C29344 control0.count\[2\] _1071_/a_1017_47# 0.00168f
C29345 _0985_/a_27_47# _1049_/a_1059_315# 0
C29346 net50 _1022_/a_1059_315# 0.0011f
C29347 _0642_/a_27_413# _0273_ 0.00383f
C29348 _0404_ _0670_/a_510_47# 0
C29349 _0399_ _0506_/a_81_21# 0
C29350 hold28/a_285_47# clkbuf_1_0__f__0464_/a_110_47# 0.0207f
C29351 _0982_/a_27_47# _0982_/a_634_159# 0.14145f
C29352 net136 _0186_ 0
C29353 _0275_ _0990_/a_1059_315# 0
C29354 net45 _0583_/a_27_297# 0
C29355 _0210_ control0.sh 0.02772f
C29356 _1049_/a_27_47# _1049_/a_193_47# 0.9692f
C29357 _0343_ _1018_/a_27_47# 0
C29358 _0725_/a_80_21# _0335_ 0
C29359 net17 _0160_ 0
C29360 _0983_/a_193_47# acc0.A\[15\] 0.00321f
C29361 clknet_1_1__leaf__0460_ _0732_/a_80_21# 0.00789f
C29362 clknet_1_1__leaf_clk _0951_/a_296_53# 0
C29363 clknet_1_1__leaf__0462_ _0350_ 0.63261f
C29364 _0228_ _0103_ 0
C29365 _0267_ _0451_ 0.03394f
C29366 _1019_/a_381_47# _0459_ 0
C29367 hold99/a_391_47# VPWR 0.19416f
C29368 net1 comp0.B\[0\] 0
C29369 _0753_/a_79_21# _0233_ 0.03271f
C29370 B[12] hold5/a_49_47# 0
C29371 _0461_ clkbuf_1_0__f__0461_/a_110_47# 0.04108f
C29372 _0530_/a_299_297# _0197_ 0.01431f
C29373 hold44/a_285_47# _0216_ 0.01441f
C29374 _0276_ _0669_/a_183_297# 0.00452f
C29375 _1054_/a_634_159# input15/a_75_212# 0
C29376 _0644_/a_129_47# _0301_ 0
C29377 _1019_/a_193_47# _0586_/a_27_47# 0
C29378 hold27/a_285_47# clknet_0__0464_ 0
C29379 VPWR _1027_/a_592_47# 0
C29380 hold98/a_49_47# hold98/a_391_47# 0.00188f
C29381 _0555_/a_512_297# _0135_ 0
C29382 hold46/a_285_47# net153 0
C29383 _0218_ net223 0.04998f
C29384 _1066_/a_27_47# _1066_/a_193_47# 0.97386f
C29385 _0473_ _1045_/a_193_47# 0
C29386 comp0.B\[7\] _0913_/a_27_47# 0
C29387 _0693_/a_68_297# _0367_ 0
C29388 net56 _1010_/a_27_47# 0.00396f
C29389 clknet_1_0__leaf__0461_ clkbuf_0__0457_/a_110_47# 0.18458f
C29390 clkbuf_1_0__f__0459_/a_110_47# _0305_ 0.01915f
C29391 net89 _0760_/a_285_47# 0
C29392 net45 _0999_/a_193_47# 0.01207f
C29393 clknet_1_1__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# 0
C29394 VPWR _1052_/a_634_159# 0.17694f
C29395 _0335_ _0128_ 0
C29396 _0330_ clkbuf_1_1__f__0462_/a_110_47# 0.01907f
C29397 _0833_/a_79_21# _0833_/a_297_297# 0.01735f
C29398 _1056_/a_891_413# acc0.A\[10\] 0.03157f
C29399 _1031_/a_27_47# acc0.A\[30\] 0.01679f
C29400 _1023_/a_193_47# _1022_/a_193_47# 0
C29401 _1023_/a_27_47# _1022_/a_634_159# 0
C29402 _0967_/a_109_93# clk 0
C29403 _1068_/a_27_47# _1068_/a_193_47# 0.96566f
C29404 net8 _1040_/a_193_47# 0
C29405 clk _0487_ 0.05857f
C29406 net157 net134 0.00312f
C29407 _0176_ _0563_/a_149_47# 0
C29408 _0174_ _1046_/a_891_413# 0.00137f
C29409 acc0.A\[25\] _1008_/a_891_413# 0
C29410 _0500_/a_27_47# VPWR 0.37936f
C29411 _1056_/a_466_413# hold67/a_49_47# 0
C29412 hold100/a_49_47# _0450_ 0
C29413 hold100/a_285_47# _0446_ 0.02508f
C29414 hold3/a_391_47# _0460_ 0
C29415 _0134_ _1036_/a_193_47# 0.00371f
C29416 _0677_/a_47_47# acc0.A\[17\] 0.05536f
C29417 clknet_1_1__leaf__0460_ _0250_ 0.05832f
C29418 net152 _1040_/a_634_159# 0
C29419 net32 _1040_/a_193_47# 0
C29420 _0205_ _1040_/a_1059_315# 0
C29421 _0487_ _1063_/a_891_413# 0
C29422 clkbuf_1_1__f__0464_/a_110_47# _1045_/a_193_47# 0
C29423 clkbuf_0__0460_/a_110_47# _0743_/a_240_47# 0
C29424 acc0.A\[14\] _0294_ 0.04103f
C29425 hold58/a_49_47# comp0.B\[5\] 0.01335f
C29426 hold58/a_391_47# comp0.B\[3\] 0.00124f
C29427 acc0.A\[8\] _0989_/a_1017_47# 0
C29428 _0231_ _0374_ 0
C29429 output57/a_27_47# _0219_ 0
C29430 _0804_/a_79_21# _0278_ 0
C29431 _1032_/a_27_47# net23 0.0291f
C29432 net36 hold18/a_49_47# 0
C29433 net44 _0676_/a_113_47# 0
C29434 _0994_/a_381_47# net80 0
C29435 _0478_ _1068_/a_27_47# 0
C29436 hold78/a_49_47# _0342_ 0
C29437 _0544_/a_51_297# _0140_ 0.10222f
C29438 _0544_/a_240_47# net198 0.04098f
C29439 _0811_/a_299_297# net37 0
C29440 net9 acc0.A\[15\] 0
C29441 VPWR _0685_/a_150_297# 0.00193f
C29442 _0358_ _0347_ 0.00409f
C29443 _0104_ _0460_ 0.04505f
C29444 _1034_/a_891_413# _1034_/a_1017_47# 0.00617f
C29445 _0557_/a_51_297# net26 0.02343f
C29446 _0110_ _0395_ 0.0032f
C29447 _0453_ acc0.A\[0\] 0
C29448 output65/a_27_47# _0989_/a_193_47# 0.00133f
C29449 _0343_ _0507_/a_373_47# 0
C29450 acc0.A\[16\] _0308_ 0
C29451 net58 _0291_ 0
C29452 hold6/a_285_47# hold6/a_391_47# 0.41909f
C29453 net68 _0782_/a_27_47# 0
C29454 _0222_ clknet_1_0__leaf__0460_ 0.0934f
C29455 _0464_ net247 0.028f
C29456 hold59/a_285_47# _0216_ 0
C29457 clkbuf_0__0464_/a_110_47# _1044_/a_193_47# 0
C29458 net242 _0350_ 0.09342f
C29459 _0200_ comp0.B\[8\] 0
C29460 hold85/a_285_47# _0477_ 0.00815f
C29461 _0389_ control0.add 0.07244f
C29462 _0789_/a_75_199# net6 0.01881f
C29463 _0570_/a_109_297# _0126_ 0.00194f
C29464 _0999_/a_193_47# _0587_/a_27_47# 0
C29465 clkbuf_0__0464_/a_110_47# net131 0.00209f
C29466 _0534_/a_81_21# _1047_/a_193_47# 0
C29467 _0534_/a_299_297# _1047_/a_27_47# 0
C29468 _0481_ hold79/a_391_47# 0.00386f
C29469 _0750_/a_27_47# _0606_/a_215_297# 0
C29470 _0176_ _1061_/a_27_47# 0
C29471 net62 _0450_ 0
C29472 _0179_ _0287_ 0.02142f
C29473 _0490_ _0468_ 0.00131f
C29474 _0129_ _0342_ 0
C29475 pp[30] net56 0
C29476 _0745_/a_109_47# _0460_ 0
C29477 _0645_/a_47_47# clkbuf_1_1__f__0459_/a_110_47# 0
C29478 hold29/a_49_47# _0379_ 0
C29479 pp[16] pp[14] 0.00649f
C29480 _1001_/a_466_413# _0352_ 0
C29481 pp[30] _1031_/a_634_159# 0.00171f
C29482 hold89/a_285_47# _0974_/a_79_199# 0
C29483 net213 VPWR 0.19487f
C29484 _0137_ net7 0
C29485 _1071_/a_891_413# _0466_ 0.003f
C29486 _1071_/a_381_47# _0488_ 0
C29487 VPWR clkbuf_1_1__f__0463_/a_110_47# 1.20818f
C29488 _0217_ _0452_ 0
C29489 _1021_/a_27_47# _0352_ 0
C29490 net81 _0995_/a_1059_315# 0
C29491 hold26/a_49_47# _0954_/a_32_297# 0
C29492 _0346_ _0264_ 0.73702f
C29493 net234 _0117_ 0
C29494 _0476_ _1062_/a_193_47# 0
C29495 _1017_/a_891_413# _1017_/a_975_413# 0.00851f
C29496 _1017_/a_27_47# net103 0.30144f
C29497 _1017_/a_381_47# _1017_/a_561_413# 0.00123f
C29498 _1058_/a_634_159# net3 0
C29499 _0753_/a_561_47# _0375_ 0.00217f
C29500 _0429_ _0621_/a_35_297# 0
C29501 _0430_ _0640_/a_215_297# 0
C29502 clknet_1_1__leaf__0463_ hold93/a_285_47# 0
C29503 _0786_/a_80_21# _0090_ 0
C29504 _0786_/a_472_297# _0422_ 0
C29505 comp0.B\[7\] _0172_ 0
C29506 net103 _1060_/a_975_413# 0
C29507 net127 net153 0.00644f
C29508 net10 _1040_/a_193_47# 0
C29509 _0179_ net9 0.98577f
C29510 _0126_ hold50/a_285_47# 0.00136f
C29511 _0831_/a_285_297# clkbuf_1_1__f__0458_/a_110_47# 0.00188f
C29512 _1006_/a_975_413# net52 0
C29513 _0507_/a_27_297# _0185_ 0.11141f
C29514 _0507_/a_109_47# net5 0.00301f
C29515 _1000_/a_891_413# net45 0.03707f
C29516 acc0.A\[5\] net154 0
C29517 _0149_ net11 0
C29518 net193 _0200_ 0.1998f
C29519 _0514_/a_109_297# _0186_ 0.01236f
C29520 _0804_/a_215_47# _0415_ 0.04718f
C29521 _0804_/a_297_297# _0416_ 0.00156f
C29522 clknet_1_1__leaf__0463_ _0214_ 0
C29523 _1010_/a_27_47# _0345_ 0
C29524 _0397_ clknet_1_1__leaf__0461_ 0.03519f
C29525 _0555_/a_51_297# _0136_ 0
C29526 net204 _0553_/a_240_47# 0
C29527 _0704_/a_68_297# _0219_ 0.00216f
C29528 _0211_ net172 0
C29529 _0476_ _0561_/a_245_297# 0.00308f
C29530 _1033_/a_193_47# _1033_/a_381_47# 0.10164f
C29531 _1033_/a_634_159# _1033_/a_891_413# 0.03684f
C29532 _1033_/a_27_47# _1033_/a_561_413# 0.00163f
C29533 _0373_ net51 0.00156f
C29534 pp[27] _0219_ 0.14249f
C29535 hold36/a_49_47# _0142_ 0
C29536 net14 clknet_1_0__leaf__0465_ 0.63207f
C29537 _0233_ clkbuf_1_0__f__0460_/a_110_47# 0
C29538 VPWR _0951_/a_368_53# 0
C29539 _0430_ _0465_ 0
C29540 VPWR A[8] 0.29324f
C29541 _1012_/a_193_47# _1012_/a_381_47# 0.0982f
C29542 _1012_/a_634_159# _1012_/a_891_413# 0.03684f
C29543 _1012_/a_27_47# _1012_/a_561_413# 0.0027f
C29544 _1039_/a_27_47# _0176_ 0.03831f
C29545 _0343_ clknet_1_1__leaf__0461_ 0.05959f
C29546 hold55/a_49_47# _1033_/a_27_47# 0
C29547 _0995_/a_634_159# net6 0
C29548 _0693_/a_68_297# _0742_/a_299_297# 0
C29549 net243 net215 0
C29550 _0629_/a_59_75# _0264_ 0
C29551 _0758_/a_215_47# _0105_ 0
C29552 _0512_/a_109_47# _0186_ 0.00291f
C29553 output47/a_27_47# A[9] 0
C29554 _0285_ _0807_/a_68_297# 0
C29555 _0107_ _1009_/a_466_413# 0.00302f
C29556 net213 net48 0.02339f
C29557 _0457_ comp0.B\[1\] 0.01178f
C29558 _0216_ _1031_/a_381_47# 0
C29559 _0233_ _0250_ 0.00223f
C29560 _0231_ _0249_ 0.00196f
C29561 pp[27] _0728_/a_59_75# 0.00121f
C29562 net66 clknet_1_1__leaf__0458_ 0.00234f
C29563 net173 _0545_/a_68_297# 0.01656f
C29564 _0642_/a_27_413# _0086_ 0
C29565 _1002_/a_193_47# hold93/a_49_47# 0
C29566 _0280_ net238 0
C29567 _1002_/a_27_47# hold93/a_285_47# 0.00104f
C29568 hold86/a_49_47# hold86/a_285_47# 0.22264f
C29569 VPWR _0738_/a_150_297# 0.00121f
C29570 net8 _0214_ 0
C29571 _0218_ _0798_/a_113_297# 0
C29572 _1072_/a_592_47# clknet_0_clk 0.00142f
C29573 _1050_/a_891_413# _1050_/a_1017_47# 0.00617f
C29574 _0275_ VPWR 0.90972f
C29575 net105 clknet_1_0__leaf__0457_ 0
C29576 _0343_ _1030_/a_193_47# 0.02983f
C29577 hold31/a_285_47# _0399_ 0
C29578 net36 _0455_ 0
C29579 hold26/a_285_47# _0540_/a_51_297# 0
C29580 _1024_/a_561_413# net50 0
C29581 _0958_/a_27_47# _0477_ 0.0867f
C29582 net214 acc0.A\[9\] 0.013f
C29583 clkbuf_1_0__f__0459_/a_110_47# _0181_ 0.04289f
C29584 net176 net110 0.1294f
C29585 hold26/a_49_47# net173 0
C29586 _0764_/a_384_47# _0462_ 0
C29587 VPWR _0837_/a_585_47# 0
C29588 _0465_ net222 0.0025f
C29589 _0458_ hold28/a_49_47# 0
C29590 _0565_/a_245_297# net201 0.00147f
C29591 _0181_ _0147_ 0
C29592 _0402_ _0347_ 0
C29593 hold74/a_49_47# VPWR 0.27552f
C29594 control0.state\[0\] _0965_/a_285_47# 0
C29595 _0517_/a_81_21# _0990_/a_1059_315# 0
C29596 _0311_ VPWR 0.59425f
C29597 net221 _0774_/a_68_297# 0
C29598 _0369_ _0830_/a_297_297# 0.00331f
C29599 _0312_ _0369_ 0
C29600 _1017_/a_193_47# net219 0
C29601 acc0.A\[27\] _0329_ 0.01745f
C29602 _0409_ _0297_ 0.02779f
C29603 _0715_/a_27_47# _0986_/a_27_47# 0
C29604 _0179_ _1054_/a_891_413# 0.07091f
C29605 _0305_ clkbuf_0__0461_/a_110_47# 0.00126f
C29606 net21 _1044_/a_891_413# 0
C29607 net83 _0219_ 0.01098f
C29608 _0180_ control0.reset 0.14749f
C29609 clknet_0__0465_ net72 0.00322f
C29610 net56 _0339_ 0.00251f
C29611 _0349_ _0568_/a_27_297# 0
C29612 _0118_ net187 0.2883f
C29613 _0241_ net219 0
C29614 net25 _0132_ 0.24511f
C29615 _0357_ hold95/a_285_47# 0
C29616 pp[30] _0345_ 0.07529f
C29617 _0143_ net184 0
C29618 _1031_/a_634_159# _0339_ 0.00639f
C29619 _1020_/a_193_47# clknet_0__0457_ 0
C29620 _1020_/a_1059_315# clkbuf_1_0__f__0457_/a_110_47# 0
C29621 _0997_/a_1059_315# _1013_/a_27_47# 0
C29622 _1024_/a_27_47# _1023_/a_891_413# 0
C29623 _1024_/a_193_47# _1023_/a_1059_315# 0
C29624 _0820_/a_215_47# _0369_ 0.09823f
C29625 clkbuf_1_1__f__0464_/a_110_47# net73 0
C29626 comp0.B\[13\] _1046_/a_891_413# 0.00123f
C29627 net193 _1046_/a_466_413# 0
C29628 _0781_/a_68_297# _0219_ 0
C29629 _0182_ _0465_ 0.05837f
C29630 clknet_1_1__leaf__0458_ _0350_ 0.18594f
C29631 _0424_ clknet_1_1__leaf__0465_ 0
C29632 _0131_ _0173_ 0.0505f
C29633 _1054_/a_1059_315# net75 0.0029f
C29634 net8 _1061_/a_1059_315# 0
C29635 _0343_ _0098_ 0
C29636 _0445_ _0840_/a_150_297# 0
C29637 _0443_ _0640_/a_215_297# 0.06566f
C29638 _1012_/a_1059_315# net98 0
C29639 _1012_/a_381_47# clknet_1_1__leaf__0461_ 0
C29640 _1046_/a_634_159# _1046_/a_1059_315# 0
C29641 _1046_/a_27_47# _1046_/a_381_47# 0.05761f
C29642 _1046_/a_193_47# _1046_/a_891_413# 0.19302f
C29643 VPWR _0604_/a_113_47# 0
C29644 pp[30] _0712_/a_381_47# 0
C29645 _0978_/a_373_47# _0466_ 0
C29646 _0991_/a_27_47# _0263_ 0.00164f
C29647 _0996_/a_27_47# net43 0
C29648 clknet_1_0__leaf__0463_ control0.sh 0
C29649 _1019_/a_1059_315# _0772_/a_215_47# 0
C29650 _0412_ _0409_ 0
C29651 net122 B[1] 0
C29652 net223 _0099_ 0
C29653 net8 _0207_ 0.02403f
C29654 net58 acc0.A\[1\] 0.00213f
C29655 acc0.A\[2\] _0182_ 0.04812f
C29656 _1016_/a_1059_315# _0115_ 0
C29657 net166 _0582_/a_109_297# 0
C29658 _1032_/a_1059_315# clknet_1_0__leaf__0457_ 0.00293f
C29659 _0221_ _0707_/a_544_297# 0.00575f
C29660 _0107_ _0310_ 0
C29661 hold68/a_49_47# net110 0.00898f
C29662 _1051_/a_193_47# _1050_/a_27_47# 0.00266f
C29663 _1051_/a_27_47# _1050_/a_193_47# 0.00266f
C29664 net86 acc0.A\[17\] 0
C29665 _0329_ _0364_ 0
C29666 _0163_ clkbuf_1_1__f_clk/a_110_47# 0.01818f
C29667 _0477_ _0132_ 0
C29668 comp0.B\[1\] _0475_ 0.00756f
C29669 _0207_ net32 0
C29670 VPWR _0583_/a_27_297# 0.29369f
C29671 _0985_/a_27_47# net175 0.00107f
C29672 clknet_0__0462_ _0352_ 0
C29673 _0186_ net73 0.00748f
C29674 _0996_/a_891_413# acc0.A\[15\] 0.01322f
C29675 clknet_1_0__leaf__0463_ _1038_/a_466_413# 0.00567f
C29676 hold64/a_391_47# acc0.A\[18\] 0
C29677 hold33/a_391_47# net180 0.15627f
C29678 net196 _0542_/a_245_297# 0.00122f
C29679 _1043_/a_381_47# net195 0.00199f
C29680 _1043_/a_891_413# net19 0
C29681 hold33/a_49_47# _0172_ 0.03879f
C29682 _0211_ _1036_/a_891_413# 0
C29683 acc0.A\[12\] hold42/a_391_47# 0
C29684 _0443_ _0465_ 0.03452f
C29685 hold38/a_391_47# _0215_ 0
C29686 _0399_ _0184_ 0
C29687 _0621_/a_35_297# clknet_1_1__leaf__0458_ 0.037f
C29688 acc0.A\[12\] _1057_/a_891_413# 0.05073f
C29689 _0998_/a_193_47# clknet_1_1__leaf__0461_ 0.00162f
C29690 VPWR _0701_/a_303_47# 0
C29691 VPWR _0603_/a_68_297# 0.15264f
C29692 _0662_/a_384_47# _0423_ 0
C29693 _0662_/a_81_21# _0401_ 0.00105f
C29694 _0662_/a_299_297# _0290_ 0.0335f
C29695 _0259_ _0815_/a_113_297# 0
C29696 _0239_ _0399_ 0
C29697 VPWR hold73/a_391_47# 0.1888f
C29698 _1033_/a_1017_47# net17 0
C29699 pp[29] _0221_ 0
C29700 _0457_ _1032_/a_634_159# 0.00851f
C29701 _0278_ _0280_ 0
C29702 VPWR _0657_/a_109_297# 0.0044f
C29703 net44 _0999_/a_891_413# 0.00438f
C29704 _0226_ _0750_/a_181_47# 0.00188f
C29705 pp[30] hold16/a_49_47# 0.00892f
C29706 net59 hold16/a_391_47# 0
C29707 _0263_ _0350_ 0.04601f
C29708 _1000_/a_1059_315# net46 0.01301f
C29709 hold54/a_285_47# net23 0
C29710 _0181_ _0584_/a_373_47# 0.0034f
C29711 net22 net157 0.24782f
C29712 _0149_ clknet_1_1__leaf__0458_ 0
C29713 _1016_/a_193_47# _0218_ 0
C29714 VPWR _0999_/a_193_47# 0.33979f
C29715 hold27/a_285_47# _0536_/a_51_297# 0
C29716 _0740_/a_113_47# _0359_ 0
C29717 _1052_/a_27_47# acc0.A\[6\] 0.04532f
C29718 _0216_ _0219_ 0.76632f
C29719 hold20/a_285_47# _0487_ 0
C29720 net88 clknet_1_0__leaf__0460_ 0.1686f
C29721 net54 hold50/a_285_47# 0
C29722 _0467_ control0.sh 0
C29723 _0581_/a_27_297# _0581_/a_109_297# 0.17136f
C29724 _0225_ _0374_ 0.22981f
C29725 clknet_0__0459_ _0645_/a_285_47# 0.00499f
C29726 _0441_ net9 0
C29727 _0983_/a_27_47# net165 0
C29728 net45 _0708_/a_150_297# 0
C29729 net136 net62 0
C29730 _0245_ _0246_ 0.02845f
C29731 net233 _0446_ 0.02203f
C29732 _1039_/a_1059_315# net8 0.04314f
C29733 _0985_/a_1059_315# _0083_ 0.06121f
C29734 hold78/a_285_47# _0195_ 0
C29735 _0216_ _0728_/a_59_75# 0.00294f
C29736 _0320_ acc0.A\[25\] 0.01883f
C29737 acc0.A\[4\] _0218_ 0.05841f
C29738 _0682_/a_68_297# VPWR 0.16126f
C29739 _1018_/a_466_413# net104 0
C29740 net232 _0967_/a_215_297# 0
C29741 hold85/a_49_47# _0476_ 0.00881f
C29742 hold67/a_391_47# clknet_1_1__leaf__0465_ 0.02119f
C29743 hold19/a_391_47# _1016_/a_381_47# 0.00142f
C29744 _0343_ _0990_/a_193_47# 0.02996f
C29745 net158 _0464_ 0.02403f
C29746 comp0.B\[14\] _1046_/a_1017_47# 0
C29747 clknet_1_0__leaf__0463_ net157 0.01169f
C29748 _0302_ _0345_ 0.00183f
C29749 _0970_/a_27_297# _0485_ 0.03447f
C29750 _0970_/a_114_47# _0484_ 0.00553f
C29751 pp[2] _0642_/a_215_297# 0
C29752 _0734_/a_129_47# _0326_ 0
C29753 _1053_/a_193_47# net15 0
C29754 _0982_/a_381_47# _0982_/a_561_413# 0.00123f
C29755 _0982_/a_27_47# net68 0.22613f
C29756 _0982_/a_891_413# _0982_/a_975_413# 0.00851f
C29757 hold88/a_285_47# _0833_/a_215_47# 0
C29758 _0174_ input30/a_75_212# 0
C29759 net45 _0114_ 0
C29760 net45 _0615_/a_109_297# 0.00157f
C29761 _1049_/a_466_413# _1049_/a_592_47# 0.00553f
C29762 _1049_/a_634_159# _1049_/a_1017_47# 0
C29763 hold65/a_391_47# _0433_ 0
C29764 control0.sh comp0.B\[0\] 0
C29765 _0334_ hold61/a_285_47# 0
C29766 net48 _0603_/a_68_297# 0.11848f
C29767 acc0.A\[8\] net47 0.02354f
C29768 net48 hold73/a_391_47# 0.06535f
C29769 control0.count\[3\] _0486_ 0.00536f
C29770 _0598_/a_79_21# _0373_ 0
C29771 net39 _0277_ 0
C29772 hold48/a_49_47# _0172_ 0
C29773 net68 _0145_ 0
C29774 _0473_ _1044_/a_27_47# 0
C29775 _1070_/a_27_47# _1070_/a_193_47# 0.97453f
C29776 net10 _1061_/a_1059_315# 0
C29777 _1053_/a_634_159# _1053_/a_466_413# 0.23992f
C29778 _1053_/a_193_47# _1053_/a_1059_315# 0.03405f
C29779 _1053_/a_27_47# _1053_/a_891_413# 0.03224f
C29780 _0269_ _0635_/a_27_47# 0
C29781 _0714_/a_512_297# _0218_ 0
C29782 net203 _0133_ 0
C29783 net192 net37 0
C29784 _0195_ _1008_/a_1059_315# 0
C29785 _0996_/a_193_47# _0181_ 0
C29786 _1066_/a_466_413# _1066_/a_592_47# 0.00553f
C29787 _1066_/a_634_159# _1066_/a_1017_47# 0
C29788 _0179_ input16/a_75_212# 0
C29789 _1046_/a_891_413# comp0.B\[9\] 0
C29790 _0339_ _0345_ 0.14468f
C29791 _0991_/a_193_47# net47 0.03112f
C29792 _1037_/a_27_47# _0176_ 0.00304f
C29793 hold34/a_285_47# A[12] 0.0019f
C29794 _1034_/a_193_47# _0175_ 0.03455f
C29795 pp[9] net2 0
C29796 pp[6] _0253_ 0.00304f
C29797 _1056_/a_193_47# _0343_ 0
C29798 net31 _1040_/a_466_413# 0
C29799 net109 _1022_/a_27_47# 0.03338f
C29800 _0833_/a_215_47# _0086_ 0.00313f
C29801 _0680_/a_300_47# _0462_ 0
C29802 _0346_ net37 0
C29803 _1068_/a_466_413# _1068_/a_592_47# 0.00553f
C29804 _1068_/a_634_159# _1068_/a_1017_47# 0
C29805 _0222_ hold94/a_285_47# 0.01187f
C29806 clkbuf_1_1__f__0464_/a_110_47# _1044_/a_27_47# 0.02569f
C29807 _1030_/a_193_47# _1030_/a_381_47# 0.09799f
C29808 _1030_/a_634_159# _1030_/a_891_413# 0.03684f
C29809 _1030_/a_27_47# _1030_/a_561_413# 0.0027f
C29810 _1041_/a_466_413# _0176_ 0
C29811 _0712_/a_381_47# _0339_ 0.01168f
C29812 clknet_1_0__leaf__0461_ _0350_ 0.31323f
C29813 _0156_ net67 0
C29814 hold74/a_49_47# clknet_1_0__leaf__0459_ 0.00847f
C29815 _0294_ _0116_ 0
C29816 VPWR _0163_ 0.30979f
C29817 _0286_ acc0.A\[10\] 0
C29818 _1017_/a_193_47# _0352_ 0
C29819 net24 _0560_/a_68_297# 0
C29820 _0461_ _0616_/a_78_199# 0.00129f
C29821 _0218_ _0807_/a_68_297# 0.18943f
C29822 hold41/a_391_47# A[12] 0
C29823 _0311_ clknet_1_0__leaf__0459_ 0
C29824 hold100/a_49_47# _0637_/a_56_297# 0
C29825 VPWR _0570_/a_27_297# 0.25572f
C29826 _0571_/a_109_297# clknet_1_1__leaf__0462_ 0
C29827 _1035_/a_561_413# clknet_1_1__leaf__0463_ 0
C29828 _1035_/a_891_413# net122 0
C29829 _0753_/a_465_47# net46 0
C29830 _0992_/a_466_413# net37 0
C29831 _0346_ hold91/a_49_47# 0.01981f
C29832 _0804_/a_215_47# _0347_ 0.08582f
C29833 net248 _0836_/a_68_297# 0.09865f
C29834 _0786_/a_80_21# _0401_ 0.20799f
C29835 _0786_/a_472_297# _0423_ 0
C29836 _0786_/a_217_297# _0290_ 0
C29837 clkbuf_0__0461_/a_110_47# _0181_ 0.00436f
C29838 _0770_/a_297_47# acc0.A\[19\] 0.00702f
C29839 _0241_ _0352_ 0.02149f
C29840 _1015_/a_891_413# _0181_ 0.02041f
C29841 _0688_/a_109_297# _0360_ 0
C29842 VPWR _0517_/a_81_21# 0.23956f
C29843 _0987_/a_193_47# _0987_/a_466_413# 0.07855f
C29844 _0987_/a_27_47# _0987_/a_1059_315# 0.04875f
C29845 clknet_0__0459_ _0507_/a_27_297# 0
C29846 acc0.A\[1\] _0262_ 0
C29847 hold64/a_391_47# net211 0.1316f
C29848 net248 net212 0.00135f
C29849 net194 _1051_/a_27_47# 0
C29850 _0579_/a_27_297# _0217_ 0.09482f
C29851 _1021_/a_27_47# net106 0
C29852 _1051_/a_1017_47# _0186_ 0
C29853 hold49/a_49_47# _1044_/a_27_47# 0
C29854 net247 _0219_ 0
C29855 _0385_ _0346_ 0.01774f
C29856 acc0.A\[27\] _1008_/a_975_413# 0
C29857 clknet_0_clk _0971_/a_299_297# 0
C29858 _0992_/a_891_413# net67 0.01206f
C29859 _1000_/a_891_413# VPWR 0.17562f
C29860 clknet_0__0459_ _0716_/a_27_47# 0
C29861 _1004_/a_27_47# _1004_/a_193_47# 0.96188f
C29862 _0483_ _0467_ 0
C29863 net162 net208 0
C29864 VPWR B[9] 0.37754f
C29865 hold16/a_49_47# _0339_ 0.0033f
C29866 _0151_ _1053_/a_634_159# 0
C29867 net45 clkload3/Y 0.0055f
C29868 control0.state\[2\] clkbuf_1_0__f_clk/a_110_47# 0
C29869 _0345_ net6 0.01921f
C29870 pp[27] hold61/a_49_47# 0.00614f
C29871 _0718_/a_47_47# net56 0
C29872 _0225_ _0249_ 0.13043f
C29873 _0608_/a_109_297# _0219_ 0
C29874 hold77/a_285_47# net96 0
C29875 clknet_1_1__leaf__0462_ _0737_/a_285_297# 0
C29876 net113 _0737_/a_35_297# 0
C29877 net9 hold83/a_49_47# 0
C29878 _0346_ _1006_/a_1017_47# 0
C29879 net58 net77 0
C29880 _1029_/a_27_47# _1029_/a_1059_315# 0.04875f
C29881 _1029_/a_193_47# _1029_/a_466_413# 0.08301f
C29882 VPWR hold50/a_49_47# 0.32783f
C29883 clknet_1_0__leaf__0459_ _0583_/a_27_297# 0.01509f
C29884 net64 net47 0.02519f
C29885 hold21/a_49_47# _0186_ 0
C29886 _0482_ hold79/a_285_47# 0
C29887 _0856_/a_79_21# _0346_ 0.19351f
C29888 _0096_ _0097_ 0
C29889 _0218_ net41 0.01904f
C29890 _0352_ _0772_/a_510_47# 0.00574f
C29891 _0770_/a_297_47# _0249_ 0
C29892 _0095_ _0406_ 0
C29893 _0844_/a_382_297# _0219_ 0
C29894 _1032_/a_592_47# clknet_1_0__leaf__0461_ 0.00107f
C29895 net240 _0487_ 0.1965f
C29896 net39 _0298_ 0.05296f
C29897 acc0.A\[12\] _0404_ 0.04613f
C29898 net175 _0197_ 0.23133f
C29899 _0805_/a_27_47# _0419_ 0.00782f
C29900 _0805_/a_181_47# _0417_ 0
C29901 net61 _0270_ 0.01884f
C29902 _0637_/a_56_297# _0450_ 0.00865f
C29903 _0343_ _0998_/a_561_413# 0
C29904 _0722_/a_510_47# clknet_1_1__leaf__0462_ 0
C29905 clkload0/a_27_47# _1072_/a_193_47# 0.0034f
C29906 hold65/a_49_47# VPWR 0.26835f
C29907 _0399_ _0580_/a_373_47# 0
C29908 _0722_/a_79_21# _0778_/a_68_297# 0
C29909 comp0.B\[13\] _1045_/a_466_413# 0
C29910 _0172_ net12 0
C29911 _1050_/a_193_47# _0085_ 0
C29912 hold33/a_391_47# hold26/a_285_47# 0.00144f
C29913 _1015_/a_27_47# _0565_/a_512_297# 0
C29914 _0716_/a_27_47# _0655_/a_109_93# 0
C29915 clknet_1_0__leaf__0465_ _0536_/a_240_47# 0
C29916 hold97/a_49_47# _0345_ 0.04665f
C29917 clknet_1_0__leaf__0463_ _0550_/a_240_47# 0.04777f
C29918 net144 net3 0.07547f
C29919 output43/a_27_47# _1013_/a_1059_315# 0.00111f
C29920 _1017_/a_1059_315# _1016_/a_891_413# 0.01084f
C29921 _1017_/a_891_413# _1016_/a_1059_315# 0.0034f
C29922 _0783_/a_297_297# net43 0
C29923 _0430_ _0254_ 0.01816f
C29924 _0998_/a_381_47# acc0.A\[17\] 0
C29925 clkbuf_1_1__f__0463_/a_110_47# _0113_ 0
C29926 net166 _1060_/a_466_413# 0
C29927 control0.reset _0495_/a_150_297# 0
C29928 _1037_/a_1059_315# clknet_1_1__leaf__0463_ 0
C29929 _1033_/a_634_159# _0956_/a_32_297# 0.00136f
C29930 _0960_/a_27_47# _0976_/a_76_199# 0
C29931 _1028_/a_27_47# _1028_/a_466_413# 0.26005f
C29932 _1028_/a_193_47# _1028_/a_634_159# 0.11072f
C29933 hold89/a_49_47# _0958_/a_27_47# 0
C29934 hold23/a_49_47# _0446_ 0
C29935 hold41/a_285_47# _1057_/a_634_159# 0
C29936 _0629_/a_59_75# _0856_/a_79_21# 0
C29937 _0657_/a_109_297# _0283_ 0
C29938 _0465_ _0495_/a_68_297# 0
C29939 clkbuf_1_0__f__0459_/a_110_47# clknet_1_1__leaf__0461_ 0
C29940 _0195_ hold60/a_49_47# 0.04489f
C29941 _0999_/a_27_47# _0783_/a_297_297# 0
C29942 _0999_/a_193_47# _0783_/a_79_21# 0
C29943 _0308_ _1009_/a_1059_315# 0
C29944 _0394_ _1009_/a_193_47# 0
C29945 _1033_/a_193_47# comp0.B\[1\] 0
C29946 _1033_/a_1059_315# _0131_ 0
C29947 _0985_/a_466_413# VPWR 0.25541f
C29948 net63 _0987_/a_891_413# 0.00652f
C29949 _0965_/a_285_47# _0478_ 0.0744f
C29950 VPWR _1018_/a_634_159# 0.17825f
C29951 _0130_ _1033_/a_381_47# 0
C29952 _0343_ _0438_ 0
C29953 VPWR _1049_/a_27_47# 0.69988f
C29954 _0953_/a_32_297# _0176_ 0
C29955 net226 _0162_ 0
C29956 _1037_/a_1059_315# net8 0
C29957 _0647_/a_47_47# clknet_1_1__leaf__0459_ 0.05494f
C29958 _0743_/a_512_297# _0366_ 0
C29959 _0743_/a_51_297# _0367_ 0.08265f
C29960 hold22/a_391_47# _0179_ 0.00312f
C29961 _1009_/a_975_413# _0219_ 0.00137f
C29962 _0234_ net46 0.23835f
C29963 net61 net233 0
C29964 VPWR _1066_/a_27_47# 0.69886f
C29965 _1050_/a_592_47# acc0.A\[4\] 0.00257f
C29966 net44 acc0.A\[17\] 0.85392f
C29967 _0833_/a_79_21# clkbuf_1_1__f__0458_/a_110_47# 0.01178f
C29968 _0107_ _0315_ 0
C29969 VPWR _1068_/a_27_47# 0.39963f
C29970 _0459_ clkbuf_0__0459_/a_110_47# 0.31483f
C29971 _1041_/a_1059_315# _0139_ 0
C29972 acc0.A\[0\] _0345_ 0
C29973 _0476_ net17 0.02965f
C29974 _0349_ _0725_/a_80_21# 0
C29975 VPWR _0677_/a_285_47# 0
C29976 hold37/a_285_47# hold37/a_391_47# 0.41909f
C29977 _0454_ _0346_ 0.22696f
C29978 hold13/a_49_47# clkbuf_0__0463_/a_110_47# 0
C29979 _0257_ hold101/a_285_47# 0.00216f
C29980 clkbuf_0__0462_/a_110_47# _0181_ 0
C29981 _0226_ _0606_/a_109_53# 0.00512f
C29982 _0230_ _0606_/a_215_297# 0
C29983 _0993_/a_27_47# _0417_ 0
C29984 _0993_/a_1059_315# net79 0
C29985 _0983_/a_1059_315# _1018_/a_1059_315# 0
C29986 VPWR _1034_/a_561_413# 0.00213f
C29987 hold66/a_49_47# _0228_ 0.02445f
C29988 clknet_1_0__leaf__0460_ _1067_/a_891_413# 0.03754f
C29989 hold42/a_285_47# _0179_ 0.05134f
C29990 _0179_ _1057_/a_1059_315# 0
C29991 _0140_ _1043_/a_27_47# 0
C29992 net18 _1043_/a_466_413# 0.01599f
C29993 net198 _1043_/a_1059_315# 0.00309f
C29994 _1004_/a_27_47# net199 0
C29995 hold34/a_285_47# _0154_ 0.00753f
C29996 VPWR hold6/a_285_47# 0.28449f
C29997 clknet_1_0__leaf__0464_ _0528_/a_81_21# 0.07721f
C29998 clknet_1_0__leaf__0465_ _1046_/a_27_47# 0.00917f
C29999 net87 _0181_ 0
C30000 _0343_ _0983_/a_466_413# 0.00369f
C30001 VPWR _0816_/a_150_297# 0.00122f
C30002 _1057_/a_27_47# _0181_ 0.00421f
C30003 _0578_/a_27_297# _0460_ 0
C30004 _0578_/a_109_47# clknet_1_0__leaf__0457_ 0
C30005 _0346_ _0505_/a_27_297# 0
C30006 acc0.A\[0\] hold2/a_49_47# 0.29408f
C30007 _1053_/a_891_413# A[5] 0
C30008 _0718_/a_47_47# _0345_ 0.00134f
C30009 _0143_ net130 0
C30010 _0399_ _0309_ 0
C30011 _1002_/a_1059_315# acc0.A\[20\] 0
C30012 _0998_/a_634_159# _0998_/a_381_47# 0
C30013 net44 net60 0
C30014 comp0.B\[15\] _0208_ 0.78234f
C30015 _0195_ hold61/a_391_47# 0
C30016 clkbuf_0__0457_/a_110_47# _0099_ 0
C30017 net64 _0988_/a_592_47# 0.00256f
C30018 net45 net104 0.00355f
C30019 _1059_/a_381_47# _0459_ 0.00147f
C30020 _0529_/a_27_297# _0186_ 0.12525f
C30021 _0779_/a_79_21# _0306_ 0
C30022 net90 acc0.A\[23\] 0
C30023 _1003_/a_1059_315# _0369_ 0.0018f
C30024 net243 clknet_1_0__leaf__0460_ 0.00218f
C30025 net205 comp0.B\[4\] 0.07202f
C30026 _0498_/a_240_47# _1061_/a_193_47# 0
C30027 VPWR _0708_/a_150_297# 0.00193f
C30028 _0122_ _1023_/a_634_159# 0
C30029 net110 _1023_/a_466_413# 0
C30030 hold56/a_391_47# _1033_/a_193_47# 0.00147f
C30031 hold56/a_49_47# _1033_/a_466_413# 0.00218f
C30032 _0662_/a_299_297# _0986_/a_1059_315# 0
C30033 _0244_ clknet_1_0__leaf__0461_ 0.04827f
C30034 clkbuf_1_1__f__0463_/a_110_47# comp0.B\[3\] 0
C30035 _0310_ _0306_ 0.01383f
C30036 _0443_ _0254_ 0.24908f
C30037 _0097_ _0395_ 0.00447f
C30038 _0176_ _0561_/a_51_297# 0
C30039 _1019_/a_634_159# _1019_/a_1059_315# 0
C30040 _1019_/a_27_47# _1019_/a_381_47# 0.05761f
C30041 _1019_/a_193_47# _1019_/a_891_413# 0.19421f
C30042 _0717_/a_209_297# _0221_ 0.08327f
C30043 hold76/a_49_47# _0216_ 0.02113f
C30044 _0578_/a_27_297# _0457_ 0
C30045 _0847_/a_109_297# _0263_ 0.00285f
C30046 _0557_/a_149_47# net171 0
C30047 _1056_/a_561_413# _0153_ 0
C30048 _0467_ _0955_/a_32_297# 0
C30049 _0227_ _0352_ 0.0366f
C30050 _0837_/a_266_47# _0172_ 0.04448f
C30051 net123 net29 0.07175f
C30052 net72 _0986_/a_27_47# 0.21487f
C30053 clknet_1_1__leaf__0458_ _0986_/a_634_159# 0
C30054 VPWR _1041_/a_1017_47# 0
C30055 VPWR _1012_/a_466_413# 0.26178f
C30056 _0231_ _0225_ 0.13857f
C30057 hold52/a_391_47# _1024_/a_1059_315# 0.00131f
C30058 _0548_/a_149_47# _1040_/a_1059_315# 0
C30059 _0475_ _0496_/a_27_47# 0.0569f
C30060 VPWR _0615_/a_109_297# 0.00696f
C30061 VPWR _0114_ 0.36448f
C30062 _0294_ _0370_ 0
C30063 _1050_/a_27_47# net184 0
C30064 _1050_/a_193_47# net131 0.00186f
C30065 clknet_1_0__leaf__0462_ net49 0.03458f
C30066 hold24/a_285_47# _0549_/a_68_297# 0
C30067 clknet_1_0__leaf__0463_ net172 0.21419f
C30068 net129 _0141_ 0
C30069 _0580_/a_109_297# _0345_ 0.00482f
C30070 net9 _1049_/a_891_413# 0.01819f
C30071 _0133_ _0176_ 0
C30072 _0289_ _0426_ 0
C30073 clknet_1_1__leaf__0459_ _0998_/a_891_413# 0.0087f
C30074 _0718_/a_47_47# hold16/a_49_47# 0
C30075 _0210_ _0474_ 0
C30076 _1001_/a_27_47# net187 0
C30077 net162 _1031_/a_193_47# 0.02645f
C30078 _0955_/a_32_297# comp0.B\[0\] 0
C30079 _0982_/a_193_47# net207 0
C30080 _0534_/a_81_21# _0178_ 0.01158f
C30081 _0758_/a_297_297# _0347_ 0
C30082 _1024_/a_891_413# net52 0.02618f
C30083 clknet_0__0458_ _0826_/a_27_53# 0.01953f
C30084 _0294_ _0991_/a_193_47# 0.03812f
C30085 _0991_/a_27_47# _0218_ 0
C30086 _0581_/a_109_297# _0116_ 0.0568f
C30087 _0990_/a_193_47# _0990_/a_381_47# 0.09799f
C30088 _0990_/a_634_159# _0990_/a_891_413# 0.03684f
C30089 _0990_/a_27_47# _0990_/a_561_413# 0.00163f
C30090 _0352_ _0687_/a_59_75# 0
C30091 _0343_ _0354_ 0.00473f
C30092 pp[28] _0703_/a_109_297# 0.00109f
C30093 _0404_ net42 0
C30094 hold81/a_49_47# _0806_/a_113_297# 0.04306f
C30095 _0790_/a_285_297# _0345_ 0.00212f
C30096 _1002_/a_193_47# clknet_1_0__leaf__0457_ 0.00254f
C30097 _0350_ _0105_ 0
C30098 _0380_ net93 0
C30099 _0343_ clknet_1_1__leaf__0465_ 0.09287f
C30100 _0747_/a_215_47# _0352_ 0.01145f
C30101 _0174_ _0546_/a_149_47# 0.02512f
C30102 acc0.A\[22\] _0228_ 0
C30103 net203 _0208_ 0.07866f
C30104 _0967_/a_215_297# _0967_/a_297_297# 0.01452f
C30105 _0967_/a_109_93# _0967_/a_403_297# 0
C30106 acc0.A\[25\] _1007_/a_1059_315# 0.00288f
C30107 _0967_/a_215_297# _0162_ 0
C30108 _0967_/a_487_297# _0485_ 0.00421f
C30109 _0466_ _0975_/a_59_75# 0
C30110 _0488_ _0975_/a_145_75# 0
C30111 hold97/a_285_47# _0329_ 0
C30112 _0695_/a_80_21# acc0.A\[24\] 0
C30113 clkbuf_1_0__f__0465_/a_110_47# _0256_ 0.00108f
C30114 _0539_/a_68_297# clknet_1_1__leaf__0464_ 0
C30115 _0179_ _0255_ 0
C30116 _0805_/a_27_47# _0992_/a_193_47# 0
C30117 hold53/a_285_47# _1025_/a_634_159# 0
C30118 hold53/a_391_47# _1025_/a_193_47# 0
C30119 _1049_/a_381_47# acc0.A\[3\] 0
C30120 _1049_/a_592_47# _0147_ 0.00188f
C30121 _0195_ clknet_1_1__leaf__0462_ 0.50267f
C30122 hold25/a_285_47# _1040_/a_381_47# 0
C30123 VPWR net98 0.40249f
C30124 hold9/a_391_47# _0739_/a_215_47# 0
C30125 _0848_/a_27_47# _0350_ 0.00471f
C30126 VPWR _0653_/a_113_47# 0
C30127 net216 _0371_ 0.45055f
C30128 _0536_/a_149_47# _0463_ 0
C30129 _0230_ hold3/a_49_47# 0
C30130 _0226_ hold3/a_285_47# 0.00201f
C30131 net243 _0576_/a_109_297# 0
C30132 net248 _0989_/a_891_413# 0
C30133 VPWR input6/a_75_212# 0.29205f
C30134 _0606_/a_215_297# _0236_ 0.16838f
C30135 _0218_ _0350_ 0.64828f
C30136 _0245_ _0774_/a_68_297# 0
C30137 _1045_/a_27_47# _1045_/a_634_159# 0.14145f
C30138 _1070_/a_466_413# _1070_/a_592_47# 0.00553f
C30139 _1070_/a_27_47# VPWR 0.67875f
C30140 _1070_/a_634_159# _1070_/a_1017_47# 0
C30141 _1052_/a_891_413# _0150_ 0.01106f
C30142 _0343_ _0693_/a_68_297# 0
C30143 pp[17] _1030_/a_891_413# 0
C30144 clkbuf_0__0461_/a_110_47# clknet_1_1__leaf__0461_ 0
C30145 clknet_1_0__leaf__0465_ _1050_/a_1017_47# 0
C30146 _0111_ _0218_ 0.18742f
C30147 net45 _0998_/a_592_47# 0
C30148 _0146_ _1061_/a_1059_315# 0
C30149 _0577_/a_109_297# net177 0
C30150 _1066_/a_381_47# control0.sh 0
C30151 hold21/a_285_47# _0518_/a_109_297# 0
C30152 _1014_/a_466_413# _0465_ 0
C30153 _0552_/a_68_297# input29/a_75_212# 0
C30154 _1062_/a_466_413# _0468_ 0
C30155 clkload3/Y VPWR 0.42401f
C30156 VPWR _1030_/a_466_413# 0.24842f
C30157 _0995_/a_466_413# net43 0
C30158 clknet_1_1__leaf__0463_ _0561_/a_240_47# 0.00193f
C30159 _0327_ net96 0
C30160 _0683_/a_113_47# net93 0
C30161 _0314_ _1007_/a_1017_47# 0
C30162 _1043_/a_27_47# _1043_/a_634_159# 0.14145f
C30163 net7 _1040_/a_466_413# 0
C30164 net1 control0.sh 0
C30165 comp0.B\[2\] _0564_/a_68_297# 0
C30166 _0217_ net36 0.02633f
C30167 A[3] input18/a_75_212# 0.00693f
C30168 input10/a_75_212# B[10] 0
C30169 net31 net174 0.00299f
C30170 _1017_/a_634_159# hold72/a_49_47# 0.00127f
C30171 _1017_/a_27_47# hold72/a_391_47# 0.00249f
C30172 _1017_/a_193_47# hold72/a_285_47# 0.00356f
C30173 net177 _1022_/a_1017_47# 0
C30174 _0997_/a_891_413# net83 0
C30175 _1038_/a_193_47# _0209_ 0.00741f
C30176 _1030_/a_193_47# _0568_/a_27_297# 0
C30177 _1030_/a_27_47# _0568_/a_109_297# 0
C30178 net236 _0975_/a_59_75# 0.00235f
C30179 clknet_1_1__leaf__0463_ _0472_ 0
C30180 _1004_/a_27_47# VPWR 0.62976f
C30181 hold67/a_285_47# _0399_ 0.00238f
C30182 _1021_/a_193_47# _1002_/a_193_47# 0
C30183 _1021_/a_634_159# _1002_/a_27_47# 0
C30184 net80 _0218_ 0.1762f
C30185 comp0.B\[2\] clknet_1_1__leaf_clk 0
C30186 _1021_/a_27_47# _1002_/a_634_159# 0
C30187 clknet_1_0__leaf__0458_ _1047_/a_634_159# 0
C30188 net138 net13 0.02502f
C30189 acc0.A\[12\] _0419_ 0
C30190 hold100/a_285_47# _0269_ 0.00448f
C30191 VPWR _0126_ 0.25857f
C30192 net182 _0517_/a_81_21# 0
C30193 _0645_/a_47_47# _0277_ 0.14441f
C30194 clknet_1_0__leaf__0465_ net63 0.03847f
C30195 _1056_/a_193_47# _1056_/a_381_47# 0.09799f
C30196 _1056_/a_634_159# _1056_/a_891_413# 0.03684f
C30197 _1056_/a_27_47# _1056_/a_561_413# 0.0027f
C30198 _0671_/a_113_297# _0303_ 0.15241f
C30199 hold28/a_49_47# acc0.A\[1\] 0
C30200 _0322_ _0315_ 0.09044f
C30201 _0294_ _0423_ 0.25223f
C30202 _0270_ _0431_ 0
C30203 clknet_0__0459_ _0185_ 0
C30204 net194 _1044_/a_193_47# 0.27488f
C30205 _0987_/a_193_47# _0085_ 0.41169f
C30206 _0987_/a_891_413# _0987_/a_1017_47# 0.00617f
C30207 clknet_1_1__leaf__0459_ _0287_ 0
C30208 _0987_/a_634_159# net73 0
C30209 hold78/a_49_47# pp[31] 0.00102f
C30210 hold74/a_391_47# _0399_ 0
C30211 hold87/a_285_47# _0241_ 0
C30212 _0366_ clknet_1_0__leaf__0460_ 0.00297f
C30213 _0327_ _0315_ 0.0258f
C30214 _0833_/a_297_297# acc0.A\[8\] 0
C30215 _0348_ hold16/a_285_47# 0
C30216 hold39/a_49_47# net24 0
C30217 _0661_/a_277_297# VPWR 0
C30218 _0849_/a_79_21# _0450_ 0
C30219 acc0.A\[1\] _1047_/a_592_47# 0
C30220 _0180_ _1047_/a_561_413# 0
C30221 _0239_ _0306_ 0.30294f
C30222 net194 net131 0.05026f
C30223 net8 _0472_ 0.08515f
C30224 _0145_ hold71/a_49_47# 0
C30225 _1041_/a_27_47# _0548_/a_512_297# 0
C30226 _0343_ _0567_/a_27_297# 0.00209f
C30227 _1004_/a_634_159# _1004_/a_1017_47# 0
C30228 _1004_/a_466_413# _1004_/a_592_47# 0.00553f
C30229 _0195_ net242 0.01189f
C30230 _1027_/a_1059_315# _1008_/a_466_413# 0
C30231 _1027_/a_634_159# _1008_/a_891_413# 0
C30232 _1027_/a_891_413# _1008_/a_634_159# 0
C30233 _1027_/a_466_413# _1008_/a_1059_315# 0
C30234 clkbuf_1_0__f__0462_/a_110_47# acc0.A\[25\] 0.0046f
C30235 net157 _1049_/a_381_47# 0
C30236 _0151_ net139 0.07095f
C30237 hold78/a_49_47# hold15/a_285_47# 0
C30238 acc0.A\[31\] _0712_/a_465_47# 0
C30239 _0196_ _0186_ 0.07026f
C30240 _1067_/a_466_413# hold93/a_285_47# 0.00105f
C30241 _0680_/a_300_47# _0312_ 0.00403f
C30242 _0098_ clkbuf_0__0461_/a_110_47# 0.00123f
C30243 _0593_/a_113_47# VPWR 0
C30244 _1029_/a_891_413# _1029_/a_1017_47# 0.00617f
C30245 _1029_/a_193_47# net191 0.2401f
C30246 clknet_1_0__leaf__0459_ _0114_ 0.49016f
C30247 _1019_/a_466_413# _0352_ 0
C30248 net1 net157 0.0486f
C30249 _0625_/a_59_75# acc0.A\[5\] 0.08092f
C30250 output46/a_27_47# net46 0.21644f
C30251 _0343_ _0800_/a_51_297# 0
C30252 hold69/a_391_47# _0250_ 0.00578f
C30253 _0535_/a_68_297# _0176_ 0.14003f
C30254 VPWR _0531_/a_109_47# 0.0014f
C30255 _0462_ acc0.A\[19\] 0.0064f
C30256 comp0.B\[13\] net184 0.00192f
C30257 acc0.A\[4\] _0987_/a_592_47# 0.00105f
C30258 net213 _0345_ 0
C30259 _0514_/a_27_297# net143 0
C30260 _1000_/a_634_159# acc0.A\[18\] 0
C30261 _1015_/a_1059_315# net201 0
C30262 hold47/a_49_47# _0180_ 0.04107f
C30263 acc0.A\[10\] net79 0
C30264 _1020_/a_634_159# _0183_ 0.00711f
C30265 _1020_/a_1059_315# _0217_ 0
C30266 clkbuf_0__0465_/a_110_47# _0271_ 0
C30267 net233 _0431_ 0
C30268 net103 _1016_/a_561_413# 0
C30269 _0292_ _0287_ 0.03881f
C30270 hold15/a_285_47# _0129_ 0.01025f
C30271 _0101_ _0596_/a_59_75# 0
C30272 _0153_ A[12] 0
C30273 net160 comp0.B\[4\] 0.13077f
C30274 _1016_/a_634_159# _1016_/a_466_413# 0.23992f
C30275 _1016_/a_193_47# _1016_/a_1059_315# 0.03405f
C30276 _1016_/a_27_47# _1016_/a_891_413# 0.02974f
C30277 hold101/a_285_47# clknet_1_1__leaf__0458_ 0.00157f
C30278 _0343_ _0829_/a_27_47# 0.00734f
C30279 hold11/a_285_47# _1061_/a_634_159# 0.00143f
C30280 _0756_/a_285_47# net109 0
C30281 clkbuf_1_0__f__0457_/a_110_47# acc0.A\[20\] 0.02614f
C30282 _0512_/a_109_297# net143 0
C30283 _0960_/a_27_47# _0488_ 0.05307f
C30284 _1028_/a_193_47# net114 0.00343f
C30285 _1028_/a_1059_315# _1028_/a_1017_47# 0
C30286 hold25/a_391_47# _1041_/a_27_47# 0
C30287 hold25/a_285_47# _1041_/a_193_47# 0
C30288 _0211_ _0549_/a_68_297# 0
C30289 hold89/a_49_47# _0477_ 0
C30290 hold41/a_49_47# net189 0
C30291 hold17/a_285_47# _1070_/a_27_47# 0
C30292 hold87/a_391_47# _0982_/a_27_47# 0
C30293 _0343_ _0996_/a_561_413# 0
C30294 hold87/a_285_47# _0982_/a_193_47# 0
C30295 _0839_/a_109_297# _0218_ 0.00144f
C30296 _1067_/a_634_159# control0.reset 0
C30297 _0369_ _0989_/a_1017_47# 0
C30298 _1057_/a_27_47# _0187_ 0.03075f
C30299 _1057_/a_634_159# net4 0
C30300 _0441_ _0255_ 0
C30301 _0593_/a_113_47# net48 0
C30302 VPWR _0990_/a_466_413# 0.26304f
C30303 _0999_/a_466_413# _0399_ 0
C30304 _0999_/a_634_159# _0096_ 0
C30305 output37/a_27_47# net67 0
C30306 hold57/a_285_47# net171 0
C30307 hold57/a_49_47# _0207_ 0
C30308 _0083_ VPWR 0.35097f
C30309 clkbuf_1_1__f__0460_/a_110_47# _0686_/a_27_53# 0
C30310 _0174_ _0176_ 0.37065f
C30311 _0514_/a_27_297# _0514_/a_109_47# 0.00393f
C30312 VPWR net104 0.36356f
C30313 pp[18] net45 0.00557f
C30314 _0130_ comp0.B\[1\] 0.05415f
C30315 _0351_ net239 0.01001f
C30316 comp0.B\[3\] _0163_ 0
C30317 _0462_ _0249_ 0.00384f
C30318 _0584_/a_27_297# _0584_/a_109_297# 0.17136f
C30319 VPWR _0651_/a_113_47# 0
C30320 _0112_ _0350_ 0
C30321 _0243_ net45 0
C30322 _0556_/a_150_297# net24 0.00133f
C30323 _0198_ _0262_ 0
C30324 _0463_ _0177_ 0
C30325 _0472_ net10 0
C30326 net217 net228 0.03719f
C30327 _1017_/a_634_159# clknet_0__0461_ 0
C30328 _1041_/a_592_47# net31 0.00266f
C30329 _0460_ _1006_/a_381_47# 0.00475f
C30330 net183 clknet_1_1__leaf__0464_ 0
C30331 _0490_ _0480_ 0
C30332 clknet_1_0__leaf__0462_ _0757_/a_68_297# 0.00467f
C30333 _0483_ _0961_/a_113_297# 0
C30334 _0170_ _1072_/a_193_47# 0.27573f
C30335 _1010_/a_891_413# clknet_1_1__leaf__0462_ 0.00425f
C30336 _0753_/a_79_21# _0754_/a_51_297# 0.00133f
C30337 hold57/a_285_47# net24 0
C30338 _0562_/a_68_297# _0213_ 0
C30339 net34 _0488_ 0.13492f
C30340 control0.state\[1\] _0466_ 0.16387f
C30341 _0738_/a_150_297# _0345_ 0.00149f
C30342 _0275_ _0345_ 0.00257f
C30343 _0783_/a_215_47# clknet_1_1__leaf__0461_ 0.00219f
C30344 _0275_ _0814_/a_27_47# 0
C30345 net123 comp0.B\[6\] 0
C30346 _0730_/a_297_297# _0195_ 0
C30347 _0601_/a_68_297# _0368_ 0
C30348 clknet_1_0__leaf__0462_ _1025_/a_193_47# 0.04215f
C30349 _1056_/a_466_413# VPWR 0.24907f
C30350 _0226_ _0238_ 0.00347f
C30351 _0175_ _0171_ 0.04288f
C30352 hold87/a_391_47# _0446_ 0
C30353 hold87/a_285_47# _0450_ 0
C30354 clknet_1_1__leaf__0463_ B[4] 0.0126f
C30355 _0195_ hold92/a_49_47# 0
C30356 net58 _0852_/a_285_297# 0
C30357 hold86/a_391_47# _0350_ 0
C30358 _1041_/a_27_47# input7/a_75_212# 0
C30359 _0244_ _0218_ 0.24397f
C30360 _0386_ _0294_ 0.002f
C30361 net18 net196 0
C30362 net54 VPWR 1.36013f
C30363 output36/a_27_47# clknet_1_0__leaf__0463_ 0.00344f
C30364 _0446_ _0529_/a_109_297# 0
C30365 hold85/a_391_47# _0468_ 0
C30366 _1028_/a_193_47# _0365_ 0
C30367 _0271_ _0824_/a_59_75# 0.15941f
C30368 _0996_/a_381_47# net5 0.0205f
C30369 _0346_ _0184_ 0
C30370 clknet_0_clk _1068_/a_1059_315# 0
C30371 acc0.A\[14\] net166 0
C30372 _0337_ _0219_ 0
C30373 _0227_ _0237_ 0.4338f
C30374 _0998_/a_381_47# net84 0.02207f
C30375 net45 _0407_ 0.00153f
C30376 comp0.B\[2\] _1015_/a_1059_315# 0
C30377 _1020_/a_891_413# control0.add 0
C30378 net178 _1055_/a_466_413# 0
C30379 _1021_/a_27_47# net220 0
C30380 clknet_1_1__leaf__0460_ acc0.A\[29\] 0.00493f
C30381 _0552_/a_68_297# net180 0
C30382 clknet_1_0__leaf__0460_ _0378_ 0.02875f
C30383 net7 _0465_ 0
C30384 _0961_/a_113_297# control0.count\[1\] 0.05194f
C30385 _0159_ _1061_/a_466_413# 0
C30386 net7 _1061_/a_381_47# 0.00842f
C30387 _1010_/a_1059_315# _0720_/a_68_297# 0
C30388 _0251_ _0825_/a_68_297# 0
C30389 _1024_/a_1017_47# acc0.A\[23\] 0
C30390 net110 net177 0
C30391 hold56/a_285_47# net119 0.01541f
C30392 VPWR _0806_/a_199_47# 0
C30393 _0984_/a_561_413# net47 0
C30394 control0.state\[1\] net236 0.11759f
C30395 clkbuf_1_0__f__0461_/a_110_47# net223 0.00203f
C30396 _0350_ _0099_ 0
C30397 _0176_ _0208_ 0.69195f
C30398 _0792_/a_80_21# net41 0.01397f
C30399 _1019_/a_1059_315# net105 0
C30400 _1019_/a_466_413# net207 0.00256f
C30401 _0714_/a_149_47# _0714_/a_240_47# 0.06872f
C30402 net58 net247 0.08215f
C30403 _0965_/a_47_47# control0.count\[3\] 0.09463f
C30404 hold18/a_391_47# _0263_ 0
C30405 net51 _1005_/a_466_413# 0
C30406 _0467_ _0474_ 0
C30407 hold98/a_285_47# _0297_ 0
C30408 net36 clknet_0__0463_ 0.01581f
C30409 _0270_ _0269_ 0
C30410 clknet_1_1__leaf__0460_ _0699_/a_68_297# 0.05396f
C30411 net126 input30/a_75_212# 0
C30412 _0725_/a_209_47# _0333_ 0
C30413 VPWR _0584_/a_27_297# 0.24873f
C30414 _0760_/a_47_47# hold3/a_285_47# 0
C30415 hold52/a_49_47# acc0.A\[24\] 0.3237f
C30416 hold83/a_285_47# net13 0.00283f
C30417 _0548_/a_240_47# net174 0
C30418 _1014_/a_27_47# clknet_1_0__leaf__0461_ 0.04214f
C30419 _0537_/a_68_297# _0537_/a_150_297# 0.00477f
C30420 clkbuf_1_0__f__0463_/a_110_47# comp0.B\[10\] 0
C30421 _0726_/a_245_297# _0355_ 0
C30422 _0726_/a_51_297# net227 0.1473f
C30423 acc0.A\[12\] _0992_/a_193_47# 0
C30424 _0172_ hold6/a_49_47# 0.00209f
C30425 _0359_ _0350_ 0.0424f
C30426 _1058_/a_1017_47# net67 0
C30427 comp0.B\[7\] _0207_ 0
C30428 _0535_/a_150_297# _0139_ 0
C30429 _1033_/a_27_47# net202 0
C30430 net119 _1032_/a_193_47# 0
C30431 net242 _1010_/a_891_413# 0.00406f
C30432 _0287_ _0655_/a_215_53# 0.12163f
C30433 _0465_ _0844_/a_297_47# 0
C30434 net34 _1064_/a_27_47# 0.42877f
C30435 control0.state\[0\] _1064_/a_634_159# 0
C30436 control0.state\[1\] _1064_/a_193_47# 0
C30437 _0178_ hold71/a_391_47# 0
C30438 _0272_ _0826_/a_219_297# 0
C30439 _0402_ hold70/a_285_47# 0.00348f
C30440 _0996_/a_193_47# clkbuf_1_1__f__0459_/a_110_47# 0
C30441 _1033_/a_27_47# clknet_1_1__leaf__0463_ 0.00692f
C30442 net44 net84 0
C30443 _0130_ _1032_/a_634_159# 0
C30444 input30/a_75_212# input8/a_75_212# 0.01223f
C30445 _1015_/a_466_413# _0584_/a_27_297# 0
C30446 _1015_/a_634_159# _0584_/a_109_297# 0
C30447 _1070_/a_466_413# _0976_/a_76_199# 0
C30448 _1050_/a_193_47# net170 0
C30449 _1001_/a_193_47# _0247_ 0
C30450 net187 _0772_/a_79_21# 0
C30451 _0951_/a_109_93# hold84/a_285_47# 0
C30452 net245 _0800_/a_512_297# 0
C30453 _0674_/a_113_47# _0219_ 0
C30454 _1059_/a_193_47# _0508_/a_299_297# 0
C30455 net8 net149 0
C30456 _0195_ _0263_ 0
C30457 _0474_ comp0.B\[0\] 0
C30458 acc0.A\[2\] _0844_/a_297_47# 0
C30459 clkbuf_1_0__f__0457_/a_110_47# _1001_/a_193_47# 0.0017f
C30460 _1020_/a_193_47# hold40/a_391_47# 0
C30461 _0127_ hold50/a_391_47# 0
C30462 clknet_1_0__leaf__0465_ _0987_/a_1017_47# 0
C30463 _0843_/a_68_297# acc0.A\[15\] 0
C30464 _1029_/a_466_413# acc0.A\[28\] 0
C30465 _0119_ _0578_/a_27_297# 0.10955f
C30466 _0195_ _1047_/a_27_47# 0
C30467 _0596_/a_59_75# net35 0
C30468 _0779_/a_79_21# _0778_/a_68_297# 0
C30469 _0950_/a_75_212# _0161_ 0.14463f
C30470 _0465_ _1048_/a_1059_315# 0.00333f
C30471 _0965_/a_285_47# VPWR 0.00153f
C30472 _0657_/a_109_297# _0345_ 0
C30473 _1054_/a_466_413# net9 0.00194f
C30474 _0293_ _0785_/a_81_21# 0.01037f
C30475 clkbuf_1_0__f__0459_/a_110_47# clknet_1_1__leaf__0465_ 0.00105f
C30476 _0990_/a_1059_315# _0088_ 0.04879f
C30477 _0216_ _1007_/a_193_47# 0
C30478 _0769_/a_81_21# _0246_ 0.00814f
C30479 _0537_/a_68_297# VPWR 0.18608f
C30480 net125 _0498_/a_149_47# 0.00758f
C30481 _0406_ _0219_ 0.42842f
C30482 _0205_ net127 0
C30483 _1002_/a_1017_47# _0460_ 0
C30484 _0982_/a_27_47# _0264_ 0.00133f
C30485 _0999_/a_193_47# _0345_ 0
C30486 acc0.A\[2\] _1048_/a_1059_315# 0.08549f
C30487 _0216_ net23 0.02163f
C30488 _0282_ clknet_1_1__leaf__0465_ 0
C30489 _0430_ _0273_ 0.09892f
C30490 _0607_/a_27_297# _1017_/a_891_413# 0
C30491 _0125_ hold8/a_49_47# 0
C30492 clknet_1_1__leaf__0459_ _0996_/a_891_413# 0
C30493 pp[19] hold29/a_49_47# 0
C30494 net46 hold29/a_391_47# 0.01397f
C30495 _0598_/a_382_297# _0382_ 0
C30496 hold65/a_391_47# _0399_ 0.06513f
C30497 _0211_ _1035_/a_27_47# 0
C30498 _0107_ _0691_/a_150_297# 0
C30499 _0564_/a_150_297# _0215_ 0
C30500 _1050_/a_891_413# _0180_ 0.01983f
C30501 _0154_ _0153_ 0
C30502 _0267_ _0845_/a_109_47# 0
C30503 _0743_/a_240_47# _0368_ 0.08035f
C30504 net233 _0269_ 0.1751f
C30505 _0958_/a_109_47# _0468_ 0
C30506 _0389_ net46 0.42818f
C30507 comp0.B\[7\] _1039_/a_1059_315# 0.13127f
C30508 clknet_1_0__leaf__0460_ acc0.A\[24\] 0.00255f
C30509 _0682_/a_68_297# _0345_ 0
C30510 _0995_/a_193_47# acc0.A\[13\] 0
C30511 _1037_/a_27_47# net28 0.00692f
C30512 _1034_/a_1059_315# comp0.B\[6\] 0.00492f
C30513 _1034_/a_891_413# comp0.B\[5\] 0
C30514 _0777_/a_377_297# clknet_1_1__leaf__0461_ 0.00128f
C30515 net57 hold80/a_285_47# 0.10679f
C30516 _1051_/a_1059_315# _1051_/a_891_413# 0.31086f
C30517 _1051_/a_193_47# _1051_/a_975_413# 0
C30518 _1051_/a_466_413# _1051_/a_381_47# 0.03733f
C30519 _1045_/a_193_47# _1044_/a_27_47# 0.01146f
C30520 _1045_/a_27_47# _1044_/a_193_47# 0.01201f
C30521 comp0.B\[14\] _1042_/a_634_159# 0
C30522 clknet_1_0__leaf__0459_ net104 0
C30523 acc0.A\[21\] _1005_/a_193_47# 0
C30524 _0227_ _1005_/a_27_47# 0.00208f
C30525 net58 _0841_/a_79_21# 0.01493f
C30526 hold15/a_285_47# hold61/a_285_47# 0
C30527 hold15/a_391_47# hold61/a_49_47# 0
C30528 _0992_/a_193_47# _0650_/a_68_297# 0
C30529 _0992_/a_27_47# _0650_/a_150_297# 0
C30530 _0411_ net6 0
C30531 acc0.A\[18\] _0242_ 0.27062f
C30532 _1070_/a_381_47# control0.count\[1\] 0
C30533 _1070_/a_592_47# _0168_ 0
C30534 net106 _1033_/a_592_47# 0
C30535 _1045_/a_891_413# _1045_/a_975_413# 0.00851f
C30536 _1045_/a_27_47# net131 0.22953f
C30537 _1045_/a_381_47# _1045_/a_561_413# 0.00123f
C30538 clkbuf_1_0__f__0464_/a_110_47# _0528_/a_81_21# 0.00788f
C30539 net1 _0462_ 0
C30540 _0979_/a_27_297# clknet_1_0__leaf_clk 0.0088f
C30541 net23 _1067_/a_27_47# 0.05974f
C30542 _0216_ _0328_ 0
C30543 _0319_ _0219_ 0
C30544 clknet_0__0458_ _0640_/a_215_297# 0
C30545 hold55/a_391_47# net106 0.05785f
C30546 VPWR _1043_/a_381_47# 0.07717f
C30547 acc0.A\[9\] _0186_ 0.40055f
C30548 _0183_ acc0.A\[23\] 0.10439f
C30549 _0852_/a_35_297# _0263_ 0
C30550 _0309_ _0306_ 0.10031f
C30551 _0209_ net29 0.16644f
C30552 _0160_ _0468_ 0
C30553 hold63/a_49_47# hold63/a_285_47# 0.22264f
C30554 _1028_/a_466_413# _0350_ 0
C30555 _0398_ _0397_ 0.12486f
C30556 _1018_/a_1059_315# _0399_ 0
C30557 _1038_/a_634_159# _0175_ 0
C30558 _1043_/a_891_413# _1043_/a_975_413# 0.00851f
C30559 _1043_/a_27_47# net129 0.22002f
C30560 _1043_/a_381_47# _1043_/a_561_413# 0.00123f
C30561 net7 net174 0.75455f
C30562 _0446_ _0264_ 0.29024f
C30563 hold18/a_285_47# _0265_ 0.00154f
C30564 VPWR _1015_/a_634_159# 0.18309f
C30565 comp0.B\[13\] _0176_ 0.10587f
C30566 clknet_1_0__leaf__0464_ _0198_ 0
C30567 hold58/a_49_47# _1037_/a_891_413# 0
C30568 _0216_ _0599_/a_113_47# 0
C30569 net103 hold72/a_49_47# 0
C30570 _0195_ clknet_1_0__leaf__0461_ 0.25442f
C30571 _0554_/a_150_297# net24 0.0013f
C30572 _1034_/a_27_47# _1065_/a_27_47# 0
C30573 _0343_ _0398_ 0.0058f
C30574 _1050_/a_27_47# _0525_/a_299_297# 0
C30575 _0176_ _1046_/a_193_47# 0
C30576 _0283_ _0651_/a_113_47# 0.00998f
C30577 _1042_/a_27_47# net153 0
C30578 _1030_/a_1059_315# net208 0
C30579 _1030_/a_193_47# _0128_ 0.00378f
C30580 _0275_ _0819_/a_81_21# 0
C30581 _0371_ _0370_ 0.24198f
C30582 _1021_/a_27_47# net88 0.04493f
C30583 _1054_/a_634_159# _1054_/a_381_47# 0
C30584 _0786_/a_472_297# _0369_ 0.00112f
C30585 hold11/a_391_47# clkbuf_0__0464_/a_110_47# 0.00124f
C30586 _0363_ clknet_1_1__leaf__0460_ 0.0102f
C30587 _1071_/a_466_413# control0.count\[0\] 0
C30588 _1015_/a_634_159# _1015_/a_466_413# 0.23992f
C30589 _1015_/a_193_47# _1015_/a_1059_315# 0.03405f
C30590 _1015_/a_27_47# _1015_/a_891_413# 0.03224f
C30591 clknet_0__0458_ _0465_ 0.30155f
C30592 _0983_/a_891_413# VPWR 0.17957f
C30593 net123 net161 0
C30594 _0814_/a_181_47# _0181_ 0
C30595 net247 _0262_ 0
C30596 clknet_1_1__leaf__0462_ _1027_/a_466_413# 0.00607f
C30597 pp[27] _0108_ 0.00123f
C30598 net113 _1027_/a_193_47# 0.016f
C30599 _0311_ net52 0.00123f
C30600 _0792_/a_209_297# _0400_ 0.03812f
C30601 _0792_/a_209_47# _0405_ 0
C30602 _0989_/a_27_47# output63/a_27_47# 0
C30603 _1014_/a_27_47# _0585_/a_27_297# 0
C30604 _1020_/a_193_47# comp0.B\[0\] 0
C30605 _1053_/a_27_47# _0180_ 0
C30606 _1038_/a_634_159# _1038_/a_1059_315# 0
C30607 _1038_/a_27_47# _1038_/a_381_47# 0.06222f
C30608 _1038_/a_193_47# _1038_/a_891_413# 0.19322f
C30609 _0446_ net170 0
C30610 clknet_0__0465_ clkbuf_1_0__f__0465_/a_110_47# 0.31944f
C30611 _0319_ _1008_/a_634_159# 0
C30612 net53 _0323_ 0
C30613 _0307_ _0219_ 0.15333f
C30614 _1041_/a_1059_315# net173 0
C30615 _1041_/a_27_47# _0138_ 0
C30616 _0655_/a_215_53# _0655_/a_297_297# 0.00494f
C30617 A[6] input14/a_75_212# 0
C30618 input13/a_75_212# A[7] 0.00206f
C30619 net55 _0350_ 0.08014f
C30620 _0343_ _0277_ 0
C30621 control0.state\[0\] _1065_/a_466_413# 0
C30622 acc0.A\[12\] net142 0
C30623 acc0.A\[8\] _0987_/a_975_413# 0
C30624 _0637_/a_56_297# _0849_/a_79_21# 0.02101f
C30625 _0446_ _0845_/a_109_297# 0.01346f
C30626 net61 _0529_/a_109_297# 0
C30627 net162 _0344_ 0.03598f
C30628 _0461_ _0766_/a_109_297# 0
C30629 net214 hold67/a_49_47# 0
C30630 _0990_/a_193_47# acc0.A\[6\] 0
C30631 _0983_/a_634_159# _0983_/a_592_47# 0
C30632 clknet_1_0__leaf__0465_ _1051_/a_561_413# 0
C30633 _0527_/a_27_297# _0142_ 0.02024f
C30634 hold59/a_49_47# _0242_ 0
C30635 _0183_ hold60/a_49_47# 0.03068f
C30636 _0217_ hold60/a_391_47# 0.00161f
C30637 net157 control0.sh 0
C30638 clknet_1_0__leaf__0465_ _1045_/a_592_47# 0
C30639 _0261_ _0844_/a_79_21# 0.00605f
C30640 _0262_ _0844_/a_382_297# 0
C30641 pp[18] VPWR 0.31114f
C30642 net40 _0995_/a_466_413# 0.00393f
C30643 net245 _0995_/a_193_47# 0.05975f
C30644 net234 _0266_ 0.04631f
C30645 _0574_/a_27_297# _0574_/a_109_47# 0.00393f
C30646 clknet_0__0461_ _0246_ 0
C30647 net207 _0352_ 0
C30648 _0286_ _0806_/a_113_297# 0.00825f
C30649 _0449_ _0186_ 0.0012f
C30650 _0985_/a_1059_315# net71 0
C30651 _0201_ comp0.B\[12\] 0.09785f
C30652 output56/a_27_47# _0336_ 0
C30653 _0243_ VPWR 0.85692f
C30654 _0369_ net47 0.02282f
C30655 _1026_/a_891_413# _0320_ 0
C30656 hold50/a_49_47# _0345_ 0
C30657 clkbuf_1_1__f__0460_/a_110_47# _0320_ 0
C30658 net71 _1049_/a_193_47# 0
C30659 _1021_/a_1059_315# _0384_ 0
C30660 net219 hold72/a_285_47# 0.0113f
C30661 _0747_/a_79_21# _1006_/a_27_47# 0.01181f
C30662 _0437_ pp[5] 0.0032f
C30663 acc0.A\[27\] clknet_0__0462_ 0.00163f
C30664 _0459_ _0505_/a_109_47# 0
C30665 _0466_ _1068_/a_634_159# 0.02169f
C30666 _1056_/a_27_47# _0154_ 0.00631f
C30667 _0189_ net143 0
C30668 net90 _1007_/a_466_413# 0
C30669 _0637_/a_311_297# _0269_ 0.004f
C30670 _0831_/a_285_47# _0369_ 0
C30671 _1048_/a_27_47# _1047_/a_193_47# 0
C30672 _1048_/a_193_47# _1047_/a_27_47# 0
C30673 _1003_/a_561_413# _0217_ 0
C30674 _1003_/a_891_413# _0183_ 0.00309f
C30675 net132 net131 0
C30676 _0280_ _0644_/a_285_47# 0
C30677 _1004_/a_634_159# net50 0
C30678 _0852_/a_117_297# net47 0
C30679 _1013_/a_975_413# _0218_ 0
C30680 _0698_/a_199_47# _0322_ 0
C30681 _0698_/a_113_297# _0329_ 0.05986f
C30682 _0081_ clknet_1_0__leaf__0461_ 0.0018f
C30683 hold10/a_285_47# acc0.A\[15\] 0.05322f
C30684 _1016_/a_634_159# net166 0.00366f
C30685 _0244_ _0581_/a_109_47# 0.00338f
C30686 _0388_ _0581_/a_27_297# 0
C30687 _0346_ control0.add 0.5596f
C30688 output48/a_27_47# pp[20] 0.15855f
C30689 net211 _0242_ 0
C30690 VPWR net227 0.45454f
C30691 _0195_ net133 0
C30692 _0192_ _0180_ 0.01252f
C30693 hold11/a_285_47# net147 0
C30694 clknet_0__0464_ net7 0
C30695 net113 _1026_/a_1059_315# 0.03008f
C30696 _0998_/a_27_47# _0399_ 0.02361f
C30697 _0998_/a_193_47# _0398_ 0.02902f
C30698 _0681_/a_113_47# _0219_ 0
C30699 net49 _0382_ 0.00101f
C30700 _0176_ comp0.B\[9\] 0.27055f
C30701 _0300_ net5 0
C30702 hold17/a_49_47# VPWR 0.30785f
C30703 _0337_ hold61/a_49_47# 0.01272f
C30704 _0354_ _0568_/a_27_297# 0
C30705 net217 _0090_ 0.0617f
C30706 VPWR _0088_ 0.28784f
C30707 net85 _0096_ 0.00118f
C30708 net19 hold51/a_285_47# 0
C30709 _0343_ _0353_ 0.09971f
C30710 VPWR _0407_ 0.35204f
C30711 _0471_ _0951_/a_209_311# 0
C30712 clknet_0__0462_ _0364_ 0
C30713 _0559_/a_51_297# VPWR 0.46512f
C30714 _0577_/a_27_297# hold4/a_285_47# 0.00104f
C30715 _0514_/a_109_47# _0189_ 0
C30716 _0430_ _0086_ 0
C30717 net39 _0994_/a_975_413# 0
C30718 acc0.A\[26\] _1008_/a_1059_315# 0
C30719 _0479_ _0976_/a_505_21# 0
C30720 _0195_ _0585_/a_27_297# 0.01258f
C30721 _0234_ _0601_/a_68_297# 0
C30722 _1059_/a_592_47# acc0.A\[14\] 0
C30723 hold54/a_285_47# _0131_ 0
C30724 _0538_/a_512_297# _0142_ 0
C30725 hold42/a_391_47# acc0.A\[11\] 0.02877f
C30726 clknet_1_1__leaf__0459_ _1057_/a_1059_315# 0
C30727 net160 _1035_/a_193_47# 0
C30728 _0210_ _1035_/a_27_47# 0
C30729 _0780_/a_285_297# _0219_ 0
C30730 _1057_/a_891_413# acc0.A\[11\] 0.00302f
C30731 _0093_ acc0.A\[13\] 0
C30732 net103 clknet_0__0461_ 0.00352f
C30733 _0729_/a_68_297# _0332_ 0
C30734 comp0.B\[4\] _1034_/a_193_47# 0
C30735 _1036_/a_193_47# comp0.B\[2\] 0
C30736 _0378_ hold94/a_285_47# 0
C30737 net53 net237 0.00634f
C30738 _1052_/a_1059_315# net65 0
C30739 _0343_ _0298_ 0
C30740 hold76/a_391_47# _0183_ 0
C30741 _0343_ _0754_/a_240_47# 0
C30742 A[11] net3 0.14648f
C30743 _0356_ hold95/a_285_47# 0
C30744 VPWR input29/a_75_212# 0.27981f
C30745 _1056_/a_466_413# net182 0.0058f
C30746 hold29/a_49_47# net176 0
C30747 _0744_/a_27_47# _0090_ 0.00225f
C30748 hold18/a_285_47# _0267_ 0
C30749 _1004_/a_193_47# net215 0
C30750 input1/a_27_47# input26/a_75_212# 0
C30751 _0179_ _0989_/a_27_47# 0.00146f
C30752 _1054_/a_592_47# VPWR 0
C30753 net76 clkbuf_0__0465_/a_110_47# 0
C30754 _0179_ hold1/a_49_47# 0
C30755 _0643_/a_337_297# _0258_ 0
C30756 _0272_ _0626_/a_150_297# 0
C30757 _0734_/a_285_47# _1009_/a_27_47# 0
C30758 _0734_/a_47_47# _1009_/a_466_413# 0
C30759 _0618_/a_510_47# net52 0
C30760 VPWR _0569_/a_109_297# 0.21242f
C30761 _1051_/a_1017_47# net73 0
C30762 net63 _0519_/a_299_297# 0.00628f
C30763 _0179_ _0992_/a_27_47# 0
C30764 clknet_1_0__leaf__0459_ _1015_/a_634_159# 0
C30765 hold34/a_285_47# net181 0.01089f
C30766 _0163_ _1065_/a_1059_315# 0
C30767 _0243_ _0390_ 0.19578f
C30768 _1038_/a_975_413# VPWR 0.00439f
C30769 clkbuf_1_0__f__0458_/a_110_47# _0263_ 0.02638f
C30770 _0335_ _0705_/a_59_75# 0
C30771 output65/a_27_47# net63 0.01431f
C30772 _1041_/a_975_413# A[15] 0
C30773 hold45/a_285_47# _0188_ 0.00533f
C30774 output64/a_27_47# _0621_/a_35_297# 0
C30775 _1018_/a_1017_47# acc0.A\[18\] 0.00171f
C30776 net186 net23 0
C30777 _0731_/a_299_297# _0359_ 0.00208f
C30778 net35 _1072_/a_193_47# 0.00716f
C30779 hold57/a_285_47# _0553_/a_51_297# 0.01258f
C30780 _1067_/a_634_159# _0460_ 0
C30781 _1067_/a_1059_315# clknet_1_0__leaf__0457_ 0.021f
C30782 hold36/a_391_47# VPWR 0.1809f
C30783 hold87/a_285_47# _0637_/a_56_297# 0
C30784 _0519_/a_81_21# _0191_ 0.18194f
C30785 acc0.A\[8\] clkbuf_1_1__f__0458_/a_110_47# 0.00361f
C30786 _0983_/a_891_413# clknet_1_0__leaf__0459_ 0
C30787 _0816_/a_150_297# _0345_ 0
C30788 _0369_ _1060_/a_1059_315# 0
C30789 net219 _0392_ 0
C30790 _0209_ _0137_ 0
C30791 clknet_0__0463_ _0563_/a_149_47# 0.00374f
C30792 _1020_/a_27_47# net118 0.01147f
C30793 _0760_/a_47_47# _0760_/a_285_47# 0.01755f
C30794 _0557_/a_245_297# net27 0
C30795 clknet_1_0__leaf__0462_ _0313_ 0.25821f
C30796 hold101/a_285_47# _0218_ 0.03907f
C30797 _1031_/a_193_47# _1030_/a_1059_315# 0
C30798 _1031_/a_27_47# _1030_/a_891_413# 0
C30799 _1031_/a_466_413# _1030_/a_634_159# 0
C30800 net106 _0352_ 0
C30801 clknet_1_0__leaf__0464_ net247 0
C30802 _0457_ _1067_/a_634_159# 0.00101f
C30803 net35 _1071_/a_1017_47# 0
C30804 net51 _0103_ 0.34035f
C30805 _0404_ net5 0.26786f
C30806 _0507_/a_109_297# _0219_ 0.00716f
C30807 comp0.B\[14\] net31 0
C30808 _0180_ _0987_/a_891_413# 0
C30809 acc0.A\[5\] acc0.A\[4\] 0.1093f
C30810 _1038_/a_466_413# _0550_/a_240_47# 0
C30811 _0627_/a_109_93# _0465_ 0.01045f
C30812 hold7/a_49_47# net148 0.13679f
C30813 _0554_/a_68_297# _1037_/a_1059_315# 0.00211f
C30814 _1025_/a_634_159# _1025_/a_1059_315# 0
C30815 _1025_/a_27_47# _1025_/a_381_47# 0.06222f
C30816 _1025_/a_193_47# _1025_/a_891_413# 0.19497f
C30817 _0237_ _0352_ 0
C30818 _0354_ _0109_ 0.02751f
C30819 net122 net25 0
C30820 _0304_ acc0.A\[13\] 0
C30821 _1012_/a_466_413# _0345_ 0
C30822 _0770_/a_297_47# _0462_ 0.00108f
C30823 hold35/a_285_47# VPWR 0.2924f
C30824 hold82/a_49_47# _0219_ 0.00106f
C30825 _0573_/a_27_47# clknet_1_0__leaf__0461_ 0
C30826 comp0.B\[1\] _1032_/a_975_413# 0
C30827 _0413_ clknet_1_1__leaf__0459_ 0.13013f
C30828 net45 _0096_ 0.04463f
C30829 _0438_ acc0.A\[6\] 0.07063f
C30830 net58 _0627_/a_215_53# 0.01226f
C30831 input34/a_27_47# clknet_1_0__leaf_clk 0.00126f
C30832 _0180_ A[5] 0
C30833 _0113_ _0584_/a_27_297# 0.113f
C30834 _1055_/a_634_159# _0181_ 0
C30835 _0433_ _0172_ 0
C30836 net61 net170 0.00516f
C30837 hold28/a_391_47# _0195_ 0.02252f
C30838 net233 _0082_ 0
C30839 VPWR _0522_/a_373_47# 0
C30840 acc0.A\[12\] output66/a_27_47# 0.00104f
C30841 _1070_/a_634_159# _0466_ 0
C30842 _1070_/a_466_413# _0488_ 0
C30843 _0168_ _0976_/a_76_199# 0.02401f
C30844 VPWR _0976_/a_218_374# 0.00217f
C30845 _0243_ clknet_1_0__leaf__0459_ 0.02483f
C30846 _0324_ acc0.A\[25\] 0.17428f
C30847 _0800_/a_512_297# VPWR 0.00705f
C30848 _0352_ hold72/a_285_47# 0.00173f
C30849 net245 _0093_ 0.2531f
C30850 _0432_ _0271_ 0.39914f
C30851 net145 _0508_/a_81_21# 0.01165f
C30852 hold54/a_49_47# _1032_/a_27_47# 0
C30853 _0333_ _0219_ 0.23823f
C30854 _1046_/a_891_413# net10 0.06739f
C30855 clknet_0__0457_ _1001_/a_592_47# 0
C30856 _0118_ hold40/a_49_47# 0
C30857 net38 _0808_/a_81_21# 0
C30858 _0982_/a_27_47# _0856_/a_79_21# 0
C30859 _0238_ _0350_ 0.02514f
C30860 _1021_/a_27_47# _1067_/a_891_413# 0.00229f
C30861 hold17/a_49_47# hold17/a_285_47# 0.22264f
C30862 net191 acc0.A\[28\] 0.03442f
C30863 clknet_0__0463_ _1061_/a_27_47# 0
C30864 _0516_/a_27_297# _0990_/a_891_413# 0
C30865 net61 _0845_/a_109_297# 0
C30866 B[8] net127 0.00231f
C30867 _1003_/a_466_413# control0.state\[2\] 0
C30868 net85 _0395_ 0
C30869 _0473_ _0540_/a_51_297# 0.00142f
C30870 _0996_/a_634_159# _0996_/a_381_47# 0
C30871 _1055_/a_27_47# _0517_/a_81_21# 0.00171f
C30872 _0483_ control0.count\[1\] 0
C30873 clknet_0__0465_ _0824_/a_145_75# 0
C30874 net169 net9 0
C30875 _0769_/a_299_297# _0352_ 0.06981f
C30876 _0227_ _0222_ 0.27642f
C30877 net45 _1031_/a_193_47# 0
C30878 net31 _0543_/a_68_297# 0
C30879 VPWR _0835_/a_292_297# 0.00854f
C30880 _0209_ comp0.B\[6\] 0.21427f
C30881 _0728_/a_59_75# _0333_ 0.14964f
C30882 _0991_/a_27_47# _0268_ 0
C30883 _0955_/a_32_297# control0.sh 0
C30884 hold11/a_285_47# _0473_ 0
C30885 _0935_/a_27_47# clknet_1_1__leaf__0457_ 0.22795f
C30886 _0465_ clkbuf_1_1__f__0457_/a_110_47# 0.01486f
C30887 clknet_1_0__leaf__0464_ _1048_/a_466_413# 0
C30888 net133 _1048_/a_193_47# 0.00122f
C30889 clknet_1_1__leaf__0457_ _1061_/a_193_47# 0
C30890 _0793_/a_240_47# _0095_ 0.00137f
C30891 net46 net50 0.09546f
C30892 acc0.A\[16\] _1017_/a_1017_47# 0
C30893 _0469_ _0477_ 0
C30894 _0376_ _0754_/a_240_47# 0.01304f
C30895 _0343_ net36 0
C30896 _0732_/a_80_21# _0219_ 0.00932f
C30897 _0559_/a_51_297# _0559_/a_245_297# 0.01218f
C30898 hold8/a_391_47# _1027_/a_27_47# 0
C30899 net64 clkbuf_1_1__f__0458_/a_110_47# 0.02812f
C30900 _1057_/a_27_47# clknet_1_1__leaf__0465_ 0.0848f
C30901 VPWR _0996_/a_592_47# 0
C30902 net66 net3 0
C30903 _0317_ _1008_/a_466_413# 0
C30904 _1065_/a_592_47# comp0.B\[0\] 0
C30905 _0726_/a_240_47# acc0.A\[29\] 0
C30906 clkbuf_1_1__f__0463_/a_110_47# net24 0.00622f
C30907 net215 net199 0.21941f
C30908 control0.count\[3\] clknet_0_clk 0.02389f
C30909 acc0.A\[9\] net62 0
C30910 _1051_/a_381_47# _0149_ 0.11943f
C30911 hold22/a_285_47# _1054_/a_1059_315# 0.00197f
C30912 hold22/a_49_47# _1054_/a_891_413# 0.01135f
C30913 _1051_/a_466_413# acc0.A\[5\] 0
C30914 hold64/a_49_47# net47 0.00181f
C30915 _0803_/a_68_297# _0802_/a_59_75# 0.00101f
C30916 _0195_ _0218_ 0.43648f
C30917 _0274_ _0252_ 0.04195f
C30918 _0992_/a_381_47# acc0.A\[10\] 0.00129f
C30919 net67 _0508_/a_81_21# 0
C30920 _0287_ clkbuf_1_1__f__0465_/a_110_47# 0
C30921 _0805_/a_27_47# _0284_ 0
C30922 clkbuf_1_0__f__0460_/a_110_47# _0219_ 0.03601f
C30923 net62 _0986_/a_592_47# 0.00266f
C30924 net22 _1040_/a_891_413# 0
C30925 _0730_/a_215_47# clkbuf_1_1__f__0460_/a_110_47# 0.00234f
C30926 _0268_ _0350_ 0.02164f
C30927 _0169_ clknet_1_0__leaf_clk 0.00502f
C30928 _0480_ control0.count\[0\] 0.45984f
C30929 _0736_/a_56_297# VPWR 0.2571f
C30930 _0399_ _0990_/a_891_413# 0.03038f
C30931 _0787_/a_80_21# _0993_/a_466_413# 0
C30932 clknet_0__0458_ _0254_ 0.04822f
C30933 _0298_ A[14] 0
C30934 _1051_/a_1059_315# _0528_/a_81_21# 0
C30935 hold49/a_49_47# _0540_/a_51_297# 0
C30936 hold47/a_391_47# clknet_1_1__leaf__0464_ 0.01596f
C30937 _0250_ _0219_ 0.07268f
C30938 _0714_/a_149_47# net117 0
C30939 _0440_ hold1/a_285_47# 0
C30940 _0715_/a_27_47# _0424_ 0
C30941 _1002_/a_381_47# net240 0
C30942 _1039_/a_27_47# clknet_0__0463_ 0.03883f
C30943 _0369_ _0796_/a_510_47# 0
C30944 _1060_/a_634_159# net229 0
C30945 _0714_/a_51_297# _1013_/a_634_159# 0
C30946 _0090_ _0350_ 0
C30947 VPWR net208 0.28376f
C30948 acc0.A\[21\] _0385_ 0
C30949 _1003_/a_1059_315# _0467_ 0
C30950 _0644_/a_47_47# net41 0.05569f
C30951 _0924_/a_27_47# VPWR 0.20062f
C30952 clknet_0__0464_ _0202_ 0
C30953 acc0.A\[20\] _0217_ 0.04582f
C30954 _1030_/a_466_413# _0345_ 0
C30955 _1072_/a_27_47# net159 0
C30956 _0972_/a_93_21# _1062_/a_193_47# 0.00525f
C30957 _0972_/a_250_297# _1062_/a_27_47# 0.00135f
C30958 hold76/a_285_47# _1000_/a_27_47# 0
C30959 hold76/a_49_47# _1000_/a_193_47# 0
C30960 _0260_ _0186_ 0.00956f
C30961 clknet_1_0__leaf__0463_ _1040_/a_891_413# 0.00351f
C30962 hold67/a_391_47# _0428_ 0.00142f
C30963 hold3/a_391_47# _1005_/a_466_413# 0
C30964 net58 pp[1] 0
C30965 _0984_/a_193_47# net233 0
C30966 _1039_/a_193_47# clknet_1_1__leaf__0457_ 0
C30967 _1032_/a_193_47# _1032_/a_592_47# 0.00135f
C30968 _1032_/a_466_413# _1032_/a_561_413# 0.00772f
C30969 _1032_/a_634_159# _1032_/a_975_413# 0
C30970 _0294_ _0240_ 0.22937f
C30971 _1054_/a_891_413# net169 0.00121f
C30972 _1054_/a_381_47# net140 0
C30973 _0429_ output63/a_27_47# 0.0018f
C30974 _1015_/a_634_159# _0113_ 0.04214f
C30975 _0712_/a_79_21# _1030_/a_891_413# 0
C30976 _1038_/a_891_413# net29 0.00207f
C30977 _0294_ _0369_ 0.22031f
C30978 hold5/a_285_47# _0176_ 0
C30979 _0569_/a_27_297# _0569_/a_373_47# 0.01338f
C30980 _0649_/a_113_47# clknet_1_1__leaf__0459_ 0
C30981 hold31/a_49_47# _0186_ 0
C30982 hold14/a_49_47# net28 0
C30983 _0146_ net149 0.00649f
C30984 _1051_/a_634_159# _0180_ 0.0026f
C30985 hold33/a_391_47# net147 0
C30986 _0352_ _0392_ 0.05295f
C30987 clknet_1_1__leaf__0462_ net156 0.04319f
C30988 net224 VPWR 0.29871f
C30989 _0252_ pp[5] 0
C30990 _0820_/a_79_21# _0990_/a_27_47# 0
C30991 _0435_ _0827_/a_109_297# 0
C30992 _0343_ _1031_/a_1017_47# 0
C30993 _0126_ _0345_ 0
C30994 _1014_/a_27_47# _0112_ 0.10355f
C30995 _0852_/a_35_297# _0848_/a_27_47# 0
C30996 _1014_/a_891_413# net149 0.03526f
C30997 VPWR net180 0.4369f
C30998 _1038_/a_466_413# net172 0.00298f
C30999 _0600_/a_253_297# _0352_ 0.00107f
C31000 _0765_/a_79_21# hold3/a_285_47# 0
C31001 init _1066_/a_1059_315# 0
C31002 net33 _1066_/a_466_413# 0.03102f
C31003 net220 _0759_/a_113_47# 0
C31004 net234 _0399_ 0
C31005 hold46/a_285_47# clknet_1_1__leaf__0464_ 0
C31006 _0573_/a_27_47# _0585_/a_27_297# 0
C31007 _0852_/a_35_297# _0218_ 0
C31008 _0319_ net94 0
C31009 _1067_/a_592_47# clknet_1_0__leaf__0461_ 0
C31010 A[0] init 0.03345f
C31011 _0551_/a_27_47# _0533_/a_27_297# 0
C31012 hold75/a_49_47# VPWR 0.29426f
C31013 net45 _0395_ 0.00225f
C31014 _0290_ _0422_ 0.00664f
C31015 _0401_ net217 0.00296f
C31016 _0661_/a_277_297# _0345_ 0
C31017 _0637_/a_311_297# _0082_ 0
C31018 net46 _0399_ 0
C31019 net54 _0697_/a_80_21# 0
C31020 _0450_ _0449_ 0
C31021 clknet_1_0__leaf__0465_ _1044_/a_975_413# 0
C31022 comp0.B\[7\] _0472_ 0
C31023 _0536_/a_51_297# net7 0
C31024 _0665_/a_109_297# _0297_ 0.01129f
C31025 net126 _0176_ 0.06518f
C31026 hold16/a_285_47# _1030_/a_634_159# 0.00139f
C31027 _1020_/a_193_47# net1 0.02631f
C31028 hold16/a_391_47# _1030_/a_193_47# 0
C31029 _0287_ _0673_/a_253_47# 0.00376f
C31030 _0175_ _0494_/a_27_47# 0.00281f
C31031 net233 clkbuf_0__0458_/a_110_47# 0
C31032 _0997_/a_634_159# net43 0.04263f
C31033 hold58/a_49_47# net27 0.01236f
C31034 _0227_ _0762_/a_297_297# 0
C31035 net198 hold51/a_49_47# 0
C31036 _0454_ _0446_ 0
C31037 VPWR _0995_/a_193_47# 0.30688f
C31038 net72 _0444_ 0
C31039 net45 _0712_/a_297_297# 0.00242f
C31040 acc0.A\[8\] _0291_ 0.05333f
C31041 _0081_ _0218_ 0
C31042 _0131_ _0562_/a_68_297# 0
C31043 _1056_/a_27_47# _0820_/a_79_21# 0
C31044 input21/a_75_212# B[13] 0.19513f
C31045 _0347_ _0986_/a_193_47# 0
C31046 _0347_ acc0.A\[25\] 0.0288f
C31047 hold45/a_391_47# _0187_ 0.00655f
C31048 _0997_/a_975_413# net42 0
C31049 _0230_ _0223_ 0.18292f
C31050 _0240_ _0775_/a_297_297# 0
C31051 net197 _1008_/a_466_413# 0
C31052 _0104_ _1006_/a_193_47# 0.20033f
C31053 net216 _1006_/a_1059_315# 0.00506f
C31054 _0354_ _0725_/a_80_21# 0.00381f
C31055 net106 _1032_/a_891_413# 0
C31056 acc0.A\[12\] _1058_/a_381_47# 0.01693f
C31057 _0488_ _0166_ 0
C31058 net90 _0105_ 0
C31059 hold32/a_391_47# _1055_/a_466_413# 0.00388f
C31060 hold32/a_49_47# _1055_/a_891_413# 0.00386f
C31061 hold32/a_285_47# _1055_/a_1059_315# 0.00108f
C31062 hold31/a_285_47# _0253_ 0.05644f
C31063 acc0.A\[12\] _0420_ 0
C31064 _1000_/a_634_159# _0461_ 0.0049f
C31065 _0186_ _0524_/a_27_297# 0.14905f
C31066 _0954_/a_304_297# comp0.B\[10\] 0
C31067 net168 net148 0.00248f
C31068 _0174_ net28 0.00102f
C31069 _0578_/a_373_47# _0352_ 0
C31070 _1061_/a_592_47# acc0.A\[15\] 0
C31071 _0546_/a_51_297# _0546_/a_512_297# 0.0116f
C31072 _0616_/a_215_47# _0246_ 0.13642f
C31073 clknet_0__0461_ _0774_/a_68_297# 0
C31074 _1036_/a_1059_315# _0175_ 0.03188f
C31075 _0163_ hold93/a_49_47# 0
C31076 _0181_ hold93/a_391_47# 0.05394f
C31077 hold101/a_49_47# net63 0.29353f
C31078 _0534_/a_81_21# _0180_ 0.00379f
C31079 _0534_/a_299_297# _0182_ 0
C31080 clknet_1_1__leaf__0462_ acc0.A\[26\] 0.04568f
C31081 _0991_/a_27_47# _0991_/a_466_413# 0.27314f
C31082 _0991_/a_193_47# _0991_/a_634_159# 0.12388f
C31083 _0534_/a_81_21# net218 0.00165f
C31084 VPWR _0516_/a_109_297# 0.19464f
C31085 _0366_ hold90/a_285_47# 0
C31086 _0315_ hold90/a_49_47# 0.02055f
C31087 clknet_1_0__leaf__0465_ _0180_ 0.05485f
C31088 net158 clknet_1_0__leaf__0464_ 0
C31089 _0356_ _1011_/a_193_47# 0
C31090 _0397_ _0308_ 0.10377f
C31091 _0241_ _0771_/a_298_297# 0.00886f
C31092 _0839_/a_109_297# _0268_ 0
C31093 hold23/a_391_47# _0180_ 0.05045f
C31094 _1041_/a_27_47# net22 0
C31095 net215 VPWR 0.30861f
C31096 _0120_ hold4/a_285_47# 0.03234f
C31097 _0210_ _0957_/a_114_297# 0
C31098 net160 _0957_/a_220_297# 0
C31099 acc0.A\[20\] _0248_ 0.00249f
C31100 _0195_ _0112_ 0
C31101 _0479_ _0466_ 0.02904f
C31102 hold46/a_49_47# net7 0
C31103 net70 _0450_ 0
C31104 clknet_1_1__leaf__0460_ acc0.A\[23\] 0
C31105 _0539_/a_68_297# B[11] 0
C31106 _0982_/a_466_413# _1014_/a_891_413# 0
C31107 _0833_/a_297_297# _0369_ 0.00431f
C31108 _0143_ _0142_ 0.02023f
C31109 _0195_ _1017_/a_975_413# 0
C31110 net104 _0345_ 0
C31111 _0179_ net11 0.20201f
C31112 _1001_/a_193_47# _0217_ 0.03897f
C31113 clkbuf_1_1__f__0462_/a_110_47# _0686_/a_27_53# 0.00586f
C31114 _0429_ _0179_ 0.00419f
C31115 hold6/a_49_47# _1040_/a_193_47# 0
C31116 hold6/a_285_47# _1040_/a_27_47# 0
C31117 _0100_ acc0.A\[21\] 0.00774f
C31118 hold39/a_285_47# _0132_ 0.00464f
C31119 _0399_ _0996_/a_27_47# 0.03263f
C31120 _0398_ _0996_/a_193_47# 0
C31121 net186 _0213_ 0
C31122 _0209_ net26 0
C31123 _0375_ clknet_1_0__leaf__0460_ 0.08809f
C31124 _1057_/a_975_413# VPWR 0.00464f
C31125 clknet_1_0__leaf__0465_ _0432_ 0.00101f
C31126 _0651_/a_113_47# _0345_ 0
C31127 _1048_/a_975_413# _0186_ 0
C31128 clkbuf_1_1__f__0462_/a_110_47# _1008_/a_891_413# 0
C31129 hold54/a_49_47# hold54/a_285_47# 0.22264f
C31130 _0579_/a_109_47# VPWR 0
C31131 hold35/a_285_47# hold35/a_391_47# 0.41909f
C31132 _1041_/a_27_47# clknet_1_0__leaf__0463_ 0.045f
C31133 hold13/a_391_47# hold57/a_285_47# 0.00144f
C31134 _0174_ _0540_/a_512_297# 0.00318f
C31135 _1058_/a_27_47# acc0.A\[10\] 0.00458f
C31136 _0296_ _0282_ 0
C31137 _0687_/a_59_75# _0364_ 0
C31138 _1067_/a_27_47# _0161_ 0
C31139 net64 _0291_ 0
C31140 _0446_ _0846_/a_51_297# 0.01542f
C31141 net53 _0320_ 0.00343f
C31142 _0181_ control0.reset 0
C31143 VPWR _0096_ 0.46068f
C31144 _0343_ pp[15] 0.27296f
C31145 _0850_/a_68_297# acc0.A\[0\] 0
C31146 _0404_ _0303_ 0
C31147 _0522_/a_109_297# acc0.A\[6\] 0.01903f
C31148 hold65/a_285_47# _0434_ 0
C31149 _0722_/a_215_47# _0347_ 0.06498f
C31150 _0257_ _0441_ 0.00544f
C31151 net28 _0208_ 0.23595f
C31152 _0800_/a_245_297# _0800_/a_240_47# 0
C31153 net61 _0856_/a_79_21# 0
C31154 _0333_ hold61/a_49_47# 0.00111f
C31155 acc0.A\[29\] _0568_/a_109_47# 0
C31156 _0476_ _0468_ 0.37222f
C31157 hold87/a_391_47# _0269_ 0
C31158 _0290_ acc0.A\[8\] 0.08799f
C31159 _0401_ net66 0
C31160 _0423_ _0291_ 0
C31161 _1017_/a_561_413# _0369_ 0
C31162 _0398_ clkbuf_0__0461_/a_110_47# 0
C31163 net236 _0479_ 0
C31164 _0225_ _1023_/a_891_413# 0
C31165 net54 _0345_ 0.09052f
C31166 _1002_/a_634_159# _0352_ 0
C31167 net44 _1031_/a_891_413# 0
C31168 _0183_ _0263_ 0
C31169 _0490_ _1068_/a_27_47# 0
C31170 _0183_ clkload4/Y 0
C31171 VPWR _0545_/a_150_297# 0.00148f
C31172 _0996_/a_193_47# _0277_ 0
C31173 VPWR _0695_/a_80_21# 0.25325f
C31174 _0179_ hold7/a_391_47# 0.05295f
C31175 _0627_/a_109_93# _0254_ 0.06129f
C31176 _1004_/a_27_47# net52 0.0429f
C31177 hold85/a_49_47# _0972_/a_93_21# 0
C31178 VPWR _1031_/a_193_47# 0.31098f
C31179 clkbuf_0__0465_/a_110_47# _0986_/a_193_47# 0.01012f
C31180 clkbuf_1_0__f__0461_/a_110_47# _0350_ 0
C31181 hold31/a_285_47# net74 0.00889f
C31182 hold9/a_391_47# _0364_ 0
C31183 _0216_ _0391_ 0.03046f
C31184 _0183_ _0582_/a_373_47# 0.00279f
C31185 _0731_/a_299_297# _0238_ 0
C31186 _0290_ _0991_/a_193_47# 0
C31187 _0401_ _0991_/a_27_47# 0
C31188 _1012_/a_381_47# _0308_ 0
C31189 _0749_/a_299_297# _0460_ 0.00998f
C31190 pp[23] _1022_/a_1059_315# 0
C31191 _0404_ _0281_ 0
C31192 hold26/a_285_47# VPWR 0.29294f
C31193 _0345_ _0806_/a_199_47# 0
C31194 comp0.B\[14\] net7 0
C31195 clkbuf_1_0__f__0458_/a_110_47# _0848_/a_27_47# 0
C31196 _1057_/a_891_413# A[12] 0
C31197 _0835_/a_78_199# _0835_/a_215_47# 0.09071f
C31198 clknet_1_0__leaf__0464_ net148 0
C31199 hold76/a_285_47# acc0.A\[19\] 0.00179f
C31200 hold35/a_285_47# net182 0.01139f
C31201 _1038_/a_891_413# _0137_ 0
C31202 _1038_/a_561_413# _0172_ 0
C31203 _1004_/a_193_47# clknet_1_0__leaf__0460_ 0.00213f
C31204 clkbuf_1_0__f__0458_/a_110_47# _0218_ 0.01746f
C31205 hold23/a_285_47# net10 0.06796f
C31206 hold25/a_391_47# net153 0
C31207 hold78/a_391_47# net60 0.00778f
C31208 clknet_1_1__leaf__0463_ comp0.B\[15\] 0
C31209 _0216_ _0581_/a_27_297# 0
C31210 net47 _0084_ 0
C31211 _1025_/a_27_47# acc0.A\[25\] 0.05281f
C31212 net49 net91 0.25027f
C31213 _0430_ _0350_ 0
C31214 _0984_/a_891_413# _0347_ 0.01003f
C31215 _1030_/a_1059_315# _0221_ 0
C31216 _0971_/a_81_21# _0880_/a_27_47# 0
C31217 hold72/a_49_47# hold72/a_391_47# 0.00188f
C31218 hold36/a_285_47# _0172_ 0.00684f
C31219 hold89/a_285_47# _0468_ 0.00181f
C31220 hold65/a_391_47# net65 0.0796f
C31221 _0982_/a_975_413# _0195_ 0
C31222 hold65/a_285_47# _0989_/a_1059_315# 0.00319f
C31223 clknet_1_0__leaf__0462_ _0321_ 0
C31224 _0168_ _0488_ 0.00961f
C31225 _1001_/a_634_159# control0.add 0
C31226 _0093_ VPWR 0.31489f
C31227 acc0.A\[12\] _0284_ 0
C31228 net67 net143 0
C31229 clkbuf_1_0__f__0457_/a_110_47# _1019_/a_193_47# 0
C31230 _0401_ _0350_ 0
C31231 clknet_1_0__leaf__0462_ clkbuf_0__0460_/a_110_47# 0
C31232 _0211_ _0173_ 0.1583f
C31233 _0559_/a_51_297# comp0.B\[3\] 0
C31234 comp0.B\[5\] _0215_ 0.00128f
C31235 VPWR net71 0.40564f
C31236 acc0.A\[11\] _0419_ 0
C31237 hold22/a_49_47# hold22/a_391_47# 0.00188f
C31238 _0190_ _0990_/a_891_413# 0
C31239 net8 comp0.B\[15\] 0.03448f
C31240 _0263_ acc0.A\[15\] 0.10892f
C31241 clkload4/Y acc0.A\[15\] 0
C31242 _0101_ control0.state\[2\] 0
C31243 net89 _0486_ 0.00226f
C31244 VPWR _0808_/a_368_297# 0.00127f
C31245 _1055_/a_466_413# _0153_ 0
C31246 _0366_ clknet_0__0462_ 0.00193f
C31247 net217 hold70/a_49_47# 0
C31248 _0218_ _0779_/a_510_47# 0.00466f
C31249 _0357_ _0332_ 0.24076f
C31250 hold77/a_391_47# VPWR 0.18492f
C31251 _1047_/a_27_47# acc0.A\[15\] 0
C31252 _0769_/a_81_21# _0769_/a_384_47# 0.00138f
C31253 net64 _0621_/a_285_297# 0.06422f
C31254 _0621_/a_35_297# _0621_/a_285_47# 0.00723f
C31255 _0233_ acc0.A\[23\] 0.01896f
C31256 clknet_0__0458_ _0625_/a_59_75# 0
C31257 _0268_ _0847_/a_109_297# 0.00224f
C31258 net222 _0350_ 0.133f
C31259 _0474_ control0.sh 0
C31260 _0183_ clknet_1_0__leaf__0461_ 0.24274f
C31261 _0575_/a_109_297# acc0.A\[23\] 0
C31262 _0153_ net181 0
C31263 _0123_ _0216_ 0.05182f
C31264 hold87/a_49_47# hold87/a_391_47# 0.00188f
C31265 hold86/a_49_47# net247 0.00125f
C31266 hold30/a_49_47# _0222_ 0
C31267 _0714_/a_240_47# _0342_ 0.01304f
C31268 acc0.A\[16\] _1016_/a_381_47# 0
C31269 _0200_ _0540_/a_51_297# 0
C31270 _0330_ _0318_ 0
C31271 clknet_1_0__leaf__0463_ _1039_/a_975_413# 0
C31272 VPWR _1036_/a_1017_47# 0
C31273 A[13] pp[13] 0.18126f
C31274 input7/a_75_212# net153 0
C31275 _0179_ clknet_1_1__leaf__0458_ 0.44808f
C31276 _0437_ _0828_/a_113_297# 0
C31277 net98 _0394_ 0
C31278 _1059_/a_27_47# clkbuf_0__0459_/a_110_47# 0.00876f
C31279 _1044_/a_634_159# _1044_/a_592_47# 0
C31280 _0178_ _1048_/a_27_47# 0
C31281 _1065_/a_634_159# _0564_/a_68_297# 0
C31282 comp0.B\[13\] _0954_/a_114_297# 0.00111f
C31283 hold11/a_285_47# _0200_ 0
C31284 net158 _0536_/a_245_297# 0
C31285 _1038_/a_891_413# comp0.B\[6\] 0.04016f
C31286 hold52/a_49_47# net199 0.00335f
C31287 hold41/a_49_47# _1058_/a_1059_315# 0.0045f
C31288 comp0.B\[8\] _0540_/a_51_297# 0
C31289 _0423_ _0290_ 0.72393f
C31290 _0149_ acc0.A\[5\] 0
C31291 hold22/a_391_47# net169 0.13101f
C31292 _0985_/a_27_47# _0465_ 0
C31293 _0971_/a_81_21# _1062_/a_27_47# 0
C31294 VPWR _0743_/a_512_297# 0.00834f
C31295 _1058_/a_27_47# _0510_/a_109_297# 0
C31296 _0441_ net11 0
C31297 _0222_ _0352_ 0.04133f
C31298 _0512_/a_373_47# net67 0
C31299 clknet_1_1__leaf_clk _1065_/a_634_159# 0.03627f
C31300 net36 _1038_/a_27_47# 0.06294f
C31301 _0226_ _0384_ 0.01304f
C31302 VPWR _0395_ 0.32827f
C31303 _0182_ _0350_ 0
C31304 _0999_/a_466_413# _0778_/a_68_297# 0.00652f
C31305 _0353_ _0568_/a_27_297# 0
C31306 _0329_ _0726_/a_51_297# 0
C31307 _0985_/a_891_413# _0629_/a_59_75# 0
C31308 _0985_/a_27_47# acc0.A\[2\] 0.00239f
C31309 _0819_/a_299_297# _0990_/a_634_159# 0
C31310 _0461_ _0242_ 0.05165f
C31311 _0237_ _1005_/a_27_47# 0
C31312 VPWR input26/a_75_212# 0.26807f
C31313 _0260_ net62 0.07061f
C31314 _1067_/a_381_47# net17 0.01253f
C31315 net46 _1023_/a_592_47# 0
C31316 _0195_ _1028_/a_466_413# 0.03272f
C31317 _0216_ _1028_/a_193_47# 0
C31318 net56 net227 0
C31319 pp[8] acc0.A\[10\] 0
C31320 _0835_/a_78_199# _0172_ 0.01506f
C31321 net203 clknet_1_1__leaf__0463_ 0.06852f
C31322 hold49/a_285_47# net20 0.04185f
C31323 _0260_ _0450_ 0
C31324 _1057_/a_634_159# _1057_/a_1059_315# 0
C31325 _1057_/a_27_47# _1057_/a_381_47# 0.06222f
C31326 _1057_/a_193_47# _1057_/a_891_413# 0.19489f
C31327 hold48/a_285_47# hold49/a_285_47# 0
C31328 _0579_/a_27_297# net87 0.06211f
C31329 pp[17] _0712_/a_465_47# 0
C31330 _0111_ _1013_/a_27_47# 0.09948f
C31331 net225 _1013_/a_634_159# 0.01176f
C31332 hold81/a_391_47# _0419_ 0
C31333 net146 net229 0
C31334 VPWR _1064_/a_634_159# 0.19394f
C31335 clknet_0__0463_ _0953_/a_32_297# 0.00782f
C31336 _0800_/a_240_47# _0995_/a_27_47# 0
C31337 _1059_/a_193_47# _1059_/a_891_413# 0.19489f
C31338 _1059_/a_27_47# _1059_/a_381_47# 0.06222f
C31339 _1059_/a_634_159# _1059_/a_1059_315# 0
C31340 VPWR _0304_ 0.29721f
C31341 _0343_ _0428_ 0.02401f
C31342 _0712_/a_297_297# VPWR 0.27507f
C31343 _0179_ _0263_ 0.01991f
C31344 _0164_ _1062_/a_27_47# 0
C31345 net231 _1062_/a_193_47# 0.01504f
C31346 _0269_ _0264_ 0
C31347 hold96/a_391_47# _0123_ 0
C31348 _0849_/a_297_297# _0082_ 0
C31349 clknet_1_0__leaf__0461_ acc0.A\[15\] 0
C31350 _1015_/a_634_159# _0345_ 0
C31351 acc0.A\[14\] net247 0
C31352 pp[15] A[14] 0
C31353 _0443_ _0350_ 0
C31354 _0179_ _1047_/a_27_47# 0.00119f
C31355 clknet_1_0__leaf__0459_ _0096_ 0
C31356 _0221_ _0726_/a_51_297# 0
C31357 _1057_/a_975_413# _0283_ 0
C31358 hold37/a_285_47# clknet_1_1__leaf__0464_ 0.01843f
C31359 _0569_/a_373_47# _0127_ 0.00133f
C31360 _1065_/a_466_413# clkbuf_1_1__f_clk/a_110_47# 0.00231f
C31361 acc0.A\[20\] _0235_ 0.03159f
C31362 _0481_ _0978_/a_109_47# 0.00167f
C31363 _0179_ _1058_/a_891_413# 0
C31364 net137 _0180_ 0.00733f
C31365 net193 _0540_/a_51_297# 0.07959f
C31366 net214 _0990_/a_1059_315# 0
C31367 _0983_/a_193_47# _0219_ 0
C31368 _0388_ _0773_/a_285_47# 0
C31369 net186 _0161_ 0
C31370 _0310_ _0245_ 0
C31371 _0783_/a_215_47# _0398_ 0.01156f
C31372 _0783_/a_79_21# _0096_ 0.05023f
C31373 _0573_/a_27_47# _0112_ 0.00123f
C31374 _0718_/a_285_47# _0336_ 0.00119f
C31375 _0349_ _0705_/a_59_75# 0
C31376 _0328_ _0319_ 0.0426f
C31377 net220 _0352_ 0.06393f
C31378 net61 _0846_/a_51_297# 0.00259f
C31379 hold86/a_285_47# _0846_/a_240_47# 0
C31380 _0551_/a_27_47# _0199_ 0
C31381 net55 _0195_ 0.13273f
C31382 acc0.A\[27\] _1028_/a_561_413# 0
C31383 comp0.B\[14\] comp0.B\[11\] 0.00116f
C31384 net40 _0994_/a_193_47# 0
C31385 _0478_ _1069_/a_891_413# 0
C31386 _0960_/a_109_47# clknet_1_0__leaf_clk 0
C31387 hold38/a_391_47# _1062_/a_27_47# 0
C31388 hold100/a_285_47# _0447_ 0
C31389 net120 net23 0
C31390 clknet_0__0461_ hold72/a_391_47# 0.00205f
C31391 _0269_ net170 0
C31392 hold17/a_391_47# _0466_ 0.06419f
C31393 clknet_1_1__leaf__0460_ clknet_1_1__leaf__0462_ 0.11038f
C31394 net57 _0347_ 0
C31395 _1052_/a_466_413# _0186_ 0
C31396 _0343_ _0715_/a_27_47# 0.21364f
C31397 _0836_/a_150_297# _0433_ 0.00159f
C31398 _0267_ _0445_ 0
C31399 _0352_ _1006_/a_592_47# 0
C31400 _0570_/a_373_47# net113 0
C31401 net101 _1015_/a_381_47# 0
C31402 net186 _1033_/a_466_413# 0
C31403 _1058_/a_27_47# _0188_ 0
C31404 net69 acc0.A\[18\] 0
C31405 _0244_ clkbuf_1_0__f__0461_/a_110_47# 0.03662f
C31406 net45 _0344_ 0.00132f
C31407 clkbuf_1_1__f__0464_/a_110_47# _0194_ 0
C31408 _0433_ _0437_ 0
C31409 clkload1/a_110_47# VPWR 0
C31410 hold22/a_49_47# _0255_ 0
C31411 _0972_/a_93_21# net17 0.06603f
C31412 clkbuf_1_0__f__0464_/a_110_47# _1048_/a_466_413# 0
C31413 acc0.A\[25\] _0106_ 0
C31414 _0305_ _1060_/a_193_47# 0
C31415 _0217_ _0585_/a_109_47# 0
C31416 net38 _0652_/a_109_297# 0.00207f
C31417 _0399_ _0794_/a_27_47# 0.01093f
C31418 _1014_/a_466_413# clkbuf_0__0457_/a_110_47# 0
C31419 VPWR _0619_/a_150_297# 0.00137f
C31420 _0280_ _0302_ 0
C31421 _0216_ net216 0.00344f
C31422 hold39/a_285_47# _0477_ 0
C31423 net180 net30 0.10314f
C31424 clknet_0__0462_ _0689_/a_68_297# 0
C31425 comp0.B\[11\] _0543_/a_68_297# 0
C31426 _0243_ _0345_ 0
C31427 hold43/a_285_47# _0126_ 0
C31428 _0533_/a_27_297# _0199_ 0.168f
C31429 _0533_/a_373_47# _0180_ 0
C31430 _0109_ _0353_ 0
C31431 net35 control0.state\[2\] 0.00456f
C31432 hold66/a_49_47# net51 0.00167f
C31433 _0349_ _0358_ 0
C31434 _0183_ _1060_/a_891_413# 0.00191f
C31435 net45 _0709_/a_113_47# 0
C31436 acc0.A\[24\] _1007_/a_561_413# 0
C31437 hold71/a_391_47# net218 0.13134f
C31438 _0555_/a_245_297# net28 0
C31439 hold32/a_391_47# net179 0.1316f
C31440 net140 _0193_ 0
C31441 hold87/a_49_47# _0264_ 0
C31442 clkbuf_0__0463_/a_110_47# _0560_/a_68_297# 0.00104f
C31443 net86 _0461_ 0.0687f
C31444 _0123_ _1024_/a_193_47# 0
C31445 clknet_1_0__leaf__0462_ _1022_/a_193_47# 0.02078f
C31446 _0186_ _0194_ 0.04494f
C31447 net11 hold83/a_49_47# 0
C31448 _0978_/a_27_297# _0484_ 0
C31449 _0369_ hold3/a_49_47# 0
C31450 _0133_ clknet_0__0463_ 0.07301f
C31451 _0375_ hold94/a_285_47# 0
C31452 _0762_/a_297_297# _0352_ 0
C31453 hold38/a_391_47# _0133_ 0.00146f
C31454 _0546_/a_51_297# _0139_ 0.10369f
C31455 _0546_/a_240_47# net152 0.04192f
C31456 hold75/a_49_47# hold75/a_285_47# 0.22264f
C31457 VPWR _1023_/a_1017_47# 0
C31458 _1047_/a_466_413# clknet_1_1__leaf__0457_ 0
C31459 control0.state\[1\] _0974_/a_79_199# 0
C31460 _0230_ _0216_ 0
C31461 net149 _0580_/a_27_297# 0.05102f
C31462 _0991_/a_27_47# _0089_ 0.09323f
C31463 _0991_/a_193_47# net77 0.00544f
C31464 _0991_/a_1059_315# _0991_/a_1017_47# 0
C31465 _0210_ _0173_ 0.08727f
C31466 _0992_/a_561_413# _0187_ 0
C31467 comp0.B\[14\] _0202_ 0.05627f
C31468 net133 acc0.A\[15\] 0.05947f
C31469 _1067_/a_193_47# _0487_ 0
C31470 net227 _0345_ 0
C31471 pp[0] VPWR 0.37565f
C31472 _0125_ _0347_ 0
C31473 acc0.A\[27\] _0352_ 0
C31474 _0441_ clknet_1_1__leaf__0458_ 0
C31475 _0722_/a_79_21# net209 0
C31476 _0370_ _1006_/a_1059_315# 0
C31477 net78 hold70/a_391_47# 0
C31478 _1043_/a_193_47# _0541_/a_68_297# 0
C31479 _0803_/a_68_297# _0414_ 0.00125f
C31480 _0817_/a_81_21# _0294_ 0.00623f
C31481 _0371_ _0369_ 0
C31482 _0814_/a_181_47# clknet_1_1__leaf__0465_ 0
C31483 net97 net191 0
C31484 _0216_ _1029_/a_561_413# 0
C31485 hold52/a_49_47# VPWR 0.36442f
C31486 clknet_1_1__leaf__0459_ _0992_/a_27_47# 0.03546f
C31487 _0344_ _0587_/a_27_47# 0
C31488 _0730_/a_79_21# _0317_ 0
C31489 _0460_ hold73/a_49_47# 0
C31490 clknet_1_0__leaf__0457_ hold73/a_391_47# 0.00843f
C31491 clknet_1_1__leaf__0460_ net242 0
C31492 _0080_ _1014_/a_891_413# 0
C31493 _0982_/a_634_159# acc0.A\[0\] 0
C31494 _0982_/a_381_47# net100 0
C31495 _0793_/a_240_47# _0219_ 0.02361f
C31496 _0407_ _0345_ 0.26586f
C31497 net245 _0997_/a_27_47# 0
C31498 _1004_/a_891_413# acc0.A\[23\] 0.00292f
C31499 _0174_ _0542_/a_51_297# 0.08913f
C31500 VPWR _1065_/a_466_413# 0.24446f
C31501 _0600_/a_103_199# _0600_/a_337_297# 0.01015f
C31502 hold64/a_285_47# _0391_ 0
C31503 net123 _1037_/a_381_47# 0.00201f
C31504 net69 hold59/a_49_47# 0
C31505 _0725_/a_209_47# acc0.A\[29\] 0.00144f
C31506 _0995_/a_27_47# _0995_/a_466_413# 0.27314f
C31507 _0995_/a_193_47# _0995_/a_634_159# 0.12729f
C31508 _0197_ _0465_ 0.00134f
C31509 _0412_ _0297_ 0.00489f
C31510 _0357_ _0701_/a_209_47# 0.0035f
C31511 _0226_ _0383_ 0.22772f
C31512 _0739_/a_215_47# _0364_ 0.05011f
C31513 _0417_ _0418_ 0.15579f
C31514 _0419_ _0281_ 0.42662f
C31515 _0543_/a_68_297# _0202_ 0.0193f
C31516 _1021_/a_592_47# _0217_ 0
C31517 _0089_ _0350_ 0
C31518 _0352_ _0364_ 0.00236f
C31519 _1060_/a_891_413# acc0.A\[15\] 0.00352f
C31520 _0174_ _0142_ 0.0343f
C31521 clknet_0__0458_ _0273_ 0
C31522 acc0.A\[2\] _0197_ 0.31873f
C31523 control0.count\[3\] hold12/a_285_47# 0
C31524 _0681_/a_113_47# _0328_ 0
C31525 hold9/a_49_47# _1027_/a_193_47# 0.00127f
C31526 hold9/a_285_47# _1027_/a_27_47# 0.01366f
C31527 _1050_/a_27_47# _0142_ 0.0011f
C31528 hold57/a_391_47# _0555_/a_149_47# 0
C31529 net53 _1007_/a_1059_315# 0.13027f
C31530 _1070_/a_1059_315# _1069_/a_634_159# 0
C31531 _1070_/a_891_413# _1069_/a_193_47# 0.0047f
C31532 _1070_/a_634_159# _1069_/a_1059_315# 0
C31533 _1070_/a_193_47# _1069_/a_891_413# 0.0047f
C31534 _0110_ _0352_ 0.03605f
C31535 net34 _1062_/a_27_47# 0
C31536 control0.state\[0\] _1062_/a_634_159# 0.00537f
C31537 control0.state\[1\] _1062_/a_193_47# 0.02535f
C31538 _0976_/a_439_47# _0488_ 0.00571f
C31539 _0217_ _0208_ 0
C31540 net46 _0576_/a_27_297# 0.00429f
C31541 net39 A[13] 0
C31542 _0280_ net6 0
C31543 _0733_/a_448_47# _0328_ 0.00878f
C31544 net16 A[12] 0
C31545 _0285_ _0179_ 0.0023f
C31546 hold74/a_391_47# net221 0.13051f
C31547 VPWR _0329_ 1.68119f
C31548 net88 _0352_ 0.00281f
C31549 net201 _0214_ 0.09101f
C31550 _0180_ _0529_/a_373_47# 0.00122f
C31551 _1011_/a_634_159# _1011_/a_1059_315# 0
C31552 _1011_/a_27_47# _1011_/a_381_47# 0.05761f
C31553 _1011_/a_193_47# _1011_/a_891_413# 0.19489f
C31554 _1016_/a_466_413# _0369_ 0
C31555 net50 _1023_/a_193_47# 0.00768f
C31556 _0643_/a_103_199# net62 0.04708f
C31557 _0179_ net133 0.12129f
C31558 hold10/a_285_47# _0171_ 0.01545f
C31559 VPWR clknet_1_0__leaf__0460_ 4.13775f
C31560 pp[27] hold62/a_391_47# 0.00157f
C31561 hold29/a_49_47# net177 0.00378f
C31562 pp[9] hold34/a_391_47# 0.02822f
C31563 _0350_ _1006_/a_891_413# 0.03515f
C31564 acc0.A\[22\] net51 0.38833f
C31565 _0295_ _0286_ 0
C31566 clknet_0__0465_ _0986_/a_561_413# 0
C31567 _0304_ _0283_ 0
C31568 net102 acc0.A\[18\] 0
C31569 net45 _0997_/a_27_47# 0.00219f
C31570 _0618_/a_297_297# _0460_ 0
C31571 _0714_/a_149_47# _0216_ 0
C31572 net39 _0279_ 0.44718f
C31573 VPWR hold51/a_391_47# 0.18992f
C31574 _0130_ _1067_/a_634_159# 0
C31575 _1021_/a_193_47# hold73/a_391_47# 0
C31576 net210 _1025_/a_27_47# 0.0011f
C31577 net56 net208 0
C31578 _0350_ _0986_/a_891_413# 0.01778f
C31579 _1020_/a_381_47# VPWR 0.07811f
C31580 _1001_/a_466_413# _0610_/a_59_75# 0
C31581 net214 VPWR 0.28211f
C31582 _0181_ _1063_/a_193_47# 0
C31583 VPWR _0221_ 2.05385f
C31584 clkbuf_0_clk/a_110_47# _0486_ 0.00542f
C31585 _0955_/a_304_297# comp0.B\[5\] 0.01462f
C31586 _0955_/a_32_297# _0474_ 0.3732f
C31587 pp[9] _0510_/a_27_297# 0
C31588 net57 hold95/a_49_47# 0
C31589 _0567_/a_109_47# _0345_ 0
C31590 hold44/a_285_47# acc0.A\[29\] 0.06676f
C31591 _0311_ _0748_/a_299_297# 0.02901f
C31592 _0680_/a_300_47# _0294_ 0
C31593 _0150_ acc0.A\[6\] 0.23459f
C31594 _0524_/a_109_47# _0987_/a_27_47# 0
C31595 net165 _0261_ 0
C31596 clknet_1_1__leaf__0459_ _0799_/a_303_47# 0
C31597 _0216_ _0116_ 0.00525f
C31598 _0252_ _0828_/a_113_297# 0
C31599 hold33/a_391_47# comp0.B\[8\] 0.00596f
C31600 hold33/a_285_47# _0206_ 0
C31601 net55 _1010_/a_891_413# 0
C31602 VPWR _0813_/a_109_297# 0.00442f
C31603 _0163_ clknet_1_0__leaf__0457_ 0
C31604 _0181_ _0460_ 0.05419f
C31605 hold21/a_285_47# _0152_ 0.00185f
C31606 hold75/a_391_47# _0399_ 0.0213f
C31607 _0165_ _1067_/a_381_47# 0.12891f
C31608 _0616_/a_78_199# _0350_ 0
C31609 clkload2/a_110_47# _0180_ 0
C31610 _1042_/a_27_47# _1042_/a_193_47# 0.96191f
C31611 _0181_ _1060_/a_193_47# 0.46782f
C31612 _0183_ _0218_ 0.05739f
C31613 control0.add _0772_/a_215_47# 0
C31614 _0172_ _0545_/a_68_297# 0.01482f
C31615 hold45/a_391_47# clknet_1_1__leaf__0465_ 0.00135f
C31616 _0516_/a_27_297# _0516_/a_373_47# 0.01338f
C31617 clknet_0__0457_ _1019_/a_592_47# 0.00175f
C31618 _0423_ _0656_/a_59_75# 0
C31619 _1010_/a_193_47# _0352_ 0.03358f
C31620 net158 clkbuf_1_0__f__0464_/a_110_47# 0
C31621 _0238_ net92 0.15576f
C31622 clknet_1_1__leaf__0460_ _0730_/a_297_297# 0
C31623 _1051_/a_1059_315# clknet_1_1__leaf__0464_ 0
C31624 _0531_/a_109_297# _1061_/a_1059_315# 0
C31625 net48 clknet_1_0__leaf__0460_ 0.0636f
C31626 hold63/a_49_47# _0216_ 0.00262f
C31627 hold63/a_285_47# net155 0.00109f
C31628 hold63/a_391_47# _0195_ 0
C31629 _1045_/a_381_47# clknet_1_1__leaf__0464_ 0
C31630 _0458_ _0844_/a_79_21# 0.00664f
C31631 _1036_/a_193_47# _1036_/a_592_47# 0.00135f
C31632 _1036_/a_466_413# _1036_/a_561_413# 0.00772f
C31633 _1036_/a_634_159# _1036_/a_975_413# 0
C31634 net179 _0153_ 0.00217f
C31635 _0457_ _0181_ 0.08162f
C31636 control0.sh _0563_/a_51_297# 0
C31637 _0314_ acc0.A\[25\] 0.01747f
C31638 _0386_ _0388_ 0.67995f
C31639 hold26/a_49_47# _0172_ 0.00242f
C31640 hold26/a_391_47# net180 0.00132f
C31641 _0517_/a_81_21# _0988_/a_1059_315# 0
C31642 _1012_/a_891_413# _0778_/a_68_297# 0
C31643 net53 clkbuf_1_0__f__0462_/a_110_47# 0.04262f
C31644 _0578_/a_27_297# net187 0.05719f
C31645 _0372_ _0772_/a_79_21# 0
C31646 net8 _0176_ 0.66082f
C31647 _1049_/a_891_413# net11 0
C31648 _0582_/a_27_297# _0242_ 0
C31649 _0347_ _1009_/a_891_413# 0
C31650 _0222_ _0237_ 0.00527f
C31651 _0725_/a_80_21# _0353_ 0.28819f
C31652 _0176_ net32 0
C31653 _1041_/a_891_413# _0204_ 0
C31654 pp[9] _0181_ 0.00476f
C31655 _0732_/a_209_297# _1007_/a_27_47# 0
C31656 _0732_/a_80_21# _1007_/a_193_47# 0
C31657 _1050_/a_1059_315# net12 0
C31658 acc0.A\[21\] net150 0.30855f
C31659 _0144_ _0138_ 0.00156f
C31660 comp0.B\[2\] _0214_ 0.01783f
C31661 _1044_/a_592_47# net130 0
C31662 pp[28] hold62/a_285_47# 0.00185f
C31663 _0369_ clkbuf_1_1__f__0458_/a_110_47# 0.03329f
C31664 clknet_1_0__leaf__0462_ _1026_/a_27_47# 0.00903f
C31665 _0483_ _0981_/a_109_297# 0.0549f
C31666 hold49/a_49_47# net195 0
C31667 _0996_/a_891_413# _0219_ 0
C31668 hold33/a_285_47# _1046_/a_1059_315# 0
C31669 hold33/a_49_47# _1046_/a_891_413# 0
C31670 _0163_ _1062_/a_466_413# 0
C31671 _0576_/a_109_297# VPWR 0.1879f
C31672 clknet_1_0__leaf__0462_ _1024_/a_1059_315# 0.00472f
C31673 _0467_ _1063_/a_1059_315# 0.00333f
C31674 _1058_/a_466_413# net4 0.03396f
C31675 _1058_/a_193_47# _0187_ 0
C31676 _0848_/a_27_47# acc0.A\[15\] 0.0024f
C31677 _0416_ net39 0
C31678 _0415_ acc0.A\[12\] 0.00757f
C31679 hold32/a_49_47# net47 0
C31680 _1021_/a_466_413# _0181_ 0.00415f
C31681 _0467_ _0959_/a_80_21# 0.21248f
C31682 _1052_/a_1059_315# _0518_/a_109_297# 0
C31683 hold19/a_285_47# _0583_/a_27_297# 0.00104f
C31684 output36/a_27_47# net172 0
C31685 _0476_ hold39/a_49_47# 0.00317f
C31686 _0218_ acc0.A\[15\] 0.03341f
C31687 _0353_ _0128_ 0
C31688 _1012_/a_634_159# net239 0
C31689 _0428_ _0990_/a_381_47# 0
C31690 _0819_/a_81_21# _0088_ 0
C31691 net233 _0447_ 0.00184f
C31692 net234 _0346_ 0
C31693 _0195_ _0721_/a_27_47# 0
C31694 _0467_ net159 0.0294f
C31695 net23 net118 0.03877f
C31696 _0736_/a_139_47# _0107_ 0.00181f
C31697 _0458_ _0846_/a_240_47# 0
C31698 _1057_/a_466_413# net189 0.03268f
C31699 _0803_/a_68_297# _0404_ 0.06202f
C31700 _0174_ clknet_0__0463_ 0.08244f
C31701 hold10/a_49_47# control0.sh 0
C31702 _0379_ net51 0.00579f
C31703 B[13] _1042_/a_1017_47# 0
C31704 _0250_ _1007_/a_193_47# 0
C31705 _1053_/a_27_47# _1052_/a_27_47# 0.00125f
C31706 _0179_ hold28/a_391_47# 0.04776f
C31707 _0216_ hold62/a_391_47# 0
C31708 _0093_ _0995_/a_634_159# 0
C31709 net46 _0346_ 0.0197f
C31710 _0789_/a_201_297# _0299_ 0.01103f
C31711 _0789_/a_208_47# _0404_ 0.00175f
C31712 _0789_/a_544_297# _0298_ 0.00733f
C31713 _1059_/a_1059_315# net145 0
C31714 _0732_/a_80_21# _0328_ 0.12336f
C31715 _0754_/a_51_297# _0754_/a_512_297# 0.0116f
C31716 control0.sh _0549_/a_68_297# 0.02283f
C31717 _0344_ VPWR 0.55185f
C31718 net165 net47 0.0288f
C31719 net208 _0345_ 0.02499f
C31720 _0959_/a_80_21# comp0.B\[0\] 0
C31721 _0470_ _0951_/a_209_311# 0.08893f
C31722 _0313_ _0737_/a_35_297# 0.03039f
C31723 _0252_ _0433_ 0
C31724 _1055_/a_634_159# clknet_1_1__leaf__0465_ 0.00312f
C31725 _0811_/a_384_47# _0283_ 0
C31726 _0855_/a_81_21# _0465_ 0.00106f
C31727 net120 _0213_ 0
C31728 _0779_/a_215_47# _0347_ 0.05719f
C31729 _0176_ _1042_/a_1059_315# 0.00683f
C31730 _0312_ _0462_ 0.07779f
C31731 _0767_/a_59_75# _0369_ 0.00401f
C31732 clknet_1_0__leaf_clk _1068_/a_1059_315# 0
C31733 _0673_/a_103_199# _0295_ 0.10278f
C31734 _0432_ _0986_/a_193_47# 0
C31735 _0352_ _0771_/a_298_297# 0
C31736 net168 hold83/a_391_47# 0.08002f
C31737 _1002_/a_1059_315# _0578_/a_109_297# 0
C31738 _1002_/a_891_413# _0578_/a_27_297# 0
C31739 comp0.B\[13\] _0142_ 0
C31740 _0407_ _0791_/a_113_297# 0.09866f
C31741 output43/a_27_47# net245 0
C31742 pp[16] hold98/a_391_47# 0
C31743 _0992_/a_193_47# _0281_ 0
C31744 _0154_ net16 0
C31745 _1046_/a_1059_315# net20 0
C31746 _0536_/a_512_297# net22 0
C31747 net47 acc0.A\[19\] 0
C31748 control0.state\[1\] hold85/a_49_47# 0.00399f
C31749 control0.state\[0\] hold85/a_285_47# 0.00914f
C31750 _0974_/a_222_93# _1068_/a_193_47# 0.00543f
C31751 _0328_ _0250_ 0.0036f
C31752 _0852_/a_35_297# _0268_ 0
C31753 _0176_ net10 0.10489f
C31754 VPWR _1008_/a_975_413# 0.00507f
C31755 _0456_ hold60/a_49_47# 0
C31756 hold43/a_49_47# VPWR 0.28833f
C31757 _0476_ hold58/a_391_47# 0.0056f
C31758 _0180_ _0148_ 0.03124f
C31759 hold11/a_391_47# net132 0
C31760 _0338_ _0723_/a_297_47# 0
C31761 _0343_ _0988_/a_193_47# 0
C31762 _1028_/a_193_47# _1027_/a_891_413# 0
C31763 _1020_/a_1059_315# net87 0
C31764 hold75/a_49_47# _0345_ 0
C31765 _0691_/a_68_297# clknet_0__0462_ 0
C31766 _0179_ _0218_ 0.02142f
C31767 acc0.A\[21\] control0.add 0
C31768 net86 _0582_/a_27_297# 0
C31769 net117 _0342_ 0
C31770 _0222_ _1005_/a_27_47# 0
C31771 clknet_0__0464_ _0197_ 0
C31772 net5 _0668_/a_297_47# 0
C31773 _0439_ _0434_ 0
C31774 _0341_ _1013_/a_466_413# 0
C31775 _0785_/a_81_21# _0427_ 0.04464f
C31776 _0305_ _1017_/a_1059_315# 0.03442f
C31777 net186 _0131_ 0.00148f
C31778 hold10/a_49_47# net157 0.04725f
C31779 VPWR _0434_ 0.62567f
C31780 clknet_1_0__leaf__0463_ _0536_/a_512_297# 0
C31781 clknet_0__0463_ _0208_ 0.68027f
C31782 _0218_ hold40/a_285_47# 0
C31783 net231 net17 0.02663f
C31784 _0183_ _0112_ 0
C31785 _0299_ _0995_/a_466_413# 0.00137f
C31786 _0589_/a_113_47# acc0.A\[29\] 0
C31787 _0695_/a_80_21# _0695_/a_217_297# 0.12661f
C31788 net104 _0634_/a_113_47# 0
C31789 _0227_ _0378_ 0.05679f
C31790 _0361_ hold90/a_285_47# 0
C31791 _0467_ _0173_ 0
C31792 net108 _0577_/a_109_297# 0
C31793 clknet_1_0__leaf__0462_ _0577_/a_373_47# 0.00183f
C31794 comp0.B\[10\] _0544_/a_51_297# 0.1157f
C31795 _1031_/a_27_47# _1031_/a_466_413# 0.27314f
C31796 _1031_/a_193_47# _1031_/a_634_159# 0.11949f
C31797 _0292_ _0818_/a_109_47# 0
C31798 clknet_1_0__leaf__0463_ _0547_/a_150_297# 0
C31799 _0982_/a_27_47# clknet_1_1__leaf__0457_ 0
C31800 _0517_/a_299_297# _0186_ 0
C31801 _0343_ net72 0
C31802 net45 _0778_/a_150_297# 0
C31803 input31/a_75_212# net152 0
C31804 _0996_/a_27_47# _0346_ 0
C31805 output43/a_27_47# net45 0.0019f
C31806 _0476_ hold57/a_285_47# 0
C31807 _0121_ hold96/a_391_47# 0
C31808 hold30/a_49_47# net243 0
C31809 control0.state\[1\] _1063_/a_975_413# 0.00184f
C31810 _1000_/a_27_47# _0294_ 0.00532f
C31811 hold53/a_49_47# acc0.A\[24\] 0
C31812 _1005_/a_634_159# _1005_/a_592_47# 0
C31813 _0813_/a_109_297# _0283_ 0
C31814 net178 hold88/a_285_47# 0
C31815 _0244_ _0616_/a_78_199# 0.00286f
C31816 _0145_ clknet_1_1__leaf__0457_ 0.02154f
C31817 _0984_/a_466_413# _0082_ 0.04689f
C31818 _0984_/a_381_47# net222 0
C31819 _0646_/a_47_47# _0646_/a_129_47# 0.00369f
C31820 _1060_/a_1059_315# _0507_/a_27_297# 0.01884f
C31821 _1013_/a_634_159# _1013_/a_381_47# 0
C31822 net149 _0117_ 0
C31823 _0125_ _0106_ 0
C31824 _1002_/a_193_47# _1002_/a_466_413# 0.07482f
C31825 _1002_/a_27_47# _1002_/a_1059_315# 0.04861f
C31826 _0144_ net134 0.01105f
C31827 comp0.B\[0\] _0173_ 0.02601f
C31828 hold64/a_391_47# clkbuf_0__0457_/a_110_47# 0.01439f
C31829 _1027_/a_193_47# _0739_/a_79_21# 0
C31830 hold26/a_285_47# hold26/a_391_47# 0.41909f
C31831 hold46/a_391_47# net22 0
C31832 _0689_/a_68_297# _0687_/a_59_75# 0.00686f
C31833 output65/a_27_47# pp[7] 0.33841f
C31834 _0415_ _0993_/a_592_47# 0
C31835 _0984_/a_27_47# clknet_1_0__leaf__0458_ 0.00471f
C31836 _1027_/a_634_159# _0347_ 0
C31837 _0177_ acc0.A\[15\] 0.04939f
C31838 _0773_/a_35_297# _0771_/a_27_413# 0
C31839 _0749_/a_299_297# _0373_ 0.00103f
C31840 net243 _0352_ 0.00134f
C31841 _0985_/a_592_47# _0261_ 0
C31842 _0607_/a_109_47# acc0.A\[16\] 0
C31843 _0286_ _0091_ 0
C31844 net165 _1060_/a_1059_315# 0
C31845 clknet_0_clk hold84/a_285_47# 0
C31846 VPWR acc0.A\[7\] 1.49405f
C31847 hold35/a_49_47# _1055_/a_193_47# 0
C31848 hold35/a_285_47# _1055_/a_27_47# 0
C31849 VPWR _0989_/a_1059_315# 0.37227f
C31850 _0183_ net240 0
C31851 VPWR _0997_/a_27_47# 0.50302f
C31852 net178 _0086_ 0.21338f
C31853 net68 acc0.A\[0\] 0.00345f
C31854 _0795_/a_81_21# _0405_ 0.06918f
C31855 _0180_ _0525_/a_384_47# 0.00128f
C31856 _1038_/a_891_413# _1040_/a_466_413# 0
C31857 _0217_ _1019_/a_193_47# 0.02083f
C31858 VPWR _0992_/a_1059_315# 0.40231f
C31859 _0600_/a_253_47# _0232_ 0.00764f
C31860 _0112_ acc0.A\[15\] 0
C31861 _0183_ _0099_ 0.00451f
C31862 _0734_/a_377_297# _0361_ 0.00284f
C31863 _1018_/a_1059_315# net221 0
C31864 control0.state\[0\] _0958_/a_27_47# 0.01426f
C31865 VPWR hold94/a_285_47# 0.27998f
C31866 comp0.B\[9\] _0142_ 0
C31867 output66/a_27_47# acc0.A\[11\] 0.00857f
C31868 _0995_/a_1059_315# _0995_/a_1017_47# 0
C31869 _0765_/a_79_21# _0765_/a_510_47# 0.00844f
C31870 _0765_/a_297_297# _0765_/a_215_47# 0
C31871 hold65/a_285_47# _0186_ 0.00211f
C31872 _0346_ _0654_/a_207_413# 0.02799f
C31873 hold46/a_391_47# clknet_1_0__leaf__0463_ 0
C31874 output56/a_27_47# _1011_/a_193_47# 0
C31875 VPWR _1061_/a_634_159# 0.19148f
C31876 hold23/a_49_47# _0447_ 0
C31877 _1015_/a_27_47# control0.reset 0
C31878 pp[28] _0350_ 0
C31879 _0983_/a_561_413# _0346_ 0
C31880 _0783_/a_297_297# _0306_ 0
C31881 _0534_/a_81_21# _1048_/a_891_413# 0
C31882 _0534_/a_299_297# _1048_/a_1059_315# 0
C31883 _1017_/a_891_413# _0675_/a_68_297# 0
C31884 _1034_/a_634_159# _0173_ 0.00236f
C31885 _1034_/a_466_413# _0213_ 0.01282f
C31886 _0679_/a_68_297# _0350_ 0
C31887 _0629_/a_145_75# VPWR 0
C31888 _0529_/a_27_297# _0449_ 0
C31889 control0.state\[1\] _0973_/a_27_297# 0.00167f
C31890 clknet_1_0__leaf__0458_ net10 0
C31891 hold87/a_49_47# _0454_ 0
C31892 _0183_ _0581_/a_109_47# 0.00137f
C31893 _1035_/a_27_47# control0.sh 0.00197f
C31894 _0605_/a_109_297# _0228_ 0.00112f
C31895 _1000_/a_27_47# _0775_/a_297_297# 0
C31896 _0139_ _1042_/a_891_413# 0
C31897 net32 _1042_/a_975_413# 0.00251f
C31898 hold54/a_49_47# _0216_ 0.00255f
C31899 _0251_ _0622_/a_193_47# 0
C31900 _0369_ _0291_ 0
C31901 hold86/a_391_47# acc0.A\[15\] 0.00503f
C31902 _1019_/a_891_413# _0580_/a_27_297# 0
C31903 _1019_/a_1059_315# _0580_/a_109_297# 0
C31904 acc0.A\[29\] _0219_ 0.09133f
C31905 _1070_/a_27_47# control0.count\[0\] 0.0023f
C31906 _1070_/a_1059_315# clknet_1_0__leaf_clk 0
C31907 control0.count\[1\] _1069_/a_27_47# 0.02178f
C31908 VPWR _1069_/a_891_413# 0.17722f
C31909 _0226_ _0749_/a_81_21# 0.02353f
C31910 _0269_ _0846_/a_51_297# 0.01708f
C31911 _0268_ _0846_/a_149_47# 0
C31912 output53/a_27_47# hold53/a_49_47# 0.02053f
C31913 hold27/a_49_47# _0138_ 0.31773f
C31914 _1034_/a_891_413# _0475_ 0
C31915 comp0.B\[12\] _1045_/a_1059_315# 0.00136f
C31916 net15 output63/a_27_47# 0
C31917 _0695_/a_80_21# _0743_/a_149_47# 0
C31918 _1052_/a_891_413# _0987_/a_27_47# 0
C31919 acc0.A\[30\] net209 0.00406f
C31920 _1011_/a_1059_315# net97 0
C31921 VPWR B[1] 0.1383f
C31922 _1011_/a_27_47# net57 0.00423f
C31923 A[10] acc0.A\[10\] 0.01219f
C31924 _0985_/a_1059_315# _0186_ 0
C31925 net166 _0369_ 0.00408f
C31926 _0316_ clkbuf_1_1__f__0460_/a_110_47# 0.07293f
C31927 _0728_/a_59_75# acc0.A\[29\] 0.0119f
C31928 net81 _0400_ 0
C31929 _1055_/a_193_47# A[9] 0
C31930 _0195_ clkbuf_1_0__f__0461_/a_110_47# 0
C31931 _0216_ _0380_ 0
C31932 _1006_/a_27_47# _1006_/a_561_413# 0.0027f
C31933 _1006_/a_634_159# _1006_/a_891_413# 0.03684f
C31934 _1006_/a_193_47# _1006_/a_381_47# 0.09503f
C31935 _0538_/a_240_47# VPWR 0.00137f
C31936 _0993_/a_634_159# _0807_/a_68_297# 0
C31937 _1049_/a_193_47# _0186_ 0
C31938 clknet_1_1__leaf__0461_ _1060_/a_193_47# 0
C31939 _0532_/a_384_47# net218 0.01033f
C31940 acc0.A\[1\] _1014_/a_193_47# 0
C31941 _0182_ _1014_/a_27_47# 0
C31942 acc0.A\[17\] _0459_ 0.01846f
C31943 net206 _0580_/a_27_297# 0.06252f
C31944 _0482_ _0480_ 0.31622f
C31945 _0984_/a_193_47# _0984_/a_466_413# 0.07482f
C31946 _0984_/a_27_47# _0984_/a_1059_315# 0.04819f
C31947 clkbuf_1_1__f__0460_/a_110_47# _0347_ 0.02747f
C31948 acc0.A\[12\] _0347_ 0.06488f
C31949 net185 _1034_/a_1059_315# 0.00183f
C31950 _0572_/a_27_297# acc0.A\[25\] 0
C31951 _0124_ _1025_/a_381_47# 0
C31952 _0808_/a_368_297# _0808_/a_266_47# 0.00153f
C31953 _1055_/a_1017_47# VPWR 0.00144f
C31954 _0399_ hold2/a_285_47# 0
C31955 _1018_/a_561_413# clknet_1_0__leaf__0461_ 0
C31956 hold66/a_285_47# hold3/a_285_47# 0.02819f
C31957 _0102_ _1024_/a_891_413# 0
C31958 _0217_ net49 0.06149f
C31959 _1003_/a_592_47# VPWR 0
C31960 _0429_ _0435_ 0.50971f
C31961 hold65/a_391_47# _0253_ 0
C31962 clkbuf_0__0464_/a_110_47# net135 0.00364f
C31963 _0441_ _0218_ 0.04494f
C31964 _1039_/a_634_159# VPWR 0.17546f
C31965 pp[9] _0187_ 0
C31966 control0.state\[0\] hold79/a_391_47# 0
C31967 _0986_/a_27_47# _0986_/a_561_413# 0.0027f
C31968 _0986_/a_634_159# _0986_/a_891_413# 0.03684f
C31969 _0986_/a_193_47# _0986_/a_381_47# 0.09503f
C31970 _0520_/a_27_297# _1054_/a_27_47# 0
C31971 _0524_/a_27_297# net73 0.01034f
C31972 net148 _0987_/a_561_413# 0
C31973 _0361_ clknet_0__0462_ 0.20034f
C31974 clkbuf_1_0__f__0458_/a_110_47# _0268_ 0.01205f
C31975 hold43/a_391_47# _0569_/a_27_297# 0.00134f
C31976 _1023_/a_634_159# _1023_/a_975_413# 0
C31977 _1023_/a_466_413# _1023_/a_561_413# 0.00772f
C31978 _1023_/a_193_47# _1023_/a_592_47# 0
C31979 _1017_/a_1059_315# _0181_ 0.02225f
C31980 net120 _0161_ 0
C31981 _0747_/a_215_47# acc0.A\[24\] 0
C31982 _0300_ _0669_/a_29_53# 0.0919f
C31983 net22 net153 0.05355f
C31984 _1042_/a_466_413# _1042_/a_592_47# 0.00553f
C31985 _1042_/a_634_159# _1042_/a_1017_47# 0
C31986 _1019_/a_634_159# control0.add 0
C31987 _0718_/a_47_47# _0723_/a_207_413# 0
C31988 _0195_ acc0.A\[5\] 0
C31989 net232 _0467_ 0
C31990 control0.state\[1\] net17 0.27442f
C31991 _0516_/a_373_47# _0190_ 0
C31992 clknet_1_1__leaf__0464_ _1044_/a_891_413# 0.03162f
C31993 _1011_/a_891_413# _0707_/a_75_199# 0
C31994 _1011_/a_1059_315# _0707_/a_201_297# 0
C31995 _1045_/a_634_159# net20 0
C31996 _0459_ net5 0.0084f
C31997 hold68/a_285_47# acc0.A\[23\] 0.01765f
C31998 hold86/a_391_47# _0179_ 0
C31999 _0179_ _1050_/a_592_47# 0
C32000 _0413_ _0219_ 0.18602f
C32001 _0347_ _0445_ 0
C32002 net125 _0493_/a_27_47# 0
C32003 _1036_/a_1059_315# comp0.B\[4\] 0.11723f
C32004 _1036_/a_561_413# net161 0
C32005 _0466_ _1064_/a_1059_315# 0.00126f
C32006 _0195_ _0528_/a_299_297# 0.05488f
C32007 _0254_ _0990_/a_27_47# 0
C32008 hold16/a_49_47# _1031_/a_193_47# 0
C32009 hold16/a_285_47# _1031_/a_27_47# 0.00329f
C32010 _0305_ _0508_/a_384_47# 0
C32011 net43 _0094_ 0
C32012 hold18/a_391_47# _0182_ 0
C32013 _0153_ _0988_/a_561_413# 0
C32014 _0984_/a_466_413# net145 0
C32015 VPWR _0421_ 0.303f
C32016 clknet_1_0__leaf__0463_ net153 0.14661f
C32017 net9 hold7/a_49_47# 0.00557f
C32018 _1059_/a_193_47# _0506_/a_299_297# 0
C32019 _1059_/a_27_47# _0506_/a_384_47# 0
C32020 _0808_/a_368_297# _0345_ 0
C32021 net165 _0848_/a_109_297# 0.0012f
C32022 _0621_/a_285_297# _0369_ 0
C32023 _1057_/a_1059_315# _0511_/a_299_297# 0
C32024 _0746_/a_299_297# _0462_ 0.01034f
C32025 pp[29] _1011_/a_466_413# 0
C32026 _1038_/a_27_47# _1037_/a_27_47# 0
C32027 VPWR _1040_/a_1017_47# 0
C32028 _0992_/a_561_413# clknet_1_1__leaf__0465_ 0
C32029 hold52/a_285_47# net215 0
C32030 _0294_ net165 0.44389f
C32031 _0997_/a_193_47# _0407_ 0
C32032 _0183_ net228 0
C32033 _0290_ _0369_ 0.27576f
C32034 _0366_ _0352_ 0
C32035 control0.reset _0215_ 0.02599f
C32036 _0426_ net47 0
C32037 _0743_/a_245_297# _0743_/a_240_47# 0
C32038 hold88/a_391_47# pp[1] 0
C32039 _0777_/a_377_297# _0308_ 0
C32040 _1002_/a_634_159# net220 0
C32041 _1054_/a_466_413# net11 0.00265f
C32042 _1019_/a_27_47# hold40/a_49_47# 0
C32043 hold85/a_391_47# _1066_/a_27_47# 0
C32044 control0.state\[0\] _0481_ 0.00123f
C32045 _0163_ _0160_ 0
C32046 _0251_ _1054_/a_891_413# 0
C32047 _0099_ hold40/a_285_47# 0
C32048 net192 _0286_ 0.0017f
C32049 _0195_ _0182_ 0.13308f
C32050 _0662_/a_81_21# _0293_ 0.1863f
C32051 _0119_ _0181_ 0.03173f
C32052 hold19/a_285_47# _0114_ 0.06875f
C32053 acc0.A\[25\] _0360_ 0.001f
C32054 clknet_0__0463_ comp0.B\[9\] 0.01156f
C32055 net215 net52 0.00763f
C32056 hold30/a_49_47# net151 0
C32057 _0999_/a_381_47# _0218_ 0.02059f
C32058 _0179_ net15 0.13305f
C32059 _0195_ _1013_/a_27_47# 0.03228f
C32060 _0346_ _0286_ 0.37653f
C32061 net33 comp0.B\[5\] 0
C32062 _0311_ _0246_ 0.09247f
C32063 clknet_1_0__leaf__0464_ _1049_/a_561_413# 0
C32064 net188 input2/a_75_212# 0
C32065 _0548_/a_51_297# net152 0
C32066 _1058_/a_381_47# acc0.A\[11\] 0
C32067 clkbuf_0__0463_/a_110_47# _0159_ 0
C32068 _0463_ net7 0
C32069 _0984_/a_561_413# net77 0
C32070 net70 _0991_/a_561_413# 0
C32071 _0363_ _0219_ 0.15762f
C32072 _0183_ hold3/a_285_47# 0
C32073 VPWR _1035_/a_891_413# 0.19679f
C32074 A[10] _0510_/a_109_297# 0
C32075 net180 _1040_/a_27_47# 0.00306f
C32076 _0754_/a_512_297# _0219_ 0
C32077 _0754_/a_149_47# net241 0.00147f
C32078 _0754_/a_240_47# _0377_ 0.04154f
C32079 _0272_ _0271_ 0.0012f
C32080 _0274_ _0256_ 0
C32081 _0275_ _0270_ 0
C32082 _0982_/a_1059_315# _0181_ 0.08209f
C32083 _0343_ _0336_ 0.21854f
C32084 VPWR _0809_/a_81_21# 0.20881f
C32085 _0179_ _1053_/a_1059_315# 0
C32086 _0992_/a_1059_315# _0283_ 0.00119f
C32087 hold27/a_49_47# net134 0
C32088 _0404_ _0669_/a_29_53# 0.00116f
C32089 _0304_ _0345_ 0.01088f
C32090 _1055_/a_193_47# _0516_/a_27_297# 0
C32091 _1064_/a_634_159# _1064_/a_466_413# 0.23992f
C32092 _1064_/a_193_47# _1064_/a_1059_315# 0.03389f
C32093 _1064_/a_27_47# _1064_/a_891_413# 0.03089f
C32094 net141 clknet_1_1__leaf__0465_ 0.18121f
C32095 _0643_/a_253_297# _0431_ 0
C32096 _1018_/a_193_47# net149 0
C32097 _0097_ _0352_ 0.07532f
C32098 clknet_1_1__leaf__0459_ _0786_/a_300_47# 0
C32099 net228 acc0.A\[15\] 0.01041f
C32100 clknet_0__0457_ acc0.A\[1\] 0.01599f
C32101 _1054_/a_466_413# hold7/a_391_47# 0
C32102 clk _1068_/a_891_413# 0
C32103 _1018_/a_1059_315# _1017_/a_27_47# 0
C32104 _1000_/a_27_47# _0581_/a_109_297# 0
C32105 net204 _0210_ 0.0022f
C32106 _0243_ _0634_/a_113_47# 0
C32107 _1047_/a_27_47# _0171_ 0
C32108 _0255_ _0826_/a_301_297# 0.00141f
C32109 _0346_ _0794_/a_27_47# 0
C32110 net226 control0.state\[2\] 0
C32111 _0435_ clknet_1_1__leaf__0458_ 0
C32112 VPWR _0778_/a_150_297# 0.00144f
C32113 clknet_1_1__leaf__0460_ _0105_ 0.00222f
C32114 _0712_/a_79_21# _0712_/a_465_47# 0
C32115 _0712_/a_297_297# _0712_/a_381_47# 0
C32116 _0574_/a_109_297# _0366_ 0
C32117 output43/a_27_47# VPWR 0.29573f
C32118 _1051_/a_1059_315# net148 0.00151f
C32119 _1051_/a_193_47# net12 0
C32120 net31 clkbuf_1_0__f__0463_/a_110_47# 0.0015f
C32121 _0144_ net22 0
C32122 VPWR _0994_/a_1017_47# 0
C32123 _0343_ _1060_/a_561_413# 0
C32124 _0520_/a_109_297# VPWR 0.19075f
C32125 net1 net159 0
C32126 _0968_/a_109_297# _0487_ 0
C32127 VPWR _0696_/a_109_297# 0.00495f
C32128 pp[31] pp[14] 0.00582f
C32129 _0373_ hold73/a_49_47# 0
C32130 _0695_/a_80_21# net52 0
C32131 clknet_0__0465_ _0841_/a_510_47# 0
C32132 clkbuf_0__0465_/a_110_47# _0445_ 0.00102f
C32133 _0946_/a_112_297# control0.state\[2\] 0
C32134 _1017_/a_891_413# _0677_/a_47_47# 0
C32135 net114 _1027_/a_1059_315# 0.00178f
C32136 net154 _0522_/a_27_297# 0
C32137 net106 _1067_/a_891_413# 0
C32138 _0553_/a_149_47# _0209_ 0.00154f
C32139 _1010_/a_975_413# _0350_ 0.00168f
C32140 output55/a_27_47# net97 0
C32141 _0399_ _0437_ 0.06527f
C32142 _0181_ _0451_ 0
C32143 _0737_/a_117_297# _0360_ 0.00777f
C32144 _0737_/a_35_297# _0321_ 0.08557f
C32145 _0317_ _0690_/a_68_297# 0.01689f
C32146 _0854_/a_79_21# _0854_/a_297_297# 0.01735f
C32147 _0259_ _0990_/a_891_413# 0
C32148 net86 _0115_ 0
C32149 clknet_1_1__leaf__0464_ _1042_/a_27_47# 0
C32150 _0216_ _0386_ 0
C32151 _0697_/a_80_21# _0329_ 0.11839f
C32152 _0697_/a_217_297# _0322_ 0.00382f
C32153 _0176_ _0492_/a_27_47# 0
C32154 net60 _0220_ 0.00133f
C32155 input21/a_75_212# comp0.B\[11\] 0.00202f
C32156 _0347_ net42 0.0015f
C32157 net157 _1061_/a_975_413# 0
C32158 net56 _0329_ 0.02796f
C32159 _0989_/a_634_159# acc0.A\[6\] 0
C32160 _0305_ _1016_/a_27_47# 0
C32161 _0420_ hold81/a_391_47# 0.00342f
C32162 clknet_1_0__leaf__0463_ _0144_ 0.00234f
C32163 _0712_/a_79_21# hold16/a_285_47# 0
C32164 _0830_/a_79_21# _0830_/a_215_47# 0.04584f
C32165 clknet_0__0458_ _0991_/a_27_47# 0
C32166 _0174_ net198 0.11241f
C32167 _0695_/a_472_297# _0327_ 0
C32168 clkbuf_1_1__f__0465_/a_110_47# _0992_/a_27_47# 0.00122f
C32169 clknet_1_0__leaf__0465_ _1052_/a_27_47# 0.00985f
C32170 _1034_/a_381_47# _1033_/a_27_47# 0
C32171 _1034_/a_27_47# _1033_/a_381_47# 0
C32172 _1037_/a_634_159# VPWR 0.19044f
C32173 _0837_/a_266_297# acc0.A\[4\] 0
C32174 _0217_ _1016_/a_381_47# 0
C32175 net175 _1047_/a_193_47# 0
C32176 _1031_/a_1059_315# _1031_/a_1017_47# 0
C32177 _0289_ _0786_/a_472_297# 0
C32178 net67 net37 0.63632f
C32179 hold30/a_49_47# _0378_ 0.00822f
C32180 A[10] _0188_ 0.00267f
C32181 _0733_/a_79_199# _0324_ 0.05551f
C32182 _1041_/a_891_413# VPWR 0.18277f
C32183 _0092_ _0403_ 0.10693f
C32184 pp[15] _0995_/a_1059_315# 0.00222f
C32185 _0179_ net228 0.28755f
C32186 _1005_/a_975_413# _0103_ 0
C32187 net17 _0565_/a_245_297# 0.00143f
C32188 _0260_ _0529_/a_27_297# 0
C32189 _0438_ _0831_/a_35_297# 0.16735f
C32190 _0388_ _0240_ 0.504f
C32191 net56 _0221_ 0.05215f
C32192 _0326_ _0315_ 0
C32193 _1066_/a_27_47# _0160_ 0.00122f
C32194 clknet_1_1__leaf_clk _1062_/a_193_47# 0.14966f
C32195 _1056_/a_193_47# pp[9] 0
C32196 acc0.A\[29\] hold61/a_49_47# 0
C32197 _0902_/a_27_47# _0346_ 0
C32198 _0082_ _0506_/a_81_21# 0
C32199 _1060_/a_381_47# net5 0
C32200 _1060_/a_1059_315# _0185_ 0.03836f
C32201 _1020_/a_27_47# _1020_/a_634_159# 0.14145f
C32202 _1002_/a_193_47# _0100_ 0.57422f
C32203 _1002_/a_891_413# _1002_/a_1017_47# 0.00617f
C32204 _1002_/a_634_159# net88 0.00468f
C32205 acc0.A\[23\] _0754_/a_51_297# 0
C32206 _0405_ _0790_/a_117_297# 0
C32207 _0792_/a_209_297# net42 0
C32208 clknet_0__0458_ _0350_ 0.19264f
C32209 net103 _0583_/a_27_297# 0
C32210 _1017_/a_634_159# _0114_ 0
C32211 _1027_/a_1059_315# _0365_ 0
C32212 _1027_/a_634_159# _0106_ 0
C32213 _0352_ _0378_ 0
C32214 _0347_ _0379_ 0.10482f
C32215 _1059_/a_1059_315# _0302_ 0
C32216 net63 _0440_ 0.45487f
C32217 net45 hold19/a_49_47# 0
C32218 control0.count\[3\] clknet_1_0__leaf_clk 0.12815f
C32219 _0983_/a_27_47# net47 0.42515f
C32220 _0343_ _0642_/a_298_297# 0.00235f
C32221 hold64/a_391_47# _0350_ 0.00321f
C32222 net53 _0324_ 0.04028f
C32223 _0217_ _0757_/a_68_297# 0
C32224 _1058_/a_193_47# clknet_1_1__leaf__0465_ 0.05172f
C32225 acc0.A\[3\] _0261_ 0
C32226 _0421_ _0283_ 0.2662f
C32227 _0957_/a_32_297# _0175_ 0
C32228 _0183_ _1019_/a_1017_47# 0
C32229 _0346_ _0673_/a_103_199# 0
C32230 _0180_ _1048_/a_27_47# 0.02534f
C32231 _0182_ _1048_/a_193_47# 0.00109f
C32232 _0998_/a_27_47# _1017_/a_27_47# 0
C32233 acc0.A\[12\] net2 0.03269f
C32234 net168 net9 0
C32235 _1001_/a_634_159# net46 0.00256f
C32236 pp[26] hold8/a_391_47# 0
C32237 _0346_ _0672_/a_79_21# 0.01736f
C32238 hold86/a_285_47# net165 0
C32239 control0.state\[0\] _0477_ 0.06605f
C32240 _1041_/a_193_47# _0550_/a_149_47# 0
C32241 _0285_ clknet_1_1__leaf__0459_ 0.21684f
C32242 _0284_ acc0.A\[11\] 0.05593f
C32243 hold88/a_49_47# _0181_ 0
C32244 _1003_/a_27_47# _0466_ 0.00302f
C32245 _0372_ _0104_ 0
C32246 VPWR net147 0.62109f
C32247 net23 _0175_ 0.00113f
C32248 _0151_ net138 0
C32249 net36 hold2/a_391_47# 0
C32250 _1021_/a_27_47# clkbuf_1_1__f_clk/a_110_47# 0
C32251 _0811_/a_384_47# _0345_ 0
C32252 _0231_ net93 0
C32253 pp[27] _0334_ 0.03579f
C32254 _0837_/a_81_21# _1051_/a_1059_315# 0
C32255 _0310_ clknet_0__0461_ 0
C32256 control0.count\[1\] _0489_ 0.14277f
C32257 control0.state\[1\] _0165_ 0.36705f
C32258 _1036_/a_27_47# B[1] 0
C32259 _0676_/a_113_47# _0347_ 0
C32260 _0172_ _0346_ 0.06677f
C32261 _0985_/a_891_413# _0446_ 0.01121f
C32262 _0413_ _0799_/a_209_297# 0.00323f
C32263 comp0.B\[12\] _1044_/a_466_413# 0
C32264 _0456_ _0263_ 0
C32265 net178 net66 0
C32266 _1066_/a_634_159# net17 0
C32267 _0534_/a_299_297# clkbuf_1_1__f__0457_/a_110_47# 0
C32268 clknet_1_1__leaf__0460_ _0690_/a_150_297# 0
C32269 VPWR input20/a_75_212# 0.22585f
C32270 _0967_/a_215_297# control0.state\[2\] 0.0662f
C32271 clknet_1_0__leaf__0458_ _1014_/a_891_413# 0
C32272 _0168_ _0167_ 0
C32273 _0486_ _0487_ 0.30016f
C32274 hold57/a_49_47# _0176_ 0
C32275 comp0.B\[2\] _0472_ 0.20362f
C32276 _0606_/a_215_297# _0374_ 0.01059f
C32277 _0414_ _0994_/a_466_413# 0
C32278 _0714_/a_51_297# net43 0
C32279 clknet_1_0__leaf__0462_ _0368_ 0.00112f
C32280 clkbuf_1_0__f__0458_/a_110_47# net222 0.00349f
C32281 _1017_/a_1059_315# clknet_1_1__leaf__0461_ 0.02722f
C32282 net69 _0465_ 0
C32283 _1000_/a_891_413# _0246_ 0
C32284 _0572_/a_27_297# net210 0.07732f
C32285 acc0.A\[14\] _0507_/a_109_297# 0.00168f
C32286 _0399_ _0301_ 0.00156f
C32287 _0216_ _1006_/a_466_413# 0.01659f
C32288 _1006_/a_891_413# net92 0
C32289 _0329_ _0345_ 0
C32290 VPWR _0974_/a_222_93# 0.08272f
C32291 acc0.A\[3\] _0509_/a_27_47# 0
C32292 net206 _0117_ 0
C32293 _0283_ _0809_/a_81_21# 0
C32294 acc0.A\[14\] hold82/a_49_47# 0
C32295 net133 _0171_ 0
C32296 clknet_1_0__leaf__0460_ _0345_ 0.00166f
C32297 hold10/a_391_47# _0137_ 0
C32298 pp[30] _0341_ 0
C32299 _0984_/a_891_413# _0984_/a_1017_47# 0.00617f
C32300 _0984_/a_634_159# net70 0
C32301 _0172_ _1061_/a_193_47# 0.0148f
C32302 _0643_/a_253_297# _0269_ 0.00613f
C32303 _0573_/a_27_47# _0182_ 0.04621f
C32304 _0352_ net112 0
C32305 _0200_ hold6/a_391_47# 0
C32306 _0984_/a_27_47# _0506_/a_299_297# 0
C32307 _0984_/a_193_47# _0506_/a_81_21# 0
C32308 _0223_ _0369_ 0
C32309 _0124_ acc0.A\[25\] 0.28022f
C32310 _0808_/a_585_47# _0091_ 0
C32311 net79 _0091_ 0.00381f
C32312 _0714_/a_51_297# _0999_/a_27_47# 0
C32313 _0439_ _0988_/a_466_413# 0.00108f
C32314 _0242_ net223 0
C32315 _0765_/a_215_47# _0369_ 0.051f
C32316 clknet_1_1__leaf__0463_ net28 0.00183f
C32317 _0352_ acc0.A\[24\] 0.04486f
C32318 _0474_ _0563_/a_51_297# 0
C32319 _0568_/a_109_297# net116 0
C32320 net180 net171 0
C32321 VPWR _0988_/a_466_413# 0.24829f
C32322 _0356_ _0332_ 0.1699f
C32323 _1015_/a_634_159# clknet_1_0__leaf__0457_ 0.01033f
C32324 net125 VPWR 0.56215f
C32325 net36 _0611_/a_68_297# 0.0031f
C32326 _0529_/a_109_297# _0447_ 0
C32327 net145 _0505_/a_27_297# 0
C32328 output66/a_27_47# A[12] 0.03379f
C32329 hold78/a_391_47# _1031_/a_891_413# 0
C32330 _0344_ _1031_/a_634_159# 0
C32331 net168 _1054_/a_891_413# 0
C32332 hold6/a_285_47# _0206_ 0
C32333 VPWR _0953_/a_220_297# 0.00505f
C32334 _0194_ net73 0
C32335 _1056_/a_1059_315# _0186_ 0.03704f
C32336 _0221_ _0345_ 0.12148f
C32337 _1023_/a_561_413# net177 0
C32338 _1023_/a_1059_315# acc0.A\[23\] 0.08418f
C32339 _0616_/a_78_199# net92 0
C32340 comp0.B\[10\] _1043_/a_27_47# 0.00187f
C32341 _0585_/a_27_297# _0171_ 0
C32342 _0294_ _0426_ 0.00273f
C32343 _1016_/a_27_47# _0181_ 0
C32344 _0581_/a_109_297# acc0.A\[19\] 0
C32345 net178 _0350_ 0
C32346 _0504_/a_27_47# clknet_1_0__leaf__0461_ 0
C32347 _0410_ acc0.A\[13\] 0
C32348 _0465_ _0840_/a_150_297# 0
C32349 _1044_/a_193_47# net20 0.03264f
C32350 hold64/a_49_47# acc0.A\[1\] 0
C32351 _0813_/a_109_297# _0345_ 0
C32352 net8 net28 0
C32353 pp[30] _0722_/a_79_21# 0
C32354 _0768_/a_109_297# _0392_ 0
C32355 net155 _0571_/a_373_47# 0
C32356 net89 clknet_0_clk 0
C32357 _0404_ _0799_/a_80_21# 0.12251f
C32358 _0457_ _1015_/a_27_47# 0.03363f
C32359 net131 net20 0
C32360 _0183_ _0721_/a_27_47# 0.04475f
C32361 VPWR _0635_/a_109_297# 0.0038f
C32362 net58 _0840_/a_68_297# 0
C32363 _0456_ clknet_1_0__leaf__0461_ 0.00131f
C32364 _0337_ hold62/a_391_47# 0
C32365 _0130_ _0181_ 0
C32366 _0258_ acc0.A\[6\] 0
C32367 _0481_ _0478_ 0.01161f
C32368 _0380_ _0756_/a_377_297# 0
C32369 _0699_/a_68_297# net94 0
C32370 _1037_/a_27_47# B[6] 0
C32371 clknet_0__0458_ _0839_/a_109_297# 0.00105f
C32372 _0294_ _0185_ 0
C32373 clkbuf_1_0__f__0463_/a_110_47# _0548_/a_240_47# 0
C32374 _1001_/a_466_413# VPWR 0.25162f
C32375 clknet_1_0__leaf__0464_ net9 0.32548f
C32376 net45 _1017_/a_193_47# 0.01025f
C32377 net163 _1031_/a_891_413# 0
C32378 net120 _0131_ 0
C32379 VPWR _1062_/a_634_159# 0.18396f
C32380 _0316_ net244 0.00141f
C32381 _0342_ _0216_ 0.02693f
C32382 _0616_/a_493_297# _0247_ 0
C32383 net145 _0506_/a_81_21# 0.02555f
C32384 _0134_ _0176_ 0
C32385 _1039_/a_193_47# _0172_ 0.00324f
C32386 _1021_/a_27_47# VPWR 0.69941f
C32387 VPWR hold90/a_285_47# 0.26918f
C32388 net193 _0204_ 0
C32389 _1018_/a_1059_315# _0245_ 0
C32390 _0762_/a_79_21# _0762_/a_215_47# 0.04584f
C32391 net167 _0466_ 0.16842f
C32392 hold52/a_49_47# hold52/a_285_47# 0.22264f
C32393 net45 _0241_ 0
C32394 hold20/a_285_47# _1068_/a_891_413# 0.01623f
C32395 hold20/a_391_47# _1068_/a_1059_315# 0.00277f
C32396 _0817_/a_81_21# _0291_ 0
C32397 _0574_/a_109_297# acc0.A\[24\] 0.0072f
C32398 _0347_ net244 0.01521f
C32399 _1041_/a_27_47# net172 0
C32400 net193 hold6/a_391_47# 0
C32401 comp0.B\[7\] _0176_ 0.00204f
C32402 _0846_/a_51_297# clkbuf_0__0458_/a_110_47# 0
C32403 acc0.A\[20\] net87 0
C32404 _0437_ _0619_/a_68_297# 0.02514f
C32405 net84 _0459_ 0
C32406 clknet_1_0__leaf__0463_ hold27/a_49_47# 0.00772f
C32407 _0216_ _0334_ 0
C32408 net53 _0347_ 0.02804f
C32409 _0243_ clknet_1_0__leaf__0457_ 0
C32410 _0395_ _0394_ 0.00431f
C32411 VPWR _0561_/a_512_297# 0.00825f
C32412 _1065_/a_193_47# _1065_/a_381_47# 0.09503f
C32413 _1065_/a_634_159# _1065_/a_891_413# 0.03684f
C32414 _1065_/a_27_47# _1065_/a_561_413# 0.00163f
C32415 net169 net11 0.02413f
C32416 _0183_ _0760_/a_285_47# 0.00603f
C32417 hold85/a_49_47# clknet_1_1__leaf_clk 0.01071f
C32418 net150 _0381_ 0.22551f
C32419 net232 _1066_/a_381_47# 0.11485f
C32420 _0121_ _0120_ 0.00353f
C32421 _0429_ net169 0
C32422 _0998_/a_466_413# _0218_ 0
C32423 _0343_ _0747_/a_79_21# 0
C32424 _1036_/a_1059_315# _1035_/a_193_47# 0.00378f
C32425 _1036_/a_891_413# _1035_/a_27_47# 0.00139f
C32426 _0532_/a_299_297# _0146_ 0.00103f
C32427 net232 net1 0
C32428 A[4] A[8] 0.26864f
C32429 _0853_/a_68_297# _0399_ 0.02182f
C32430 _0707_/a_75_199# _0707_/a_315_47# 0.02023f
C32431 net31 _0548_/a_245_297# 0
C32432 _1033_/a_27_47# net201 0
C32433 _1033_/a_891_413# _0565_/a_240_47# 0
C32434 hold79/a_49_47# _1070_/a_466_413# 0
C32435 _1014_/a_27_47# _1014_/a_466_413# 0.27314f
C32436 _1014_/a_193_47# _1014_/a_634_159# 0.11072f
C32437 net33 hold84/a_49_47# 0.00307f
C32438 net152 _0540_/a_149_47# 0
C32439 _0268_ acc0.A\[15\] 0.01354f
C32440 VPWR _1047_/a_1059_315# 0.41546f
C32441 clknet_1_1__leaf__0460_ _0359_ 0.03309f
C32442 _0627_/a_369_297# clknet_0__0465_ 0
C32443 VPWR _0473_ 1.29782f
C32444 hold3/a_49_47# _0374_ 0
C32445 output55/a_27_47# pp[30] 0
C32446 pp[27] output59/a_27_47# 0
C32447 _1052_/a_27_47# net137 0
C32448 _0239_ clknet_0__0461_ 0
C32449 _0399_ _0252_ 0.00448f
C32450 VPWR _1007_/a_561_413# 0.00345f
C32451 _0341_ _0339_ 0.04027f
C32452 net236 net167 0.00107f
C32453 _0753_/a_79_21# _0230_ 0
C32454 hold34/a_285_47# A[11] 0
C32455 _0312_ _0746_/a_299_297# 0
C32456 net61 hold65/a_391_47# 0.02243f
C32457 _1021_/a_27_47# net48 0
C32458 _0734_/a_377_297# VPWR 0.00367f
C32459 net245 _0410_ 0.00191f
C32460 VPWR clkbuf_1_1__f__0464_/a_110_47# 1.24001f
C32461 _1055_/a_466_413# net16 0.00389f
C32462 _1055_/a_193_47# _0190_ 0
C32463 clknet_1_1__leaf__0465_ _1060_/a_193_47# 0.00165f
C32464 acc0.A\[27\] _0364_ 0
C32465 _0344_ _0345_ 0.00258f
C32466 hold78/a_285_47# _0219_ 0
C32467 _0830_/a_79_21# _0989_/a_27_47# 0.00841f
C32468 _0357_ _0355_ 0
C32469 output52/a_27_47# pp[24] 0.15955f
C32470 _0350_ net110 0
C32471 _1018_/a_634_159# net103 0
C32472 _1000_/a_1059_315# net206 0
C32473 pp[27] _0724_/a_113_297# 0.01886f
C32474 hold41/a_391_47# A[11] 0
C32475 clknet_1_1__leaf__0459_ _0218_ 0.1631f
C32476 clknet_1_1__leaf_clk _1063_/a_975_413# 0
C32477 _0837_/a_585_47# _0085_ 0
C32478 net16 net181 0.00251f
C32479 net112 _1025_/a_466_413# 0
C32480 clkbuf_1_0__f__0463_/a_110_47# net7 0
C32481 _0243_ _1001_/a_1059_315# 0.00373f
C32482 _0088_ _0988_/a_1059_315# 0
C32483 _0959_/a_80_21# control0.sh 0
C32484 _0554_/a_68_297# _0176_ 0
C32485 VPWR _0748_/a_81_21# 0.23732f
C32486 _0343_ _1017_/a_1017_47# 0
C32487 _0375_ _0227_ 0.26502f
C32488 _0151_ hold83/a_285_47# 0.00862f
C32489 _0264_ _0447_ 0
C32490 _1025_/a_466_413# acc0.A\[24\] 0
C32491 _0439_ _0186_ 0.02612f
C32492 clknet_1_0__leaf__0462_ _0753_/a_465_47# 0
C32493 _0693_/a_68_297# _0460_ 0
C32494 VPWR _0186_ 6.69881f
C32495 _0985_/a_891_413# net61 0.01459f
C32496 _1013_/a_891_413# _0339_ 0.00109f
C32497 net25 _1066_/a_193_47# 0
C32498 hold49/a_49_47# VPWR 0.32405f
C32499 clknet_1_0__leaf__0460_ net52 0.0051f
C32500 _0981_/a_27_297# _0981_/a_109_47# 0.00393f
C32501 _0284_ _0281_ 0.39221f
C32502 _0686_/a_219_297# _0219_ 0
C32503 net154 _0193_ 0
C32504 _0457_ _0215_ 0.18791f
C32505 pp[9] clknet_1_1__leaf__0465_ 0.0027f
C32506 _0118_ net211 0
C32507 _0222_ _1022_/a_466_413# 0
C32508 _0855_/a_384_47# net149 0.01033f
C32509 _0481_ _1070_/a_193_47# 0
C32510 VPWR hold19/a_49_47# 0.30705f
C32511 _0854_/a_215_47# _0081_ 0.00423f
C32512 _1037_/a_193_47# _1036_/a_193_47# 0
C32513 _1037_/a_634_159# _1036_/a_27_47# 0
C32514 _1037_/a_27_47# _1036_/a_634_159# 0
C32515 _0082_ _0184_ 0
C32516 _0384_ net92 0
C32517 _0179_ _0268_ 0.01991f
C32518 _0642_/a_27_413# _0435_ 0.00293f
C32519 hold21/a_391_47# net12 0
C32520 _0600_/a_253_297# _0366_ 0
C32521 _0817_/a_81_21# _0290_ 0.00115f
C32522 _0297_ _0668_/a_79_21# 0.03207f
C32523 hold22/a_49_47# clknet_1_1__leaf__0458_ 0.00186f
C32524 _0346_ net79 0.00427f
C32525 _0999_/a_634_159# _0352_ 0.00224f
C32526 _0983_/a_27_47# _0294_ 0
C32527 net78 acc0.A\[10\] 0.00203f
C32528 _0830_/a_510_47# _0087_ 0
C32529 _0251_ _0255_ 0
C32530 _0841_/a_215_47# _0986_/a_193_47# 0
C32531 _0841_/a_79_21# _0986_/a_466_413# 0
C32532 clknet_1_1__leaf__0460_ _1028_/a_466_413# 0
C32533 _0640_/a_109_53# _0255_ 0.14001f
C32534 _0179_ _0090_ 0
C32535 clknet_0__0458_ _0847_/a_109_297# 0
C32536 pp[8] hold35/a_49_47# 0
C32537 net170 _0447_ 0
C32538 _0274_ clknet_0__0465_ 0.43893f
C32539 _1038_/a_1059_315# _0553_/a_240_47# 0
C32540 _1038_/a_27_47# _0174_ 0
C32541 comp0.B\[2\] _1033_/a_27_47# 0.36075f
C32542 net36 _1040_/a_634_159# 0
C32543 hold44/a_285_47# clknet_1_1__leaf__0462_ 0
C32544 _0577_/a_27_297# _1005_/a_891_413# 0
C32545 net190 _1028_/a_27_47# 0.07694f
C32546 _0216_ _1014_/a_193_47# 0
C32547 _0195_ _1014_/a_466_413# 0
C32548 A[13] A[14] 0.17942f
C32549 _0684_/a_145_75# clknet_0__0460_ 0.00165f
C32550 _0180_ _0524_/a_373_47# 0.0019f
C32551 VPWR clknet_0__0462_ 1.95677f
C32552 _0289_ _0294_ 0
C32553 _0292_ _0218_ 0
C32554 output67/a_27_47# _1057_/a_27_47# 0
C32555 hold33/a_49_47# _0176_ 0
C32556 _0845_/a_109_297# _0447_ 0
C32557 net43 _0405_ 0
C32558 _0837_/a_266_47# clknet_0__0465_ 0
C32559 _0340_ net99 0
C32560 _0972_/a_93_21# _0468_ 0.1441f
C32561 control0.state\[0\] hold89/a_49_47# 0.00554f
C32562 net101 _0461_ 0.0219f
C32563 _0179_ net3 0
C32564 _1001_/a_193_47# net87 0.01325f
C32565 acc0.A\[27\] _1010_/a_193_47# 0
C32566 _1018_/a_193_47# net206 0.02183f
C32567 B[8] input7/a_75_212# 0.00436f
C32568 input31/a_75_212# A[15] 0
C32569 _1008_/a_634_159# _1008_/a_1059_315# 0
C32570 _1008_/a_27_47# _1008_/a_381_47# 0.06222f
C32571 _1008_/a_193_47# _1008_/a_891_413# 0.19489f
C32572 _0976_/a_218_374# control0.count\[0\] 0.0094f
C32573 net169 clknet_1_1__leaf__0458_ 0
C32574 _0290_ _0084_ 0.00139f
C32575 _0172_ clkbuf_0__0464_/a_110_47# 0.15167f
C32576 _0092_ acc0.A\[13\] 0
C32577 hold56/a_49_47# comp0.B\[0\] 0.01009f
C32578 _0718_/a_47_47# _1011_/a_1059_315# 0
C32579 _0718_/a_285_47# _1011_/a_193_47# 0
C32580 output43/a_27_47# _0995_/a_634_159# 0
C32581 _1020_/a_381_47# _1020_/a_561_413# 0.00123f
C32582 _1020_/a_891_413# _1020_/a_975_413# 0.00851f
C32583 acc0.A\[0\] _0264_ 0
C32584 net53 _1025_/a_27_47# 0.01551f
C32585 acc0.A\[23\] _0219_ 0.04029f
C32586 _1035_/a_891_413# comp0.B\[3\] 0.00352f
C32587 net103 _0114_ 0.03134f
C32588 _0559_/a_51_297# _0561_/a_149_47# 0
C32589 _1035_/a_27_47# _0474_ 0
C32590 _0559_/a_149_47# _0561_/a_51_297# 0
C32591 _0175_ _0213_ 0.08205f
C32592 net58 _0255_ 0.00409f
C32593 _0239_ _0607_/a_373_47# 0
C32594 _0229_ _0234_ 0.00378f
C32595 _0724_/a_113_297# _0724_/a_199_47# 0
C32596 _0255_ hold7/a_49_47# 0
C32597 output59/a_27_47# _0216_ 0.02704f
C32598 net59 net57 0
C32599 _0230_ _0732_/a_80_21# 0
C32600 net216 clkbuf_1_0__f__0460_/a_110_47# 0.00871f
C32601 hold28/a_285_47# acc0.A\[3\] 0.052f
C32602 hold85/a_285_47# VPWR 0.29374f
C32603 acc0.A\[27\] _1009_/a_634_159# 0
C32604 clknet_0__0458_ _0986_/a_634_159# 0.00208f
C32605 net64 pp[1] 0
C32606 _0343_ output58/a_27_47# 0
C32607 net55 clknet_1_1__leaf__0460_ 0.37593f
C32608 _0183_ clkbuf_1_0__f__0461_/a_110_47# 0.02233f
C32609 clknet_0__0457_ _1014_/a_634_159# 0
C32610 hold34/a_285_47# net66 0.00344f
C32611 pp[8] A[9] 0.69757f
C32612 control0.sh _0173_ 0.5998f
C32613 net216 _0250_ 0.0473f
C32614 _0513_/a_81_21# net3 0
C32615 _1054_/a_27_47# _0518_/a_109_297# 0
C32616 _1054_/a_193_47# _0518_/a_27_297# 0
C32617 _0502_/a_27_47# _0465_ 0.02229f
C32618 _1013_/a_381_47# net99 0
C32619 hold14/a_391_47# VPWR 0.17493f
C32620 _0275_ _0815_/a_113_297# 0
C32621 _1032_/a_27_47# comp0.B\[0\] 0
C32622 _0313_ _0367_ 0.28594f
C32623 _1041_/a_1059_315# _0172_ 0.00335f
C32624 _1041_/a_634_159# _0137_ 0
C32625 _0404_ _0997_/a_1059_315# 0
C32626 _0997_/a_27_47# _0345_ 0.03406f
C32627 _0483_ net159 0
C32628 pp[28] _0195_ 0.00251f
C32629 _0109_ hold80/a_391_47# 0
C32630 _0992_/a_1059_315# _0345_ 0
C32631 _0230_ clkbuf_1_0__f__0460_/a_110_47# 0
C32632 net111 _0352_ 0
C32633 hold94/a_285_47# _0345_ 0.02977f
C32634 hold21/a_285_47# A[8] 0.08117f
C32635 _0216_ _0724_/a_113_297# 0.00171f
C32636 _0570_/a_109_297# _0352_ 0
C32637 _0991_/a_466_413# acc0.A\[15\] 0
C32638 _0984_/a_193_47# _0184_ 0
C32639 _0346_ hold2/a_285_47# 0.00141f
C32640 _0476_ _0163_ 0
C32641 _0992_/a_381_47# _0295_ 0
C32642 _0982_/a_27_47# net234 0
C32643 net102 _0582_/a_27_297# 0.00162f
C32644 _0982_/a_1059_315# _0855_/a_299_297# 0
C32645 _0982_/a_891_413# _0855_/a_81_21# 0
C32646 _0212_ _0175_ 0.0228f
C32647 net161 input24/a_75_212# 0.00121f
C32648 _1010_/a_193_47# _0110_ 0
C32649 _0578_/a_109_297# _0217_ 0.01259f
C32650 _0093_ _0411_ 0.001f
C32651 VPWR _0497_/a_68_297# 0.14718f
C32652 clknet_1_1__leaf_clk net17 0.20295f
C32653 _0596_/a_59_75# _0369_ 0
C32654 _0781_/a_68_297# _0369_ 0
C32655 net168 hold22/a_391_47# 0.05018f
C32656 done control0.count\[2\] 0
C32657 _1000_/a_381_47# _0352_ 0.01924f
C32658 _1000_/a_592_47# _0347_ 0
C32659 _0576_/a_109_47# clknet_1_0__leaf__0460_ 0
C32660 _0701_/a_80_21# _0350_ 0.01995f
C32661 _0602_/a_113_47# _0219_ 0
C32662 net210 _0124_ 0.02561f
C32663 net155 _0216_ 0.86826f
C32664 net44 _1017_/a_891_413# 0
C32665 clknet_1_0__leaf__0462_ clknet_0__0460_ 0
C32666 hold13/a_285_47# VPWR 0.27737f
C32667 _1016_/a_27_47# clknet_1_1__leaf__0461_ 0.08368f
C32668 net72 acc0.A\[6\] 0
C32669 _0820_/a_79_21# net142 0
C32670 net46 pp[23] 0.00111f
C32671 pp[19] net51 0
C32672 VPWR _1017_/a_193_47# 0.28068f
C32673 _0739_/a_215_47# hold50/a_285_47# 0
C32674 _0432_ _0445_ 0
C32675 _1037_/a_27_47# comp0.B\[5\] 0.00387f
C32676 _0378_ _1005_/a_27_47# 0
C32677 clk clkbuf_1_0__f_clk/a_110_47# 0
C32678 clkbuf_0_clk/a_110_47# clknet_0_clk 1.73133f
C32679 _0984_/a_381_47# net229 0
C32680 _0316_ clkbuf_1_1__f__0462_/a_110_47# 0.04417f
C32681 _0548_/a_245_297# _0548_/a_240_47# 0
C32682 VPWR _1060_/a_592_47# 0
C32683 clkload3/Y net103 0
C32684 _1015_/a_193_47# net149 0
C32685 _1056_/a_634_159# A[10] 0
C32686 _1043_/a_193_47# net153 0
C32687 _0177_ _0171_ 0.0017f
C32688 _0241_ VPWR 0.45857f
C32689 clknet_0_clk _1063_/a_634_159# 0
C32690 net145 _0184_ 0.04491f
C32691 clkbuf_1_1__f__0462_/a_110_47# _0347_ 0.03273f
C32692 net14 net140 0
C32693 acc0.A\[4\] _0197_ 0
C32694 VPWR _1050_/a_634_159# 0.18321f
C32695 clknet_1_0__leaf__0459_ hold19/a_49_47# 0.03769f
C32696 net157 _1047_/a_1017_47# 0
C32697 _0216_ _0240_ 0.00443f
C32698 hold21/a_391_47# pp[5] 0
C32699 acc0.A\[14\] _0998_/a_891_413# 0
C32700 _0252_ _0619_/a_68_297# 0
C32701 _0216_ _0369_ 0.11392f
C32702 VPWR _0958_/a_27_47# 0.39047f
C32703 hold45/a_285_47# net192 0.02539f
C32704 _1010_/a_27_47# _1010_/a_634_159# 0.14145f
C32705 _0179_ _0991_/a_466_413# 0
C32706 clknet_0__0457_ _0216_ 0.25669f
C32707 _0644_/a_377_297# net42 0.00324f
C32708 _0644_/a_47_47# acc0.A\[15\] 0.06276f
C32709 _0348_ _1011_/a_891_413# 0
C32710 _0670_/a_297_297# _0302_ 0
C32711 _0183_ _0182_ 0.02149f
C32712 _0784_/a_113_47# acc0.A\[15\] 0
C32713 net57 _0335_ 0.19512f
C32714 _0198_ _1048_/a_634_159# 0
C32715 _0536_/a_512_297# net157 0.00203f
C32716 _0618_/a_79_21# _0350_ 0.0015f
C32717 VPWR _0973_/a_109_297# 0.19654f
C32718 hold96/a_285_47# _0216_ 0.068f
C32719 _0195_ _0852_/a_285_47# 0
C32720 _1002_/a_27_47# _0217_ 0.02803f
C32721 _1002_/a_193_47# net150 0
C32722 _0746_/a_81_21# _0746_/a_384_47# 0.00138f
C32723 input21/a_75_212# input32/a_75_212# 0
C32724 net76 _0181_ 0
C32725 hold88/a_49_47# _0990_/a_193_47# 0
C32726 hold88/a_285_47# _0990_/a_27_47# 0
C32727 _0749_/a_299_297# _1006_/a_193_47# 0
C32728 _1020_/a_466_413# _0461_ 0
C32729 _1018_/a_381_47# _0347_ 0
C32730 _0309_ clknet_0__0461_ 0
C32731 net222 acc0.A\[15\] 0.02137f
C32732 _0280_ _0651_/a_113_47# 0
C32733 net36 control0.reset 0
C32734 net191 hold50/a_49_47# 0
C32735 acc0.A\[12\] hold70/a_285_47# 0
C32736 hold91/a_49_47# net6 0
C32737 _0421_ _0345_ 0.0101f
C32738 _0106_ net244 0
C32739 net212 _0434_ 0
C32740 _1000_/a_1059_315# _0773_/a_35_297# 0
C32741 _1000_/a_634_159# _0773_/a_285_297# 0
C32742 _0575_/a_27_297# _0347_ 0
C32743 _1009_/a_27_47# _1009_/a_1059_315# 0.04875f
C32744 _1009_/a_193_47# _1009_/a_466_413# 0.08261f
C32745 _0698_/a_199_47# acc0.A\[28\] 0
C32746 VPWR _0518_/a_109_47# 0
C32747 net36 _1061_/a_891_413# 0
C32748 _0376_ net49 0
C32749 _0576_/a_27_297# _0576_/a_373_47# 0.01338f
C32750 _0645_/a_47_47# _1059_/a_193_47# 0
C32751 _0645_/a_377_297# _1059_/a_27_47# 0
C32752 clknet_1_0__leaf__0460_ hold93/a_49_47# 0
C32753 hold100/a_49_47# VPWR 0.2696f
C32754 net32 _0542_/a_51_297# 0
C32755 net139 hold83/a_391_47# 0.00374f
C32756 _0387_ net43 0
C32757 clknet_1_1__leaf__0460_ _0325_ 0.00546f
C32758 _0236_ clkbuf_1_0__f__0460_/a_110_47# 0
C32759 hold35/a_391_47# _0186_ 0
C32760 _1065_/a_193_47# control0.reset 0.00112f
C32761 hold5/a_285_47# net198 0
C32762 hold5/a_49_47# net18 0
C32763 acc0.A\[17\] _0347_ 0.06654f
C32764 VPWR _0132_ 0.52626f
C32765 net232 control0.sh 0.00677f
C32766 _0982_/a_193_47# VPWR 0.30516f
C32767 _0476_ _1066_/a_27_47# 0.03726f
C32768 net213 _1005_/a_193_47# 0
C32769 _0260_ _0449_ 0.04807f
C32770 _1036_/a_466_413# net121 0.02244f
C32771 _1036_/a_634_159# _0133_ 0
C32772 net111 _1025_/a_466_413# 0
C32773 net7 _0548_/a_245_297# 0.0012f
C32774 _0236_ _0250_ 0
C32775 _0305_ clkbuf_0__0459_/a_110_47# 0.02011f
C32776 net1 _0162_ 0
C32777 net89 _0228_ 0
C32778 _0819_/a_299_297# _0346_ 0.01866f
C32779 _0707_/a_208_47# _0339_ 0
C32780 _0182_ acc0.A\[15\] 0.12772f
C32781 comp0.B\[1\] _0565_/a_149_47# 0.00139f
C32782 hold79/a_49_47# _0168_ 0.01384f
C32783 hold79/a_391_47# VPWR 0.18127f
C32784 comp0.B\[11\] _1042_/a_1017_47# 0.00125f
C32785 _0390_ _0241_ 0.00922f
C32786 _1014_/a_193_47# net100 0.03103f
C32787 _1014_/a_1059_315# _1014_/a_1017_47# 0
C32788 _0959_/a_80_21# _0955_/a_32_297# 0.00194f
C32789 _1071_/a_634_159# _1071_/a_381_47# 0
C32790 net59 _1010_/a_1059_315# 0
C32791 _0996_/a_27_47# net238 0.0455f
C32792 pp[30] acc0.A\[30\] 0.05641f
C32793 _1015_/a_891_413# _0208_ 0.04754f
C32794 _0333_ hold62/a_391_47# 0
C32795 _0327_ _0729_/a_68_297# 0.00832f
C32796 hold96/a_285_47# hold96/a_391_47# 0.41909f
C32797 _0985_/a_592_47# _0458_ 0.00116f
C32798 _1013_/a_193_47# net42 0
C32799 net54 _0687_/a_145_75# 0
C32800 _0852_/a_35_297# _0852_/a_285_47# 0.00723f
C32801 _0717_/a_209_297# pp[29] 0
C32802 net168 _0255_ 0
C32803 _0179_ _0401_ 0.01739f
C32804 _0179_ acc0.A\[5\] 0.00491f
C32805 _0983_/a_193_47# acc0.A\[14\] 0
C32806 _0251_ _0830_/a_215_47# 0
C32807 _0343_ _0792_/a_209_47# 0
C32808 hold53/a_49_47# VPWR 0.36575f
C32809 _1035_/a_634_159# net26 0.01568f
C32810 hold39/a_49_47# hold39/a_391_47# 0.00188f
C32811 _0195_ _0844_/a_297_47# 0
C32812 _0175_ _0161_ 0
C32813 VPWR _0200_ 0.73782f
C32814 clknet_1_1__leaf__0460_ _0238_ 0.18691f
C32815 VPWR _0410_ 0.5118f
C32816 _1039_/a_1017_47# comp0.B\[6\] 0
C32817 _0670_/a_297_297# net6 0.0082f
C32818 _0439_ net62 0.02475f
C32819 net179 net16 0.04052f
C32820 clknet_0__0457_ net247 0
C32821 _0216_ _1024_/a_27_47# 0
C32822 net65 _0437_ 0.51302f
C32823 _0809_/a_81_21# _0345_ 0.01608f
C32824 _0087_ _0989_/a_193_47# 0.18376f
C32825 _0437_ _0989_/a_466_413# 0.01657f
C32826 _0856_/a_79_21# _0447_ 0
C32827 _0305_ _1059_/a_381_47# 0
C32828 VPWR net62 1.10412f
C32829 _0179_ net222 0
C32830 hold98/a_285_47# pp[14] 0.02505f
C32831 net45 net219 0.25431f
C32832 VPWR _0450_ 0.38879f
C32833 _1015_/a_1059_315# net17 0
C32834 _0186_ _0523_/a_81_21# 0.07419f
C32835 VPWR comp0.B\[8\] 0.67055f
C32836 _1026_/a_1017_47# acc0.A\[25\] 0
C32837 _0295_ _0809_/a_384_47# 0.00884f
C32838 net36 _1039_/a_891_413# 0.04152f
C32839 _0787_/a_80_21# _0808_/a_81_21# 0.00103f
C32840 _0195_ _1048_/a_1059_315# 0.01431f
C32841 _0100_ _1067_/a_1059_315# 0
C32842 net88 _1067_/a_891_413# 0
C32843 _1042_/a_1059_315# _0542_/a_51_297# 0
C32844 _1002_/a_193_47# control0.add 0
C32845 _1012_/a_1059_315# _0352_ 0.01376f
C32846 _1012_/a_561_413# _0347_ 0
C32847 _0608_/a_109_297# _0240_ 0
C32848 clknet_1_0__leaf__0460_ hold94/a_391_47# 0.00137f
C32849 net182 _0186_ 0
C32850 acc0.A\[25\] _0122_ 0
C32851 clknet_1_1__leaf__0462_ _0219_ 0.46075f
C32852 _0343_ _1016_/a_381_47# 0.00226f
C32853 _1033_/a_193_47# _0215_ 0.03929f
C32854 clknet_1_0__leaf__0459_ _1017_/a_193_47# 0.00788f
C32855 _0609_/a_109_297# _0462_ 0
C32856 hold30/a_49_47# _0375_ 0
C32857 _0083_ net233 0
C32858 _0369_ _0825_/a_68_297# 0
C32859 hold25/a_285_47# net7 0
C32860 acc0.A\[31\] _0340_ 0.13274f
C32861 _0728_/a_59_75# clknet_1_1__leaf__0462_ 0
C32862 _0433_ _0987_/a_1059_315# 0
C32863 _1052_/a_381_47# _0180_ 0
C32864 hold54/a_285_47# comp0.B\[0\] 0
C32865 _1016_/a_891_413# acc0.A\[17\] 0
C32866 _0241_ clknet_1_0__leaf__0459_ 0.02627f
C32867 hold89/a_49_47# _0478_ 0
C32868 _0222_ net151 0
C32869 _0456_ _0112_ 0
C32870 _0225_ _0606_/a_215_297# 0.19883f
C32871 _0481_ VPWR 0.85253f
C32872 _0179_ _0182_ 0.00122f
C32873 hold20/a_391_47# control0.count\[3\] 0
C32874 hold20/a_49_47# _0483_ 0
C32875 hold42/a_49_47# pp[10] 0.00167f
C32876 clknet_1_1__leaf__0459_ net228 0.02848f
C32877 _0255_ _0831_/a_285_297# 0
C32878 net9 clkbuf_1_0__f__0464_/a_110_47# 0.03391f
C32879 net62 output62/a_27_47# 0.22668f
C32880 _0459_ acc0.A\[18\] 0.05519f
C32881 net85 _0352_ 0.02994f
C32882 _1030_/a_193_47# hold62/a_49_47# 0
C32883 _1030_/a_27_47# hold62/a_285_47# 0.00329f
C32884 _0305_ _0731_/a_81_21# 0
C32885 input28/a_75_212# net28 0.10856f
C32886 _0985_/a_27_47# _0350_ 0.00204f
C32887 _0975_/a_59_75# _0468_ 0
C32888 _0498_/a_240_47# _0159_ 0.00162f
C32889 net22 _0205_ 0.04089f
C32890 _0375_ _0352_ 0.02071f
C32891 _0445_ _0986_/a_381_47# 0
C32892 _0084_ _0986_/a_1059_315# 0
C32893 _0579_/a_27_297# _0457_ 0
C32894 net10 _0142_ 0
C32895 _0227_ VPWR 1.0782f
C32896 _0108_ acc0.A\[29\] 0
C32897 hold97/a_285_47# acc0.A\[27\] 0.00416f
C32898 hold96/a_391_47# _1024_/a_27_47# 0
C32899 hold96/a_285_47# _1024_/a_193_47# 0
C32900 hold96/a_49_47# _1024_/a_634_159# 0
C32901 _0258_ _0826_/a_219_297# 0
C32902 _0551_/a_27_47# _0565_/a_51_297# 0
C32903 _0224_ net49 0
C32904 net14 input14/a_75_212# 0.1077f
C32905 net168 A[7] 0
C32906 clknet_1_0__leaf__0462_ output46/a_27_47# 0.00139f
C32907 net197 net114 0.24342f
C32908 _0266_ net149 0
C32909 net193 VPWR 0.178f
C32910 clknet_1_1__leaf__0462_ _1008_/a_634_159# 0.00188f
C32911 _0955_/a_32_297# _0173_ 0
C32912 comp0.B\[3\] _0561_/a_512_297# 0
C32913 comp0.B\[5\] _0561_/a_51_297# 0.00131f
C32914 _1032_/a_193_47# _0565_/a_240_47# 0
C32915 _0165_ clknet_1_1__leaf_clk 0.04127f
C32916 VPWR _1046_/a_466_413# 0.24057f
C32917 _1022_/a_193_47# _1022_/a_891_413# 0.19549f
C32918 _1022_/a_27_47# _1022_/a_381_47# 0.06222f
C32919 _1022_/a_634_159# _1022_/a_1059_315# 0
C32920 acc0.A\[31\] _1013_/a_381_47# 0
C32921 net162 _1013_/a_1059_315# 0
C32922 net231 _0468_ 0
C32923 _0856_/a_79_21# acc0.A\[0\] 0.02062f
C32924 _0717_/a_80_21# acc0.A\[30\] 0
C32925 _1003_/a_1017_47# clknet_1_0__leaf__0460_ 0
C32926 _0686_/a_27_53# _0318_ 0.03507f
C32927 _1059_/a_1017_47# acc0.A\[15\] 0
C32928 clknet_1_0__leaf__0463_ _0205_ 0
C32929 _0855_/a_81_21# clkbuf_0__0457_/a_110_47# 0
C32930 _1008_/a_891_413# _0318_ 0
C32931 clknet_0__0463_ clknet_1_1__leaf__0463_ 0.18932f
C32932 _0272_ _0986_/a_193_47# 0
C32933 net211 _1001_/a_27_47# 0.09091f
C32934 _0957_/a_114_297# _0474_ 0.01124f
C32935 _1018_/a_592_47# _0116_ 0
C32936 _0957_/a_304_297# comp0.B\[6\] 0.00137f
C32937 hold38/a_391_47# clknet_1_1__leaf__0463_ 0.00424f
C32938 _0339_ acc0.A\[30\] 0.37201f
C32939 _1055_/a_466_413# _1055_/a_561_413# 0.00772f
C32940 _1055_/a_634_159# _1055_/a_975_413# 0
C32941 _0505_/a_27_297# net6 0.19125f
C32942 hold74/a_391_47# clknet_0__0461_ 0
C32943 VPWR _0759_/a_113_47# 0
C32944 hold43/a_49_47# hold43/a_285_47# 0.22264f
C32945 hold24/a_285_47# hold24/a_391_47# 0.41909f
C32946 _1020_/a_1017_47# _0118_ 0
C32947 _0771_/a_215_297# _0771_/a_382_47# 0.01048f
C32948 _0133_ comp0.B\[5\] 0.02622f
C32949 _0559_/a_149_47# _0208_ 0.02272f
C32950 hold14/a_391_47# _1036_/a_27_47# 0
C32951 hold14/a_285_47# _1036_/a_193_47# 0
C32952 hold14/a_49_47# _1036_/a_634_159# 0
C32953 _0466_ _1063_/a_27_47# 0
C32954 net89 hold12/a_285_47# 0.01395f
C32955 _1003_/a_634_159# _1003_/a_381_47# 0
C32956 hold97/a_285_47# _0364_ 0.0018f
C32957 net166 net165 0
C32958 clkload2/Y _0142_ 0.00175f
C32959 _1001_/a_891_413# _0399_ 0
C32960 VPWR _0687_/a_59_75# 0.2127f
C32961 hold64/a_49_47# _0216_ 0.0465f
C32962 _0292_ net228 0
C32963 _0626_/a_68_297# _0346_ 0
C32964 _0466_ _0974_/a_448_47# 0
C32965 clknet_0__0457_ net100 0.04099f
C32966 clknet_0__0463_ net8 0.62019f
C32967 net185 _0955_/a_220_297# 0.00107f
C32968 _0558_/a_68_297# comp0.B\[5\] 0.00301f
C32969 _0212_ _0955_/a_114_297# 0
C32970 hold55/a_391_47# _0584_/a_109_297# 0
C32971 _0227_ net48 0.05101f
C32972 _0176_ _0203_ 0.08501f
C32973 net87 _0208_ 0
C32974 _0233_ _0238_ 0
C32975 _0346_ _0301_ 0.25699f
C32976 net22 _1042_/a_193_47# 0
C32977 VPWR _0747_/a_215_47# 0.00204f
C32978 _1054_/a_193_47# _0191_ 0.03352f
C32979 _1054_/a_466_413# net15 0
C32980 _0556_/a_68_297# net28 0.00569f
C32981 _0556_/a_150_297# B[5] 0
C32982 _0830_/a_79_21# clknet_1_1__leaf__0458_ 0.00654f
C32983 _0181_ clkbuf_0__0459_/a_110_47# 0.00555f
C32984 _0997_/a_561_413# _0219_ 0
C32985 _0764_/a_299_297# _0384_ 0.10107f
C32986 _0465_ _0843_/a_150_297# 0
C32987 _0844_/a_79_21# _0844_/a_382_297# 0.00145f
C32988 _1004_/a_1059_315# _0347_ 0.00325f
C32989 _1004_/a_193_47# _0352_ 0.01747f
C32990 _1004_/a_27_47# _0102_ 0.12289f
C32991 _0855_/a_384_47# net206 0
C32992 hold59/a_49_47# _0459_ 0
C32993 net53 _0314_ 0.22823f
C32994 net197 _0365_ 0.02844f
C32995 _0534_/a_81_21# _0531_/a_27_297# 0
C32996 clknet_1_1__leaf__0461_ _0400_ 0
C32997 _0089_ acc0.A\[15\] 0
C32998 _0441_ acc0.A\[5\] 0
C32999 _0966_/a_27_47# clk 0.00265f
C33000 _1054_/a_466_413# _1053_/a_1059_315# 0
C33001 _0506_/a_81_21# net6 0.00107f
C33002 VPWR hold9/a_391_47# 0.16509f
C33003 _0799_/a_209_297# _0799_/a_303_47# 0
C33004 _0982_/a_975_413# _0456_ 0.00116f
C33005 net102 _0115_ 0.06181f
C33006 _1012_/a_27_47# _0350_ 0
C33007 _0222_ _0378_ 0.0662f
C33008 _0330_ _0350_ 0.07125f
C33009 _0467_ _0950_/a_75_212# 0.011f
C33010 VPWR _0987_/a_634_159# 0.20496f
C33011 _0271_ _0636_/a_59_75# 0
C33012 _1024_/a_27_47# _1024_/a_193_47# 0.97441f
C33013 _1058_/a_1059_315# net189 0.00903f
C33014 _0276_ _0788_/a_68_297# 0
C33015 _0557_/a_51_297# net160 0.07877f
C33016 net48 _0759_/a_113_47# 0
C33017 _0370_ _0250_ 0.30267f
C33018 _0516_/a_109_47# _0186_ 0.00145f
C33019 hold64/a_285_47# clknet_0__0457_ 0.00291f
C33020 _0218_ _0095_ 0
C33021 net45 _0352_ 0.01272f
C33022 VPWR input12/a_75_212# 0.19472f
C33023 _0464_ net133 0
C33024 _1000_/a_634_159# _0244_ 0.0019f
C33025 _1000_/a_27_47# _0388_ 0.012f
C33026 _1000_/a_193_47# _0386_ 0.00701f
C33027 VPWR _1029_/a_634_159# 0.19626f
C33028 _0294_ _0462_ 0.03159f
C33029 _0367_ _0321_ 0
C33030 hold59/a_285_47# clknet_1_0__leaf__0461_ 0.00582f
C33031 _0128_ _0336_ 0.009f
C33032 _0982_/a_193_47# _0453_ 0
C33033 _0982_/a_1059_315# _0452_ 0.01413f
C33034 clkbuf_0__0460_/a_110_47# _0367_ 0.00101f
C33035 hold61/a_49_47# hold61/a_391_47# 0.00188f
C33036 clknet_1_0__leaf_clk _1064_/a_381_47# 0
C33037 _1048_/a_634_159# _1048_/a_466_413# 0.23992f
C33038 _1048_/a_193_47# _1048_/a_1059_315# 0.03405f
C33039 _1048_/a_27_47# _1048_/a_891_413# 0.03224f
C33040 net211 _0459_ 0.02487f
C33041 comp0.B\[0\] _0950_/a_75_212# 0
C33042 _0348_ output56/a_27_47# 0
C33043 _0398_ _0796_/a_79_21# 0
C33044 _1037_/a_1017_47# comp0.B\[6\] 0
C33045 _0607_/a_27_297# _0780_/a_35_297# 0
C33046 _0350_ _0242_ 0.40163f
C33047 VPWR net25 1.24491f
C33048 _0563_/a_240_47# _0214_ 0
C33049 _0846_/a_51_297# _0447_ 0.01513f
C33050 _0339_ _0779_/a_79_21# 0
C33051 _0555_/a_149_47# VPWR 0.00856f
C33052 _0312_ _1007_/a_634_159# 0
C33053 _0092_ VPWR 0.34253f
C33054 _0713_/a_27_47# net149 0
C33055 hold11/a_49_47# hold11/a_391_47# 0.00188f
C33056 _0680_/a_80_21# clkbuf_0__0460_/a_110_47# 0
C33057 init B[15] 0
C33058 _0083_ hold23/a_49_47# 0
C33059 hold59/a_391_47# net47 0.02018f
C33060 _0243_ _0246_ 0.0396f
C33061 _0337_ _0334_ 0
C33062 clkbuf_1_1__f__0462_/a_110_47# _0106_ 0
C33063 hold55/a_391_47# VPWR 0.18581f
C33064 _0518_/a_27_297# acc0.A\[6\] 0.06173f
C33065 VPWR net136 0.43128f
C33066 net36 _1041_/a_975_413# 0
C33067 hold76/a_49_47# hold76/a_391_47# 0.00188f
C33068 _0349_ _0722_/a_215_47# 0.05119f
C33069 VPWR _0477_ 0.398f
C33070 _1010_/a_891_413# _1010_/a_975_413# 0.00851f
C33071 _1010_/a_27_47# net96 0.2288f
C33072 _1010_/a_381_47# _1010_/a_561_413# 0.00123f
C33073 _0179_ _0089_ 0
C33074 clknet_1_0__leaf__0462_ _1004_/a_1017_47# 0
C33075 _0153_ net66 0
C33076 _1056_/a_891_413# _0514_/a_27_297# 0.01252f
C33077 _1056_/a_1059_315# _0514_/a_109_297# 0
C33078 hold6/a_49_47# _0546_/a_149_47# 0
C33079 _0130_ _1015_/a_27_47# 0
C33080 hold55/a_49_47# _1015_/a_891_413# 0.01135f
C33081 hold55/a_285_47# _1015_/a_1059_315# 0.00197f
C33082 hold92/a_49_47# _0219_ 0.0135f
C33083 _1040_/a_634_159# _1040_/a_975_413# 0
C33084 _1040_/a_466_413# _1040_/a_561_413# 0.00772f
C33085 _0587_/a_27_47# _0352_ 0
C33086 net69 net146 0
C33087 _0146_ _1048_/a_1017_47# 0.00109f
C33088 net232 _0955_/a_32_297# 0
C33089 _0432_ _0440_ 0
C33090 _0443_ _0441_ 0
C33091 hold19/a_391_47# _0399_ 0
C33092 _0144_ net157 0.44257f
C33093 net135 net132 0.00186f
C33094 _1072_/a_27_47# _1072_/a_193_47# 0.96976f
C33095 hold88/a_49_47# clknet_1_1__leaf__0465_ 0.00433f
C33096 _0216_ _1027_/a_1059_315# 0.0666f
C33097 _0853_/a_68_297# _0346_ 0.03868f
C33098 VPWR _1019_/a_466_413# 0.24163f
C33099 _0273_ _0829_/a_109_297# 0
C33100 comp0.B\[7\] net28 0
C33101 control0.state\[0\] _0469_ 0.0017f
C33102 _0749_/a_81_21# net92 0
C33103 _0635_/a_109_297# _0345_ 0
C33104 _1014_/a_27_47# clkbuf_1_1__f__0457_/a_110_47# 0
C33105 _0118_ _0461_ 0.00435f
C33106 acc0.A\[14\] _0996_/a_891_413# 0.01932f
C33107 _0537_/a_150_297# _1045_/a_193_47# 0
C33108 net45 _1016_/a_975_413# 0
C33109 _1067_/a_193_47# _1067_/a_592_47# 0
C33110 _1067_/a_466_413# _1067_/a_561_413# 0.00772f
C33111 _1067_/a_634_159# _1067_/a_975_413# 0
C33112 net9 _0987_/a_561_413# 0
C33113 control0.state\[1\] _0468_ 0.3834f
C33114 hold1/a_285_47# net154 0
C33115 _0821_/a_113_47# acc0.A\[7\] 0
C33116 _1001_/a_466_413# _0345_ 0.01705f
C33117 _0251_ _0989_/a_27_47# 0.0046f
C33118 _0800_/a_149_47# _0410_ 0
C33119 _1002_/a_27_47# _0235_ 0
C33120 hold35/a_49_47# A[10] 0.04165f
C33121 hold12/a_49_47# net35 0.32121f
C33122 _1071_/a_193_47# _0169_ 0.23007f
C33123 _1050_/a_193_47# _0172_ 0
C33124 acc0.A\[1\] net165 0.0012f
C33125 _0985_/a_1059_315# _0529_/a_27_297# 0.00131f
C33126 _0985_/a_466_413# _0529_/a_109_297# 0
C33127 net38 net246 0.23204f
C33128 net199 _0352_ 0
C33129 hold90/a_285_47# _0345_ 0.00863f
C33130 VPWR net219 0.62299f
C33131 _1009_/a_891_413# _1009_/a_1017_47# 0.00617f
C33132 net65 _0252_ 0.14423f
C33133 _0717_/a_80_21# _0717_/a_209_47# 0.01013f
C33134 _0252_ _0989_/a_466_413# 0.03408f
C33135 net65 _0989_/a_381_47# 0
C33136 _0588_/a_113_47# _0395_ 0
C33137 control0.state\[1\] _1002_/a_193_47# 0.00252f
C33138 _0989_/a_1059_315# _0989_/a_891_413# 0.31086f
C33139 _0989_/a_193_47# _0989_/a_975_413# 0
C33140 _0989_/a_466_413# _0989_/a_381_47# 0.03733f
C33141 _0997_/a_27_47# _0997_/a_193_47# 0.95992f
C33142 _1020_/a_27_47# clknet_1_0__leaf__0461_ 0
C33143 comp0.B\[4\] _0957_/a_32_297# 0
C33144 clknet_1_0__leaf__0462_ hold29/a_391_47# 0.01013f
C33145 net190 _0350_ 0
C33146 _0697_/a_80_21# clknet_0__0462_ 0
C33147 comp0.B\[15\] net201 0.17119f
C33148 _0181_ _0986_/a_193_47# 0.00139f
C33149 _0544_/a_51_297# _1042_/a_634_159# 0.00153f
C33150 _0992_/a_1059_315# _0992_/a_891_413# 0.31086f
C33151 _0992_/a_193_47# _0992_/a_975_413# 0
C33152 _0992_/a_466_413# _0992_/a_381_47# 0.03733f
C33153 net161 net121 0.22698f
C33154 _0315_ _1009_/a_193_47# 0
C33155 _0718_/a_47_47# acc0.A\[30\] 0
C33156 comp0.B\[4\] net23 0
C33157 VPWR _1045_/a_193_47# 0.29952f
C33158 acc0.A\[16\] net43 0.49616f
C33159 _0402_ _0808_/a_81_21# 0.0855f
C33160 VPWR _1053_/a_975_413# 0.00477f
C33161 _0125_ _1027_/a_561_413# 0
C33162 acc0.A\[27\] _1027_/a_1017_47# 0
C33163 net54 _0739_/a_510_47# 0.00108f
C33164 _0355_ _1029_/a_1059_315# 0
C33165 _0109_ _1029_/a_27_47# 0
C33166 acc0.A\[1\] acc0.A\[19\] 0.00711f
C33167 _1014_/a_975_413# acc0.A\[0\] 0.00142f
C33168 hold94/a_285_47# hold94/a_391_47# 0.41909f
C33169 _0263_ _0219_ 0.02303f
C33170 clkload4/Y _0219_ 0
C33171 net187 _0181_ 0
C33172 _0963_/a_35_297# _0466_ 0
C33173 hold10/a_391_47# _0465_ 0.00648f
C33174 _0983_/a_193_47# _0116_ 0
C33175 hold54/a_391_47# _0565_/a_240_47# 0
C33176 _1061_/a_193_47# _1061_/a_1059_315# 0.03414f
C33177 _1061_/a_27_47# _1061_/a_891_413# 0.03224f
C33178 _1061_/a_634_159# _1061_/a_466_413# 0.23992f
C33179 _0680_/a_80_21# _1009_/a_27_47# 0
C33180 _0742_/a_384_47# _0360_ 0
C33181 _0458_ acc0.A\[3\] 0.00774f
C33182 net66 _0990_/a_27_47# 0.02607f
C33183 net21 _0541_/a_68_297# 0.00552f
C33184 pp[21] VPWR 0.20649f
C33185 acc0.A\[16\] _0999_/a_27_47# 0
C33186 net121 net26 0
C33187 _0554_/a_68_297# net28 0.00756f
C33188 _0626_/a_150_297# _0258_ 0
C33189 _0572_/a_373_47# net112 0
C33190 _0216_ _1026_/a_561_413# 0
C33191 _1007_/a_466_413# _0219_ 0
C33192 A[10] A[9] 0.00712f
C33193 _0174_ comp0.B\[5\] 0
C33194 _0689_/a_68_297# _0364_ 0.07822f
C33195 _0313_ _0570_/a_373_47# 0
C33196 _0648_/a_205_297# _0277_ 0
C33197 clknet_1_1__leaf__0458_ _0826_/a_301_297# 0
C33198 _0190_ _0988_/a_891_413# 0
C33199 net199 _0574_/a_109_297# 0.00211f
C33200 clkbuf_0__0459_/a_110_47# hold82/a_391_47# 0
C33201 clkbuf_1_1__f__0462_/a_110_47# _1011_/a_27_47# 0
C33202 _0217_ _1014_/a_891_413# 0.04933f
C33203 _0183_ _1014_/a_466_413# 0
C33204 _0787_/a_209_297# _0419_ 0
C33205 _1042_/a_891_413# net19 0
C33206 _0977_/a_75_212# _1069_/a_466_413# 0
C33207 _0489_ _1069_/a_27_47# 0.13831f
C33208 _1065_/a_466_413# clknet_1_0__leaf__0457_ 0
C33209 VPWR _0637_/a_56_297# 0.21984f
C33210 clkbuf_1_0__f__0458_/a_110_47# clknet_0__0458_ 0.42181f
C33211 _0131_ _0175_ 0.05686f
C33212 _0627_/a_215_53# _0369_ 0
C33213 _0984_/a_592_47# acc0.A\[15\] 0
C33214 _0195_ clkbuf_1_1__f__0457_/a_110_47# 0.01817f
C33215 net76 _0990_/a_193_47# 0.00436f
C33216 clknet_1_1__leaf__0459_ _0090_ 0.03601f
C33217 _0375_ _0237_ 0
C33218 _0130_ _0215_ 0
C33219 VPWR _1028_/a_561_413# 0.00253f
C33220 _1069_/a_634_159# _1069_/a_592_47# 0
C33221 _1056_/a_27_47# net66 0
C33222 net2 acc0.A\[11\] 0
C33223 net44 hold62/a_285_47# 0
C33224 VPWR _0723_/a_27_413# 0.24317f
C33225 net45 _0613_/a_109_297# 0
C33226 VPWR _0812_/a_510_47# 0
C33227 net204 control0.sh 0.12978f
C33228 _0320_ _0318_ 0.00246f
C33229 _0718_/a_129_47# pp[30] 0
C33230 VPWR _0514_/a_109_297# 0.19254f
C33231 clknet_0__0465_ _0990_/a_634_159# 0
C33232 _0402_ _0296_ 0.21f
C33233 _0673_/a_253_47# _0218_ 0
C33234 _1059_/a_466_413# acc0.A\[13\] 0
C33235 _1059_/a_27_47# net5 0
C33236 hold69/a_391_47# _0359_ 0
C33237 hold69/a_285_47# _0324_ 0
C33238 pp[16] hold78/a_285_47# 0
C33239 _0954_/a_220_297# comp0.B\[12\] 0.0133f
C33240 _0399_ net149 0.01437f
C33241 _0555_/a_51_297# net29 0
C33242 net203 net201 0.00235f
C33243 net84 _0347_ 0
C33244 _1041_/a_1059_315# _1040_/a_193_47# 0.00269f
C33245 _1041_/a_891_413# _1040_/a_27_47# 0.00461f
C33246 _1031_/a_891_413# _0220_ 0.04975f
C33247 net213 _0762_/a_215_47# 0.08365f
C33248 _0426_ _0291_ 0
C33249 B[8] net22 0.00159f
C33250 _0997_/a_27_47# _0411_ 0
C33251 _0398_ _1017_/a_1059_315# 0
C33252 hold55/a_49_47# net87 0
C33253 pp[10] net189 0
C33254 net48 pp[21] 0.00111f
C33255 pp[20] net49 0.00556f
C33256 hold64/a_49_47# hold64/a_285_47# 0.22264f
C33257 output66/a_27_47# net181 0.19879f
C33258 comp0.B\[2\] comp0.B\[15\] 0
C33259 _0990_/a_27_47# _0350_ 0.00512f
C33260 B[1] net24 0.0034f
C33261 B[12] hold51/a_49_47# 0.00244f
C33262 _1030_/a_891_413# net209 0
C33263 _1027_/a_193_47# _1026_/a_27_47# 0
C33264 _1027_/a_27_47# _1026_/a_193_47# 0
C33265 _0596_/a_145_75# _0183_ 0
C33266 _0244_ _0242_ 0.113f
C33267 _1018_/a_1059_315# clknet_0__0461_ 0
C33268 VPWR _0512_/a_109_47# 0
C33269 _1051_/a_1059_315# net9 0.02355f
C33270 net180 _0206_ 0
C33271 net30 comp0.B\[8\] 0
C33272 _1002_/a_891_413# _0181_ 0
C33273 hold96/a_49_47# net110 0
C33274 net139 net9 0
C33275 hold12/a_285_47# clkbuf_0_clk/a_110_47# 0.00254f
C33276 _0217_ _1022_/a_193_47# 0
C33277 acc0.A\[22\] _1022_/a_27_47# 0.00547f
C33278 clknet_1_0__leaf__0460_ clknet_1_0__leaf__0457_ 0.06421f
C33279 _0561_/a_51_297# hold84/a_49_47# 0
C33280 _0538_/a_51_297# net183 0.09172f
C33281 hold75/a_285_47# _0450_ 0.01104f
C33282 hold75/a_391_47# _0446_ 0
C33283 hold6/a_49_47# _0176_ 0.00549f
C33284 _1037_/a_1017_47# net26 0
C33285 clknet_1_1__leaf__0462_ net94 0.10825f
C33286 hold30/a_49_47# VPWR 0.29402f
C33287 comp0.B\[5\] _0208_ 0.12551f
C33288 _0474_ _0173_ 0.14618f
C33289 comp0.B\[3\] _0132_ 0.08204f
C33290 net194 _0172_ 0.01593f
C33291 hold67/a_49_47# acc0.A\[9\] 0
C33292 clknet_1_0__leaf__0463_ B[8] 0.01456f
C33293 hold20/a_285_47# _0966_/a_27_47# 0
C33294 _1022_/a_466_413# net151 0.00881f
C33295 clknet_1_1__leaf__0463_ _0565_/a_512_297# 0
C33296 hold22/a_49_47# net15 0
C33297 _0646_/a_47_47# _0218_ 0
C33298 net53 _0572_/a_27_297# 0
C33299 _1065_/a_193_47# _1062_/a_891_413# 0
C33300 clknet_1_0__leaf__0459_ _1019_/a_466_413# 0.00453f
C33301 net87 _1019_/a_193_47# 0.00178f
C33302 _0992_/a_891_413# _0421_ 0
C33303 clknet_0__0462_ _0345_ 0.04512f
C33304 clkbuf_0__0459_/a_110_47# clknet_1_1__leaf__0461_ 0
C33305 _0987_/a_27_47# acc0.A\[6\] 0
C33306 _0328_ _0686_/a_219_297# 0.01384f
C33307 net199 _1025_/a_466_413# 0
C33308 _0994_/a_193_47# _0994_/a_592_47# 0
C33309 _0994_/a_466_413# _0994_/a_561_413# 0.00772f
C33310 _0994_/a_634_159# _0994_/a_975_413# 0
C33311 _0662_/a_81_21# _0427_ 0
C33312 _0259_ _0819_/a_299_297# 0.00787f
C33313 _1020_/a_381_47# clknet_1_0__leaf__0457_ 0.01216f
C33314 _0275_ _0986_/a_1017_47# 0
C33315 hold12/a_391_47# _0460_ 0.0016f
C33316 _0357_ _0327_ 0.23074f
C33317 net211 _0772_/a_79_21# 0
C33318 _0779_/a_297_297# _0396_ 0
C33319 _0287_ _0422_ 0
C33320 _0292_ _0090_ 0.00387f
C33321 _0328_ _1008_/a_1059_315# 0
C33322 _1056_/a_27_47# _0350_ 0
C33323 _0260_ _0643_/a_103_199# 0.13341f
C33324 net6 _0184_ 0.01549f
C33325 VPWR _0739_/a_215_47# 0.00329f
C33326 _1023_/a_193_47# pp[23] 0
C33327 _1023_/a_466_413# net51 0.0124f
C33328 _0349_ net57 0
C33329 _0133_ hold84/a_49_47# 0
C33330 _0835_/a_78_199# _0256_ 0.10954f
C33331 _0855_/a_81_21# _0350_ 0.00105f
C33332 VPWR _0352_ 8.72224f
C33333 _1003_/a_381_47# net89 0.00201f
C33334 _1003_/a_891_413# _0101_ 0.05263f
C33335 clknet_0__0465_ _0433_ 0.17547f
C33336 _0954_/a_32_297# net20 0.00406f
C33337 _0954_/a_304_297# _0202_ 0
C33338 _0279_ _0789_/a_544_297# 0
C33339 _0648_/a_277_297# _0404_ 0
C33340 _0993_/a_27_47# _0993_/a_193_47# 0.97453f
C33341 _1058_/a_27_47# net192 0.02845f
C33342 _0459_ _0611_/a_150_297# 0
C33343 clknet_1_0__leaf__0459_ net219 0.25237f
C33344 _1039_/a_634_159# _1039_/a_466_413# 0.23992f
C33345 _1039_/a_193_47# _1039_/a_1059_315# 0.03384f
C33346 _1039_/a_27_47# _1039_/a_891_413# 0.02996f
C33347 _0251_ _0257_ 0
C33348 _0257_ _0640_/a_109_53# 0.03543f
C33349 hold33/a_285_47# net173 0
C33350 _1020_/a_1059_315# _0457_ 0
C33351 net46 _0757_/a_150_297# 0
C33352 _0785_/a_81_21# clkbuf_0__0465_/a_110_47# 0
C33353 net169 net15 0.21333f
C33354 _0985_/a_466_413# net170 0
C33355 _0346_ _0809_/a_384_47# 0.00124f
C33356 _0172_ _1046_/a_634_159# 0.011f
C33357 _0498_/a_512_297# clknet_1_1__leaf__0457_ 0.00225f
C33358 _1049_/a_193_47# _0196_ 0
C33359 _0684_/a_59_75# net224 0
C33360 _1026_/a_27_47# _1026_/a_1059_315# 0.04875f
C33361 _1026_/a_193_47# _1026_/a_466_413# 0.08301f
C33362 net33 _1062_/a_891_413# 0
C33363 _0733_/a_79_199# _0360_ 0.12003f
C33364 _0985_/a_634_159# clknet_1_0__leaf__0458_ 0.00511f
C33365 net203 comp0.B\[2\] 0.06748f
C33366 _1021_/a_193_47# clknet_1_0__leaf__0460_ 0.01502f
C33367 _0603_/a_68_297# _0385_ 0
C33368 net23 _1065_/a_1017_47# 0.00159f
C33369 hold59/a_285_47# _0218_ 0.00247f
C33370 net140 _1053_/a_891_413# 0.00743f
C33371 net169 _1053_/a_1059_315# 0.01047f
C33372 _0385_ hold73/a_391_47# 0.01818f
C33373 pp[9] _0515_/a_81_21# 0
C33374 clknet_0_clk _0487_ 0.06776f
C33375 _1032_/a_1059_315# clknet_1_1__leaf_clk 0.00828f
C33376 VPWR net73 0.4931f
C33377 net150 _1067_/a_1059_315# 0
C33378 _0217_ _1067_/a_466_413# 0
C33379 _0328_ acc0.A\[23\] 0
C33380 _1024_/a_466_413# _1024_/a_592_47# 0.00553f
C33381 _1024_/a_634_159# _1024_/a_1017_47# 0
C33382 net45 hold72/a_285_47# 0.0214f
C33383 net227 _0723_/a_207_413# 0
C33384 _0183_ _0383_ 0
C33385 _0426_ _0290_ 0
C33386 _0995_/a_1059_315# A[13] 0.00165f
C33387 net188 net67 0.02104f
C33388 net58 _0257_ 0
C33389 _1021_/a_1059_315# _1020_/a_466_413# 0
C33390 _1021_/a_891_413# _1020_/a_634_159# 0
C33391 clknet_1_1__leaf__0464_ _0542_/a_149_47# 0
C33392 _0195_ _0701_/a_80_21# 0
C33393 _0266_ net206 0.05184f
C33394 net48 _0352_ 0.30537f
C33395 _1036_/a_193_47# B[2] 0.00111f
C33396 net61 _0835_/a_215_47# 0.00477f
C33397 _0083_ hold71/a_49_47# 0
C33398 acc0.A\[23\] _0599_/a_113_47# 0
C33399 hold97/a_49_47# hold97/a_391_47# 0.00188f
C33400 net86 _0244_ 0
C33401 VPWR net115 0.52728f
C33402 _0574_/a_109_297# VPWR 0.19595f
C33403 hold89/a_49_47# VPWR 0.2658f
C33404 VPWR _0659_/a_150_297# 0.00155f
C33405 _0786_/a_80_21# _0992_/a_193_47# 0
C33406 _0786_/a_217_297# _0992_/a_27_47# 0
C33407 _0180_ _1049_/a_1059_315# 0.02643f
C33408 _0182_ _1049_/a_891_413# 0
C33409 _0540_/a_240_47# _0202_ 0
C33410 _0540_/a_245_297# net20 0
C33411 _0953_/a_114_297# _1040_/a_193_47# 0
C33412 _0080_ _0266_ 0
C33413 clk _1064_/a_561_413# 0
C33414 control0.add _0771_/a_215_297# 0
C33415 _1048_/a_466_413# net134 0
C33416 net53 _0360_ 0.04701f
C33417 _0402_ _0811_/a_81_21# 0.12202f
C33418 _1034_/a_1017_47# clknet_1_1__leaf__0463_ 0
C33419 _0464_ _0177_ 0
C33420 B[13] _1043_/a_27_47# 0
C33421 _0399_ _0094_ 0.02333f
C33422 VPWR _1016_/a_975_413# 0.00418f
C33423 _0731_/a_384_47# _0250_ 0.00884f
C33424 _1068_/a_634_159# _0468_ 0.03971f
C33425 _0343_ _1013_/a_634_159# 0.00173f
C33426 net1 acc0.A\[1\] 0.00428f
C33427 _1032_/a_891_413# clkbuf_1_1__f_clk/a_110_47# 0
C33428 _0234_ _0751_/a_29_53# 0.0128f
C33429 clknet_1_0__leaf__0458_ _0816_/a_68_297# 0
C33430 _0195_ _0675_/a_68_297# 0
C33431 _0415_ _0803_/a_68_297# 0.02869f
C33432 _0390_ _0352_ 0.06458f
C33433 _0748_/a_81_21# net52 0
C33434 acc0.A\[27\] _0698_/a_113_297# 0
C33435 _0340_ _0708_/a_68_297# 0.1605f
C33436 _1015_/a_193_47# comp0.B\[15\] 0
C33437 _0341_ _0708_/a_150_297# 0
C33438 _1060_/a_891_413# _0219_ 0
C33439 _0623_/a_109_297# _0255_ 0.01313f
C33440 net76 _0438_ 0
C33441 _0191_ acc0.A\[6\] 0.21298f
C33442 _0804_/a_510_47# _0404_ 0.00132f
C33443 _0223_ _0249_ 0.00125f
C33444 _0241_ _0345_ 0
C33445 net1 _0950_/a_75_212# 0.039f
C33446 _0539_/a_150_297# net21 0
C33447 clkbuf_1_0__f__0457_/a_110_47# hold73/a_285_47# 0
C33448 net32 net198 0.05244f
C33449 net152 net18 0.03682f
C33450 net167 _0974_/a_79_199# 0
C33451 _0490_ _0974_/a_222_93# 0
C33452 _0607_/a_109_297# acc0.A\[17\] 0.01696f
C33453 output58/a_27_47# acc0.A\[6\] 0.01107f
C33454 _1051_/a_466_413# _0522_/a_27_297# 0
C33455 _1051_/a_634_159# _0522_/a_109_297# 0
C33456 hold16/a_391_47# _0336_ 0.04431f
C33457 clkbuf_1_0__f__0460_/a_110_47# _1006_/a_466_413# 0.00102f
C33458 clknet_0__0460_ _1006_/a_27_47# 0
C33459 hold55/a_391_47# _0113_ 0
C33460 hold69/a_285_47# _0104_ 0
C33461 hold6/a_285_47# _0139_ 0.08305f
C33462 _1056_/a_891_413# _0189_ 0.0191f
C33463 hold26/a_391_47# _0200_ 0.00135f
C33464 _0830_/a_79_21# _0218_ 0
C33465 _0836_/a_68_297# _0186_ 0
C33466 net44 _0350_ 0
C33467 _1057_/a_27_47# _0512_/a_27_297# 0
C33468 _0622_/a_193_47# acc0.A\[8\] 0
C33469 _0294_ _0312_ 0.0034f
C33470 _1017_/a_592_47# acc0.A\[18\] 0
C33471 net44 _0111_ 0
C33472 _0249_ _1006_/a_1059_315# 0
C33473 _0250_ _1006_/a_466_413# 0
C33474 _0273_ _0827_/a_27_47# 0.05349f
C33475 _1072_/a_466_413# _1072_/a_592_47# 0.00553f
C33476 _1072_/a_634_159# _1072_/a_1017_47# 0
C33477 net212 _0186_ 0.07701f
C33478 _0343_ _0984_/a_27_47# 0.02515f
C33479 _0841_/a_79_21# _0084_ 0.0506f
C33480 _0841_/a_215_47# _0445_ 0.01154f
C33481 _0841_/a_510_47# _0444_ 0.00459f
C33482 clknet_0__0463_ _0492_/a_27_47# 0
C33483 VPWR net207 0.48008f
C33484 hold39/a_391_47# clkbuf_1_1__f__0463_/a_110_47# 0
C33485 _0251_ _0429_ 0.49451f
C33486 _0640_/a_215_297# _0640_/a_465_297# 0.00827f
C33487 _1020_/a_27_47# _0218_ 0
C33488 _1013_/a_193_47# net60 0.00442f
C33489 hold36/a_49_47# clknet_1_0__leaf__0465_ 0.007f
C33490 _0471_ _1062_/a_27_47# 0
C33491 VPWR _1025_/a_466_413# 0.24645f
C33492 _1067_/a_1059_315# control0.add 0.08524f
C33493 hold49/a_285_47# hold51/a_391_47# 0
C33494 hold49/a_391_47# hold51/a_285_47# 0
C33495 acc0.A\[27\] _0691_/a_68_297# 0
C33496 hold54/a_391_47# _0171_ 0
C33497 _0573_/a_27_47# clkbuf_1_1__f__0457_/a_110_47# 0.03805f
C33498 comp0.B\[4\] _0213_ 0
C33499 _0155_ net67 0
C33500 _0104_ _0617_/a_68_297# 0
C33501 _1041_/a_891_413# net171 0
C33502 _1041_/a_1059_315# _0207_ 0
C33503 net81 net42 0.07058f
C33504 _1012_/a_193_47# _0722_/a_215_47# 0
C33505 _1012_/a_466_413# _0722_/a_79_21# 0
C33506 _0285_ _0511_/a_299_297# 0
C33507 clknet_1_1__leaf__0459_ _0644_/a_47_47# 0.00129f
C33508 _0476_ _0559_/a_51_297# 0.01869f
C33509 net45 _0392_ 0
C33510 clknet_1_1__leaf__0460_ _1006_/a_891_413# 0.00171f
C33511 _0334_ _0333_ 1.0038f
C33512 _0473_ _1040_/a_27_47# 0
C33513 _0217_ _1024_/a_1059_315# 0
C33514 _1004_/a_561_413# _0380_ 0
C33515 _1004_/a_975_413# _0350_ 0.00116f
C33516 _0717_/a_303_47# _0348_ 0
C33517 clknet_1_0__leaf__0459_ _0352_ 0.00584f
C33518 clknet_1_0__leaf__0462_ net50 0.24121f
C33519 hold75/a_49_47# net233 0.00355f
C33520 hold75/a_391_47# net61 0
C33521 _0997_/a_466_413# _0997_/a_592_47# 0.00553f
C33522 _0997_/a_634_159# _0997_/a_1017_47# 0
C33523 _1053_/a_27_47# _0150_ 0
C33524 _0640_/a_465_297# _0465_ 0
C33525 _1037_/a_634_159# net24 0
C33526 _0583_/a_27_297# _0505_/a_27_297# 0
C33527 clknet_1_1__leaf__0459_ _0401_ 0.00199f
C33528 _0664_/a_79_21# _0346_ 0.00127f
C33529 _0371_ _0462_ 0.00724f
C33530 _0140_ _1042_/a_27_47# 0.11267f
C33531 net18 _1042_/a_466_413# 0
C33532 net198 _1042_/a_1059_315# 0.01052f
C33533 VPWR _1044_/a_27_47# 0.66574f
C33534 hold100/a_49_47# _0345_ 0.01677f
C33535 VPWR _1051_/a_1017_47# 0
C33536 _0517_/a_299_297# acc0.A\[9\] 0.00436f
C33537 _0349_ _1010_/a_1059_315# 0.0424f
C33538 net7 acc0.A\[15\] 0.00169f
C33539 _0356_ _0355_ 0
C33540 _0183_ net229 0
C33541 _0982_/a_193_47# _0345_ 0.00179f
C33542 _0783_/a_79_21# _0352_ 0.10308f
C33543 _0783_/a_510_47# _0347_ 0
C33544 VPWR _0613_/a_109_297# 0.00571f
C33545 _0756_/a_47_47# _0756_/a_377_297# 0.00899f
C33546 _1000_/a_27_47# _0216_ 0
C33547 _0151_ net13 0.08355f
C33548 net106 _0584_/a_109_297# 0
C33549 _0793_/a_149_47# _0408_ 0.00727f
C33550 _1001_/a_27_47# _0461_ 0.01374f
C33551 net243 _0378_ 0
C33552 VPWR _0551_/a_27_47# 0.25364f
C33553 _1027_/a_1059_315# _1027_/a_891_413# 0.31086f
C33554 _1027_/a_193_47# _1027_/a_975_413# 0
C33555 _1027_/a_466_413# _1027_/a_381_47# 0.03733f
C33556 _0606_/a_109_53# _0754_/a_51_297# 0
C33557 hold87/a_49_47# net234 0
C33558 _0212_ comp0.B\[4\] 0.02894f
C33559 _0253_ _0437_ 0
C33560 clknet_1_0__leaf__0463_ _0548_/a_149_47# 0
C33561 net193 hold26/a_391_47# 0.00114f
C33562 VPWR _0849_/a_79_21# 0.46137f
C33563 net10 net198 0.14895f
C33564 _0996_/a_381_47# net41 0
C33565 _0465_ _1061_/a_1017_47# 0
C33566 VPWR _1032_/a_891_413# 0.19058f
C33567 _0362_ _0776_/a_109_297# 0
C33568 _0217_ _1072_/a_1059_315# 0
C33569 clknet_1_0__leaf__0465_ _0522_/a_109_297# 0.00302f
C33570 _1061_/a_466_413# net147 0.00181f
C33571 comp0.B\[3\] net25 0.08488f
C33572 _0305_ _1009_/a_891_413# 0
C33573 net51 net241 0.00418f
C33574 _0555_/a_245_297# comp0.B\[5\] 0.00262f
C33575 _0555_/a_51_297# comp0.B\[6\] 0.00159f
C33576 clknet_0__0460_ _0737_/a_35_297# 0
C33577 _0581_/a_373_47# acc0.A\[18\] 0
C33578 hold21/a_49_47# VPWR 0.30154f
C33579 _1054_/a_592_47# A[4] 0
C33580 _0105_ _0219_ 0.02558f
C33581 _0982_/a_193_47# hold2/a_49_47# 0.00209f
C33582 _0982_/a_27_47# hold2/a_285_47# 0.00178f
C33583 B[3] B[0] 0.01301f
C33584 net64 _0622_/a_193_47# 0
C33585 _0307_ _0240_ 0
C33586 A[1] input29/a_75_212# 0
C33587 input8/a_75_212# B[6] 0
C33588 _0369_ _0307_ 0.03336f
C33589 acc0.A\[27\] _0570_/a_109_297# 0
C33590 _0571_/a_109_297# net190 0
C33591 _1035_/a_634_159# _1035_/a_592_47# 0
C33592 _0346_ _1060_/a_27_47# 0
C33593 _0410_ _0345_ 0.16273f
C33594 _0470_ _1065_/a_193_47# 0
C33595 hold76/a_49_47# clknet_1_0__leaf__0461_ 0
C33596 net17 _1064_/a_1059_315# 0
C33597 _1000_/a_193_47# _0240_ 0
C33598 _1000_/a_1059_315# _0247_ 0.07325f
C33599 net36 _0136_ 0.2835f
C33600 _0477_ comp0.B\[3\] 0
C33601 hold7/a_49_47# hold7/a_391_47# 0.00188f
C33602 _0977_/a_75_212# _0167_ 0.10895f
C33603 _0809_/a_81_21# _0809_/a_299_297# 0.08213f
C33604 net62 _0345_ 0
C33605 _0172_ _1045_/a_27_47# 0.03653f
C33606 VPWR _0533_/a_27_297# 0.22687f
C33607 _0292_ _0401_ 0.09169f
C33608 _0289_ _0290_ 0.0998f
C33609 _0287_ _0423_ 0
C33610 net33 net27 0
C33611 _0450_ _0345_ 0.03718f
C33612 _1048_/a_1059_315# acc0.A\[15\] 0
C33613 _0727_/a_277_47# acc0.A\[29\] 0
C33614 clknet_1_1__leaf__0459_ _1013_/a_27_47# 0.00122f
C33615 _1010_/a_1059_315# _0701_/a_209_297# 0
C33616 _1010_/a_891_413# _0701_/a_80_21# 0
C33617 net158 net134 0
C33618 _0718_/a_47_47# _0718_/a_129_47# 0.00369f
C33619 clkbuf_1_0__f__0465_/a_110_47# acc0.A\[6\] 0
C33620 VPWR _0546_/a_245_297# 0.006f
C33621 _1054_/a_891_413# acc0.A\[8\] 0.01471f
C33622 _0218_ _0219_ 0.27557f
C33623 acc0.A\[15\] net229 0.00555f
C33624 _0127_ _1029_/a_1059_315# 0
C33625 acc0.A\[29\] _1029_/a_561_413# 0
C33626 _0569_/a_109_297# net191 0.0033f
C33627 _1011_/a_466_413# _0726_/a_51_297# 0
C33628 hold57/a_49_47# clknet_0__0463_ 0
C33629 _1069_/a_891_413# control0.count\[0\] 0.02861f
C33630 _1033_/a_193_47# _1065_/a_193_47# 0
C33631 _1016_/a_193_47# net102 0.01325f
C33632 _1033_/a_27_47# _1065_/a_634_159# 0
C33633 _0430_ _0435_ 0.00402f
C33634 _1052_/a_634_159# _0524_/a_109_297# 0
C33635 _1052_/a_466_413# _0524_/a_27_297# 0
C33636 _0157_ acc0.A\[13\] 0
C33637 _0231_ _0223_ 0.0615f
C33638 _0343_ _0232_ 0.00221f
C33639 _0642_/a_215_297# _0826_/a_27_53# 0
C33640 _1041_/a_634_159# net174 0.00214f
C33641 _0857_/a_27_47# control0.reset 0
C33642 acc0.A\[27\] hold50/a_285_47# 0.0765f
C33643 net125 _1061_/a_466_413# 0.01867f
C33644 _0723_/a_207_413# net208 0
C33645 _0398_ _1016_/a_27_47# 0
C33646 _0488_ _0485_ 0
C33647 _0466_ _0484_ 0
C33648 _0985_/a_27_47# _0195_ 0
C33649 hold64/a_391_47# _0183_ 0.01621f
C33650 _0577_/a_109_297# _0183_ 0.00759f
C33651 VPWR net106 0.38236f
C33652 _0251_ clknet_1_1__leaf__0458_ 0.00242f
C33653 _0640_/a_109_53# clknet_1_1__leaf__0458_ 0
C33654 _0182_ _0171_ 0.00134f
C33655 _0750_/a_181_47# _0219_ 0
C33656 _0461_ _0459_ 0.00696f
C33657 _0467_ _1067_/a_27_47# 0
C33658 hold20/a_285_47# clkload0/a_27_47# 0
C33659 _0470_ net33 0.21557f
C33660 hold15/a_285_47# hold15/a_391_47# 0.41909f
C33661 net243 acc0.A\[24\] 0
C33662 _0311_ _0310_ 0.00373f
C33663 _0663_/a_27_413# VPWR 0.19567f
C33664 comp0.B\[2\] _0176_ 0
C33665 _0426_ net77 0
C33666 _0563_/a_51_297# _0173_ 0.08441f
C33667 _0208_ hold84/a_49_47# 0
C33668 _0201_ _0143_ 0
C33669 hold58/a_49_47# _1034_/a_27_47# 0
C33670 _0227_ _0345_ 0.02031f
C33671 _0328_ clknet_1_1__leaf__0462_ 0
C33672 VPWR _0237_ 0.7341f
C33673 clknet_1_0__leaf__0463_ net247 0.00561f
C33674 _0524_/a_27_297# _0194_ 0.12192f
C33675 _0673_/a_253_47# net228 0.00478f
C33676 pp[25] _0216_ 0
C33677 net53 _0124_ 0.00537f
C33678 _1065_/a_466_413# _0160_ 0
C33679 hold75/a_285_47# _0637_/a_56_297# 0
C33680 clknet_1_0__leaf__0459_ net207 0.03891f
C33681 net104 _0264_ 0
C33682 _0475_ _0563_/a_149_47# 0.004f
C33683 _0995_/a_193_47# output41/a_27_47# 0
C33684 net211 _1019_/a_27_47# 0.00901f
C33685 _0217_ _0580_/a_27_297# 0.09314f
C33686 _0404_ _0798_/a_113_297# 0.07539f
C33687 _0800_/a_51_297# _0400_ 0
C33688 hold50/a_285_47# _0364_ 0
C33689 _0982_/a_1059_315# net36 0.12351f
C33690 _0520_/a_27_297# _0520_/a_373_47# 0.01338f
C33691 VPWR hold72/a_285_47# 0.29769f
C33692 _1067_/a_27_47# comp0.B\[0\] 0
C33693 hold24/a_391_47# clknet_1_0__leaf__0463_ 0
C33694 net45 _1013_/a_1059_315# 0.02187f
C33695 _1018_/a_193_47# _0247_ 0.00246f
C33696 _0780_/a_285_297# _0240_ 0
C33697 _0179_ _1048_/a_1059_315# 0
C33698 _0238_ _0617_/a_150_297# 0
C33699 _0361_ acc0.A\[27\] 0.00228f
C33700 net58 clknet_1_1__leaf__0458_ 0.31664f
C33701 net177 net51 0.13393f
C33702 _1043_/a_27_47# _1042_/a_634_159# 0.00117f
C33703 _1043_/a_193_47# _1042_/a_193_47# 0
C33704 _1043_/a_634_159# _1042_/a_27_47# 0.00117f
C33705 _0858_/a_27_47# net71 0
C33706 _0181_ _1048_/a_27_47# 0
C33707 _0777_/a_129_47# _0347_ 0
C33708 _1055_/a_193_47# net74 0
C33709 _0803_/a_68_297# _0347_ 0
C33710 net236 _0484_ 0.13366f
C33711 hold7/a_49_47# clknet_1_1__leaf__0458_ 0.04975f
C33712 _0375_ _0222_ 0.61273f
C33713 _0179_ net229 0.19925f
C33714 _0769_/a_299_297# VPWR 0.19529f
C33715 clknet_0__0458_ acc0.A\[15\] 0.0049f
C33716 _1019_/a_891_413# _0399_ 0
C33717 A[12] net2 0
C33718 _0993_/a_466_413# _0993_/a_592_47# 0.00553f
C33719 _0993_/a_634_159# _0993_/a_1017_47# 0
C33720 _0426_ _0656_/a_59_75# 0
C33721 hold33/a_49_47# _0142_ 0
C33722 hold87/a_285_47# VPWR 0.29391f
C33723 _0437_ output61/a_27_47# 0
C33724 _1039_/a_466_413# net125 0
C33725 _0180_ net175 0.05424f
C33726 _0199_ _0531_/a_373_47# 0
C33727 _0134_ clknet_0__0463_ 0
C33728 VPWR _0529_/a_27_297# 0.21861f
C33729 _0280_ _0304_ 0.00143f
C33730 net175 net218 0
C33731 _1038_/a_891_413# _0463_ 0
C33732 _0973_/a_109_47# clknet_1_0__leaf__0460_ 0.00152f
C33733 _0673_/a_337_297# _0347_ 0.00284f
C33734 _0146_ _0530_/a_81_21# 0
C33735 _0343_ _0707_/a_75_199# 0.00601f
C33736 _0083_ net170 0
C33737 hold20/a_285_47# _0981_/a_27_297# 0
C33738 _0209_ clkbuf_1_0__f__0463_/a_110_47# 0.00101f
C33739 _0724_/a_113_297# _0333_ 0.0494f
C33740 _0172_ net132 0
C33741 _0159_ clknet_1_1__leaf__0457_ 0.08647f
C33742 _0714_/a_51_297# _1031_/a_27_47# 0
C33743 net48 _0237_ 0.41941f
C33744 _0399_ net206 0.0283f
C33745 comp0.B\[7\] clknet_0__0463_ 0
C33746 _0485_ _1064_/a_27_47# 0.00222f
C33747 net73 _0523_/a_81_21# 0.00115f
C33748 _0549_/a_68_297# _0173_ 0.00192f
C33749 clknet_1_1__leaf__0463_ _0564_/a_150_297# 0.00125f
C33750 _0624_/a_59_75# clkbuf_1_0__f__0465_/a_110_47# 0
C33751 _1026_/a_634_159# net112 0
C33752 _1026_/a_891_413# _1026_/a_1017_47# 0.00617f
C33753 _1059_/a_466_413# VPWR 0.25261f
C33754 net107 hold93/a_391_47# 0
C33755 _0985_/a_1059_315# _0449_ 0
C33756 _0465_ _1047_/a_193_47# 0.01037f
C33757 _0133_ control0.reset 0
C33758 _0480_ _0975_/a_59_75# 0
C33759 _0234_ net91 0
C33760 _0999_/a_193_47# _0779_/a_79_21# 0
C33761 _1072_/a_27_47# control0.state\[2\] 0
C33762 _0172_ hold5/a_391_47# 0.00171f
C33763 _0472_ _1061_/a_193_47# 0
C33764 _0195_ _0330_ 0.02873f
C33765 _0697_/a_300_47# _0324_ 0.0019f
C33766 _0080_ _0399_ 0
C33767 _0817_/a_81_21# _0817_/a_266_297# 0.01575f
C33768 net58 _0263_ 0.0657f
C33769 _0718_/a_285_47# _0348_ 0.06696f
C33770 _0181_ _1009_/a_891_413# 0.00106f
C33771 _0156_ _0186_ 0
C33772 _0347_ acc0.A\[18\] 0.0472f
C33773 A[5] _0150_ 0
C33774 _1024_/a_592_47# _0122_ 0
C33775 _1024_/a_381_47# acc0.A\[24\] 0
C33776 _0455_ _1018_/a_193_47# 0
C33777 _0346_ _0586_/a_27_47# 0.01367f
C33778 hold30/a_391_47# net50 0
C33779 hold9/a_391_47# _0345_ 0
C33780 _0670_/a_79_21# acc0.A\[13\] 0
C33781 hold47/a_49_47# _0527_/a_27_297# 0.0441f
C33782 _0230_ _0754_/a_512_297# 0
C33783 net168 net11 0.47373f
C33784 _0642_/a_215_297# _0087_ 0
C33785 _0376_ _0232_ 0
C33786 clknet_1_1__leaf__0459_ hold70/a_49_47# 0.01043f
C33787 hold99/a_49_47# pp[11] 0.00284f
C33788 _0429_ net168 0.00345f
C33789 hold36/a_391_47# net131 0
C33790 hold36/a_285_47# net184 0
C33791 _0174_ _1040_/a_634_159# 0.01246f
C33792 net34 _0978_/a_27_297# 0
C33793 _1037_/a_634_159# _1037_/a_466_413# 0.23992f
C33794 _1037_/a_193_47# _1037_/a_1059_315# 0.03112f
C33795 _1037_/a_27_47# _1037_/a_891_413# 0.03224f
C33796 hold53/a_49_47# net52 0
C33797 acc0.A\[22\] _0756_/a_285_47# 0
C33798 _0767_/a_59_75# _0462_ 0
C33799 comp0.B\[10\] _1040_/a_1059_315# 0.06421f
C33800 _0369_ _0507_/a_109_297# 0.00576f
C33801 _0186_ _0989_/a_891_413# 0
C33802 _0835_/a_78_199# clknet_0__0465_ 0
C33803 _0473_ net24 0.02336f
C33804 _0785_/a_299_297# _0401_ 0.0135f
C33805 clknet_1_1__leaf_clk _0468_ 0.06288f
C33806 clknet_0__0458_ _0179_ 0.1209f
C33807 _0195_ _0242_ 0
C33808 _0216_ acc0.A\[19\] 0.17608f
C33809 acc0.A\[1\] control0.sh 0.01034f
C33810 _0242_ net92 0.00391f
C33811 VPWR _1005_/a_27_47# 0.73106f
C33812 _0790_/a_35_297# net42 0.22438f
C33813 _0369_ hold82/a_49_47# 0.01443f
C33814 _1041_/a_634_159# _1041_/a_592_47# 0
C33815 VPWR _0991_/a_561_413# 0.00314f
C33816 _0504_/a_27_47# _0182_ 0.2159f
C33817 _1054_/a_634_159# _0180_ 0.02168f
C33818 hold30/a_49_47# _1023_/a_27_47# 0
C33819 _0555_/a_51_297# net26 0.00166f
C33820 _0390_ _0769_/a_299_297# 0
C33821 VPWR _0392_ 0.95171f
C33822 _0243_ hold87/a_391_47# 0
C33823 _1002_/a_975_413# net1 0.00163f
C33824 VPWR _0600_/a_253_297# 0.00196f
C33825 _1057_/a_193_47# net2 0
C33826 _1038_/a_27_47# net8 0
C33827 _0176_ _1043_/a_891_413# 0
C33828 _0337_ hold15/a_285_47# 0
C33829 _1057_/a_891_413# A[11] 0
C33830 _1039_/a_466_413# _0473_ 0.0129f
C33831 _1039_/a_193_47# _0472_ 0.02507f
C33832 hold9/a_49_47# _1008_/a_27_47# 0
C33833 _0625_/a_59_75# _0989_/a_193_47# 0
C33834 _0469_ clkbuf_1_1__f_clk/a_110_47# 0
C33835 _0366_ net112 0
C33836 _0149_ _0522_/a_27_297# 0.00107f
C33837 hold86/a_391_47# _0219_ 0.06065f
C33838 acc0.A\[29\] hold62/a_391_47# 0
C33839 _0366_ acc0.A\[24\] 0.4057f
C33840 clkbuf_0__0459_/a_110_47# clknet_1_1__leaf__0465_ 0
C33841 clknet_1_1__leaf__0460_ _0679_/a_68_297# 0
C33842 _0216_ _0249_ 0
C33843 VPWR _1011_/a_466_413# 0.2435f
C33844 _0195_ _0197_ 0.17961f
C33845 hold59/a_49_47# _0347_ 0.00201f
C33846 _0234_ _0762_/a_510_47# 0.00111f
C33847 _0752_/a_27_413# _0383_ 0.00305f
C33848 _0479_ _0468_ 0
C33849 _1055_/a_27_47# net62 0
C33850 _1029_/a_27_47# _1008_/a_27_47# 0.00214f
C33851 _0300_ net41 0.00196f
C33852 _0963_/a_35_297# _1069_/a_1059_315# 0
C33853 hold65/a_391_47# net248 0
C33854 _0195_ _1030_/a_27_47# 0.03524f
C33855 _1030_/a_193_47# net57 0
C33856 _0465_ _0265_ 0.00953f
C33857 _0252_ _0253_ 0.22825f
C33858 _0226_ _0228_ 0.03482f
C33859 _0640_/a_465_297# _0254_ 0.00112f
C33860 net48 _1005_/a_27_47# 0.01536f
C33861 _0369_ net4 0
C33862 _0108_ clknet_1_1__leaf__0462_ 0
C33863 net215 _0102_ 0
C33864 A[10] _0515_/a_299_297# 0.0054f
C33865 _0292_ _0089_ 0
C33866 _0891_/a_27_47# _1033_/a_27_47# 0
C33867 _1019_/a_466_413# _0345_ 0.03311f
C33868 _0361_ _1009_/a_634_159# 0
C33869 _0467_ net186 0
C33870 output67/a_27_47# _1058_/a_193_47# 0
C33871 _0985_/a_193_47# _0846_/a_512_297# 0
C33872 _0764_/a_81_21# hold73/a_49_47# 0
C33873 net247 net165 0.00594f
C33874 net67 hold81/a_49_47# 0
C33875 acc0.A\[1\] net157 0.02778f
C33876 clknet_1_0__leaf__0459_ hold72/a_285_47# 0.01812f
C33877 _1012_/a_1059_315# _0110_ 0
C33878 _0369_ clkbuf_1_0__f__0460_/a_110_47# 0.00705f
C33879 clknet_0__0457_ net118 0
C33880 _0412_ pp[14] 0
C33881 acc0.A\[22\] _0122_ 0
C33882 _0183_ net110 0
C33883 hold33/a_49_47# clknet_0__0463_ 0
C33884 _0272_ _0445_ 0
C33885 net213 net150 0
C33886 _0218_ _0799_/a_209_297# 0.00865f
C33887 _0195_ net190 0.3014f
C33888 _0216_ net197 0.3138f
C33889 _0578_/a_373_47# VPWR 0
C33890 _0147_ net10 0
C33891 _0487_ _1065_/a_27_47# 0
C33892 _0369_ _0250_ 0.30231f
C33893 net69 _0350_ 0.00386f
C33894 _0579_/a_373_47# _0352_ 0
C33895 net158 net22 0
C33896 _0359_ _0219_ 0.33655f
C33897 _0146_ _1049_/a_466_413# 0.00218f
C33898 clknet_1_0__leaf__0464_ net11 0
C33899 net186 comp0.B\[0\] 0
C33900 _0225_ _0223_ 0.12491f
C33901 net95 _1009_/a_27_47# 0.22685f
C33902 net12 _0142_ 0
C33903 _0154_ net2 0
C33904 net101 clkbuf_0__0457_/a_110_47# 0.00221f
C33905 _0262_ _0263_ 0.10421f
C33906 _0289_ _0656_/a_59_75# 0
C33907 _1003_/a_27_47# acc0.A\[21\] 0
C33908 _0756_/a_285_47# _0379_ 0.04387f
C33909 net86 _0195_ 0
C33910 _0495_/a_68_297# _0171_ 0.07338f
C33911 _0461_ _0772_/a_79_21# 0.00384f
C33912 _1035_/a_1059_315# _0561_/a_240_47# 0
C33913 _1035_/a_27_47# _0173_ 0
C33914 clkbuf_1_1__f__0465_/a_110_47# _0090_ 0.00141f
C33915 _0606_/a_109_53# _0219_ 0.00555f
C33916 _1027_/a_381_47# net156 0.12224f
C33917 net178 _0179_ 0.11892f
C33918 _0643_/a_253_47# _0272_ 0.03027f
C33919 _0643_/a_253_297# _0275_ 0.00228f
C33920 _0643_/a_337_297# _0274_ 0.00121f
C33921 pp[17] _0340_ 0.03072f
C33922 _0985_/a_27_47# clkbuf_1_0__f__0458_/a_110_47# 0
C33923 comp0.B\[8\] _1040_/a_27_47# 0.08236f
C33924 VPWR _0196_ 0.38039f
C33925 net168 clknet_1_1__leaf__0458_ 0
C33926 hold76/a_49_47# _0218_ 0
C33927 hold97/a_285_47# _0698_/a_113_297# 0.00163f
C33928 net158 clknet_1_0__leaf__0463_ 0.01078f
C33929 _1059_/a_466_413# clknet_1_0__leaf__0459_ 0
C33930 _0697_/a_80_21# _0352_ 0
C33931 _0957_/a_32_297# _0957_/a_220_297# 0.00132f
C33932 _0749_/a_384_47# _0248_ 0.00921f
C33933 _0749_/a_299_297# _0372_ 0.05215f
C33934 net56 _0352_ 0
C33935 clknet_1_0__leaf__0462_ _1023_/a_592_47# 0
C33936 VPWR net122 0.4261f
C33937 control0.sh _0562_/a_68_297# 0
C33938 _0346_ net149 0.02468f
C33939 _0855_/a_81_21# _1014_/a_27_47# 0
C33940 hold23/a_49_47# net71 0
C33941 _0478_ _1071_/a_1059_315# 0
C33942 _1007_/a_27_47# _1007_/a_1059_315# 0.04875f
C33943 _1007_/a_193_47# _1007_/a_466_413# 0.0751f
C33944 _1052_/a_634_159# _1052_/a_1059_315# 0
C33945 _1052_/a_27_47# _1052_/a_381_47# 0.05761f
C33946 _1052_/a_193_47# _1052_/a_891_413# 0.19489f
C33947 net202 _1015_/a_891_413# 0
C33948 acc0.A\[20\] _0460_ 0.06303f
C33949 _0991_/a_1017_47# clknet_1_1__leaf__0465_ 0
C33950 _1035_/a_975_413# _0133_ 0
C33951 _1035_/a_592_47# net121 0
C33952 _0469_ VPWR 0.23425f
C33953 hold87/a_285_47# _0453_ 0.00197f
C33954 net33 _0485_ 0
C33955 net186 _1034_/a_634_159# 0.00122f
C33956 net121 B[15] 0
C33957 _0330_ _1010_/a_891_413# 0
C33958 _0108_ net242 0
C33959 _0973_/a_27_297# hold93/a_285_47# 0.00119f
C33960 _1058_/a_634_159# _1058_/a_381_47# 0
C33961 net139 A[7] 0.02618f
C33962 _0570_/a_27_297# _1027_/a_27_47# 0.00955f
C33963 hold14/a_391_47# net24 0
C33964 control0.state\[1\] _0480_ 0
C33965 _1051_/a_592_47# _0172_ 0.00248f
C33966 _0312_ _0371_ 0.11291f
C33967 _0404_ net41 0
C33968 _0399_ _0405_ 0.04048f
C33969 VPWR _0199_ 0.23106f
C33970 _0585_/a_109_297# _0465_ 0
C33971 _0680_/a_217_297# _0305_ 0.02394f
C33972 hold12/a_285_47# _0487_ 0.03317f
C33973 acc0.A\[12\] _0510_/a_27_297# 0.13821f
C33974 _0261_ _0509_/a_27_47# 0
C33975 _0252_ net74 0.00515f
C33976 acc0.A\[20\] _0457_ 0
C33977 clkbuf_0_clk/a_110_47# clknet_1_0__leaf_clk 0.0021f
C33978 _1011_/a_381_47# _0354_ 0.01345f
C33979 _1011_/a_891_413# _0355_ 0.02219f
C33980 _1011_/a_1059_315# net227 0.00496f
C33981 _1011_/a_193_47# _0109_ 0.41262f
C33982 VPWR _1013_/a_1059_315# 0.39929f
C33983 clknet_0__0465_ _0516_/a_27_297# 0
C33984 _0243_ _0264_ 0.00133f
C33985 clknet_1_0__leaf__0465_ _0150_ 0.00764f
C33986 net119 _1065_/a_27_47# 0
C33987 _1002_/a_634_159# VPWR 0.18117f
C33988 clkbuf_1_1__f__0457_/a_110_47# acc0.A\[15\] 0
C33989 _0174_ control0.reset 0
C33990 _0949_/a_59_75# clknet_0_clk 0.01537f
C33991 _0781_/a_68_297# clkbuf_1_1__f__0461_/a_110_47# 0.00133f
C33992 _1052_/a_466_413# _0194_ 0
C33993 _0983_/a_193_47# _0854_/a_79_21# 0
C33994 clknet_1_0__leaf__0459_ _0392_ 0
C33995 _0538_/a_245_297# comp0.B\[14\] 0.0012f
C33996 clkload4/a_110_47# hold19/a_49_47# 0
C33997 _0831_/a_285_297# clknet_1_1__leaf__0458_ 0.00337f
C33998 _0812_/a_510_47# _0345_ 0
C33999 _0362_ _0318_ 0.06179f
C34000 acc0.A\[9\] _0990_/a_1059_315# 0.01122f
C34001 _1027_/a_381_47# acc0.A\[26\] 0.00137f
C34002 _0252_ output61/a_27_47# 0
C34003 net58 _0988_/a_1017_47# 0
C34004 hold13/a_285_47# net24 0
C34005 _0277_ _0400_ 0
C34006 _1038_/a_561_413# _0176_ 0
C34007 _0231_ _0216_ 0.00919f
C34008 net23 clknet_1_0__leaf__0461_ 0.81055f
C34009 hold70/a_285_47# _0281_ 0
C34010 net228 _0219_ 0
C34011 pp[18] _0341_ 0.00687f
C34012 _0974_/a_79_199# _0974_/a_448_47# 0.04614f
C34013 _0197_ _1048_/a_193_47# 0
C34014 net205 _1034_/a_1059_315# 0
C34015 _0257_ _0625_/a_145_75# 0.00152f
C34016 net106 _0113_ 0
C34017 hold11/a_391_47# _1049_/a_27_47# 0
C34018 net47 _0261_ 0
C34019 _0984_/a_634_159# VPWR 0.18036f
C34020 _0880_/a_27_47# _0460_ 0.11344f
C34021 _0172_ _0546_/a_51_297# 0.20526f
C34022 _0746_/a_81_21# _0359_ 0.05746f
C34023 _0994_/a_1059_315# _0218_ 0.003f
C34024 _0216_ net1 0.02786f
C34025 net59 _1012_/a_561_413# 0
C34026 _0267_ _0465_ 0.01189f
C34027 acc0.A\[12\] _0181_ 0.1088f
C34028 net61 _0836_/a_150_297# 0
C34029 _0414_ net80 0.01223f
C34030 net78 _0399_ 0
C34031 _0399_ clknet_0__0465_ 0.09921f
C34032 net111 _1026_/a_634_159# 0
C34033 _0217_ _0117_ 0
C34034 _0520_/a_109_47# _0186_ 0.00438f
C34035 _0201_ _0174_ 0.11535f
C34036 _0776_/a_109_297# _0347_ 0
C34037 clkbuf_1_0__f__0462_/a_110_47# _1007_/a_27_47# 0.01244f
C34038 _1002_/a_634_159# net48 0
C34039 VPWR _1042_/a_381_47# 0.0711f
C34040 _0251_ _0642_/a_27_413# 0.26689f
C34041 net61 _0437_ 0.04555f
C34042 _0982_/a_466_413# _0346_ 0.02079f
C34043 _0343_ _0795_/a_81_21# 0.0026f
C34044 net35 done 0.00955f
C34045 _0544_/a_51_297# _0202_ 0
C34046 _0195_ _0855_/a_81_21# 0.00446f
C34047 net55 _0219_ 0.05118f
C34048 net183 comp0.B\[10\] 0
C34049 pp[26] _0572_/a_109_47# 0
C34050 output54/a_27_47# _0195_ 0
C34051 _1043_/a_27_47# net128 0
C34052 VPWR _0763_/a_193_47# 0
C34053 _0998_/a_1059_315# net83 0
C34054 clknet_0__0460_ _1009_/a_1059_315# 0
C34055 _1030_/a_466_413# acc0.A\[30\] 0.02579f
C34056 _0642_/a_382_47# _0252_ 0
C34057 _0682_/a_150_297# _0366_ 0
C34058 _0682_/a_68_297# _0315_ 0
C34059 hold89/a_391_47# _0466_ 0.07918f
C34060 _0273_ _0989_/a_193_47# 0.00208f
C34061 _0179_ clkbuf_1_1__f__0457_/a_110_47# 0
C34062 _0500_/a_27_47# clknet_1_1__leaf__0457_ 0.06471f
C34063 _0988_/a_193_47# _0988_/a_381_47# 0.09642f
C34064 _0988_/a_634_159# _0988_/a_891_413# 0.03684f
C34065 _0988_/a_27_47# _0988_/a_561_413# 0.0027f
C34066 hold3/a_285_47# _0219_ 0.00237f
C34067 control0.reset _0208_ 0.02813f
C34068 _0352_ _0345_ 0.30296f
C34069 _0313_ clkbuf_0__0462_/a_110_47# 0
C34070 _1039_/a_27_47# _0136_ 0
C34071 _1039_/a_891_413# _0174_ 0.0011f
C34072 net49 net109 0
C34073 VPWR _0560_/a_150_297# 0.002f
C34074 _0368_ _0367_ 0.11064f
C34075 _0278_ _0301_ 0
C34076 net1 _1067_/a_27_47# 0
C34077 _0730_/a_297_297# _0108_ 0.00157f
C34078 _0730_/a_510_47# _0358_ 0.00286f
C34079 _0699_/a_150_297# _0350_ 0
C34080 hold64/a_285_47# acc0.A\[19\] 0.09248f
C34081 _0343_ _0338_ 0.00117f
C34082 hold20/a_285_47# _0170_ 0
C34083 _0255_ acc0.A\[8\] 0.00144f
C34084 _0629_/a_59_75# hold100/a_391_47# 0.01341f
C34085 _0678_/a_68_297# _0780_/a_35_297# 0.01292f
C34086 _0542_/a_149_47# _0542_/a_240_47# 0.06872f
C34087 _0542_/a_51_297# _0203_ 0.11476f
C34088 _0822_/a_109_297# _0399_ 0
C34089 net225 _1031_/a_27_47# 0
C34090 net63 _0087_ 0.10854f
C34091 _0162_ _1064_/a_975_413# 0
C34092 _0857_/a_27_47# _0457_ 0.11023f
C34093 _1026_/a_592_47# acc0.A\[26\] 0
C34094 _0157_ VPWR 0.37155f
C34095 _0982_/a_466_413# _0629_/a_59_75# 0
C34096 _0179_ input15/a_75_212# 0
C34097 _1001_/a_466_413# clknet_1_0__leaf__0457_ 0.00279f
C34098 _0999_/a_634_159# _0097_ 0.00105f
C34099 _0460_ _1062_/a_27_47# 0.00135f
C34100 net112 acc0.A\[24\] 0
C34101 _0817_/a_585_47# _0424_ 0
C34102 clknet_1_1__leaf__0460_ _1009_/a_592_47# 0
C34103 _0222_ VPWR 1.06149f
C34104 _0118_ net223 0
C34105 _1035_/a_466_413# net27 0
C34106 _1021_/a_27_47# clknet_1_0__leaf__0457_ 0.01442f
C34107 net87 net202 0
C34108 net19 net20 0.04452f
C34109 _0141_ _0202_ 0.02746f
C34110 _0454_ net104 0
C34111 _0251_ _0218_ 0
C34112 hold48/a_391_47# net195 0.13067f
C34113 _0640_/a_109_53# _0218_ 0
C34114 hold36/a_285_47# net130 0
C34115 _1038_/a_891_413# clkbuf_1_0__f__0463_/a_110_47# 0
C34116 net236 hold89/a_391_47# 0.13866f
C34117 net40 pp[13] 0.01375f
C34118 _0279_ _0994_/a_634_159# 0
C34119 _0278_ _0994_/a_193_47# 0
C34120 _0299_ _0405_ 0
C34121 _0792_/a_80_21# _0219_ 0.0635f
C34122 _0363_ _0370_ 0.00197f
C34123 _0305_ _0372_ 0
C34124 _0347_ _1008_/a_193_47# 0.02993f
C34125 _0228_ _0760_/a_47_47# 0
C34126 _1037_/a_634_159# _0135_ 0.04448f
C34127 net111 _0366_ 0
C34128 _0531_/a_27_297# _1048_/a_27_47# 0.01072f
C34129 _0997_/a_891_413# _0218_ 0.00558f
C34130 hold38/a_285_47# clkbuf_1_1__f__0463_/a_110_47# 0
C34131 _0195_ _0998_/a_381_47# 0.01241f
C34132 _0604_/a_113_47# control0.add 0
C34133 output67/a_27_47# pp[9] 0.37481f
C34134 clknet_1_0__leaf__0462_ _0576_/a_27_297# 0.02102f
C34135 net231 _0951_/a_368_53# 0
C34136 pp[30] _1030_/a_891_413# 0.0131f
C34137 _0779_/a_215_47# clknet_1_1__leaf__0461_ 0
C34138 net115 _0345_ 0.03522f
C34139 _0635_/a_109_297# _0635_/a_27_47# 0
C34140 net36 clknet_1_0__leaf__0465_ 0
C34141 _0285_ _0786_/a_217_297# 0
C34142 net58 _0848_/a_27_47# 0
C34143 net171 comp0.B\[8\] 0
C34144 _1039_/a_891_413# _0208_ 0
C34145 hold24/a_49_47# _0209_ 0.01405f
C34146 _0985_/a_634_159# _0448_ 0
C34147 _0985_/a_891_413# _0447_ 0
C34148 _0959_/a_217_297# net23 0
C34149 net140 _0180_ 0.01575f
C34150 net58 _0218_ 0.65408f
C34151 pp[12] _0994_/a_891_413# 0.00271f
C34152 _1001_/a_27_47# _1001_/a_561_413# 0.0027f
C34153 _1001_/a_634_159# _1001_/a_891_413# 0.03684f
C34154 _1001_/a_193_47# _1001_/a_381_47# 0.09503f
C34155 _0705_/a_59_75# hold80/a_391_47# 0
C34156 _0442_ net148 0
C34157 net48 _0222_ 0.0328f
C34158 _1062_/a_634_159# _1062_/a_466_413# 0.23992f
C34159 _1062_/a_193_47# _1062_/a_1059_315# 0.03405f
C34160 _1062_/a_27_47# _1062_/a_891_413# 0.03224f
C34161 VPWR net220 0.2141f
C34162 _0239_ _0677_/a_285_47# 0
C34163 _1020_/a_193_47# _1032_/a_27_47# 0
C34164 _1020_/a_27_47# _1032_/a_193_47# 0
C34165 net81 net5 0
C34166 _0341_ _0567_/a_109_47# 0
C34167 _0340_ _0567_/a_109_297# 0
C34168 clknet_1_0__leaf__0458_ _0266_ 0.01981f
C34169 _1011_/a_193_47# _0725_/a_80_21# 0
C34170 _1011_/a_27_47# _0725_/a_209_297# 0.00119f
C34171 _0183_ _0486_ 0
C34172 _0473_ _0953_/a_304_297# 0
C34173 _0461_ _0178_ 0.00113f
C34174 _1021_/a_27_47# _1021_/a_193_47# 0.96682f
C34175 _0149_ _0193_ 0
C34176 _0343_ net99 0
C34177 hold90/a_285_47# hold90/a_391_47# 0.41909f
C34178 _1003_/a_193_47# net49 0.00432f
C34179 net61 _0626_/a_68_297# 0.01809f
C34180 net44 _0195_ 0.24879f
C34181 _0575_/a_27_297# _1024_/a_466_413# 0
C34182 hold41/a_49_47# hold41/a_285_47# 0.22264f
C34183 clkbuf_1_1__f__0465_/a_110_47# _0401_ 0
C34184 _0419_ _0807_/a_68_297# 0.10661f
C34185 net64 _0255_ 0
C34186 net235 _0434_ 0
C34187 _1049_/a_1059_315# _1048_/a_891_413# 0
C34188 _1049_/a_466_413# _1048_/a_381_47# 0
C34189 _0227_ hold94/a_391_47# 0.05913f
C34190 _0758_/a_510_47# acc0.A\[23\] 0.00213f
C34191 VPWR _1006_/a_592_47# 0
C34192 _0248_ hold73/a_285_47# 0
C34193 VPWR acc0.A\[9\] 1.34799f
C34194 _0284_ _0787_/a_209_297# 0.00707f
C34195 _1000_/a_634_159# _0183_ 0
C34196 hold43/a_391_47# _1029_/a_193_47# 0
C34197 hold43/a_49_47# _1029_/a_466_413# 0
C34198 _0963_/a_117_297# _0167_ 0
C34199 _0963_/a_285_297# clknet_1_0__leaf_clk 0.05102f
C34200 hold47/a_49_47# _0143_ 0
C34201 hold4/a_49_47# net51 0.01088f
C34202 net78 _0295_ 0
C34203 clknet_1_1__leaf__0464_ _1043_/a_193_47# 0.46397f
C34204 net207 _0345_ 0.00335f
C34205 _0083_ _0846_/a_51_297# 0.1022f
C34206 _0742_/a_299_297# _0368_ 0.00661f
C34207 _0325_ _0219_ 0.02171f
C34208 VPWR _0670_/a_79_21# 0.49229f
C34209 _0280_ _0992_/a_1059_315# 0
C34210 _1020_/a_27_47# _0721_/a_27_47# 0.0026f
C34211 _0092_ _0994_/a_27_47# 0.10191f
C34212 _0388_ _0462_ 0.00126f
C34213 _0186_ _0988_/a_1059_315# 0
C34214 _0371_ _0746_/a_299_297# 0
C34215 _1004_/a_381_47# _0216_ 0.00487f
C34216 _0460_ net107 0.00661f
C34217 _0224_ _1022_/a_193_47# 0
C34218 net225 _0712_/a_79_21# 0
C34219 _0361_ _0366_ 0
C34220 _0561_/a_245_297# _0561_/a_240_47# 0
C34221 _0221_ _0723_/a_207_413# 0.00245f
C34222 net48 net220 0.13298f
C34223 _1072_/a_634_159# _1068_/a_891_413# 0
C34224 _1072_/a_466_413# _1068_/a_1059_315# 0
C34225 _0476_ _1065_/a_466_413# 0
C34226 VPWR _0762_/a_297_297# 0.01069f
C34227 _0251_ _0833_/a_215_47# 0
C34228 _0230_ acc0.A\[23\] 0.00429f
C34229 _0662_/a_384_47# _0294_ 0.00137f
C34230 _0146_ _0147_ 0
C34231 _0404_ net80 0
C34232 hold41/a_391_47# _0179_ 0.05619f
C34233 _0346_ _0256_ 0
C34234 net82 _0459_ 0.00257f
C34235 hold30/a_285_47# clknet_1_0__leaf__0460_ 0.00178f
C34236 pp[0] A[1] 0.15395f
C34237 _0352_ net52 0.67516f
C34238 acc0.A\[27\] VPWR 1.8034f
C34239 comp0.B\[13\] _0201_ 0.32683f
C34240 _1036_/a_27_47# net122 0.23091f
C34241 _1036_/a_634_159# clknet_1_1__leaf__0463_ 0.01399f
C34242 _0346_ _0987_/a_1059_315# 0.00111f
C34243 net71 hold71/a_49_47# 0
C34244 VPWR _0707_/a_544_297# 0.00635f
C34245 _0461_ _1019_/a_27_47# 0.042f
C34246 _0538_/a_149_47# _1046_/a_891_413# 0
C34247 _0238_ _0219_ 0.00447f
C34248 _1041_/a_27_47# net153 0.09539f
C34249 _1041_/a_193_47# net127 0.00655f
C34250 _1047_/a_1059_315# _1047_/a_891_413# 0.31086f
C34251 _1047_/a_193_47# _1047_/a_975_413# 0
C34252 _1047_/a_466_413# _1047_/a_381_47# 0.03733f
C34253 net1 net100 0
C34254 _1030_/a_891_413# _0339_ 0
C34255 net16 net66 0.00969f
C34256 hold1/a_391_47# _0987_/a_891_413# 0
C34257 _0157_ clknet_1_0__leaf__0459_ 0
C34258 net83 _0793_/a_149_47# 0
C34259 _1041_/a_975_413# _0174_ 0
C34260 clknet_1_0__leaf__0460_ _0102_ 0.03988f
C34261 _0664_/a_297_47# _0284_ 0.04856f
C34262 pp[29] VPWR 0.33366f
C34263 _0229_ hold94/a_49_47# 0
C34264 _0133_ _0475_ 0
C34265 hold85/a_49_47# _1063_/a_27_47# 0
C34266 output56/a_27_47# _0355_ 0
C34267 _0985_/a_27_47# _0183_ 0
C34268 VPWR _0449_ 0.36335f
C34269 hold52/a_285_47# _0574_/a_109_297# 0
C34270 hold52/a_391_47# _0574_/a_27_297# 0.00108f
C34271 net58 _0833_/a_215_47# 0.00789f
C34272 _0195_ _0566_/a_27_47# 0
C34273 comp0.B\[6\] _0496_/a_27_47# 0.00176f
C34274 _0797_/a_207_413# net5 0.00287f
C34275 _0217_ _1018_/a_193_47# 0.03145f
C34276 net234 _1014_/a_381_47# 0
C34277 _0570_/a_109_297# _0689_/a_68_297# 0
C34278 _1007_/a_634_159# net93 0
C34279 _1007_/a_193_47# _0105_ 0.25861f
C34280 _1007_/a_891_413# _1007_/a_1017_47# 0.00617f
C34281 _0324_ _0318_ 0.00243f
C34282 net243 _1004_/a_193_47# 0.05876f
C34283 VPWR _0364_ 0.34672f
C34284 _0622_/a_193_47# _0369_ 0
C34285 clknet_1_0__leaf__0464_ net133 0.10809f
C34286 _0372_ _0181_ 0
C34287 _0837_/a_81_21# _0442_ 0.12034f
C34288 _0837_/a_368_297# _0440_ 0.00311f
C34289 _0837_/a_266_297# _0441_ 0
C34290 _0165_ hold93/a_285_47# 0.03157f
C34291 _1058_/a_381_47# net144 0
C34292 _0287_ _0369_ 0.12165f
C34293 _0126_ _1027_/a_27_47# 0
C34294 net197 _1027_/a_891_413# 0.00142f
C34295 _0178_ _0465_ 0.03464f
C34296 net48 _0762_/a_297_297# 0.0014f
C34297 VPWR _0498_/a_149_47# 0.00165f
C34298 _0625_/a_145_75# clknet_1_1__leaf__0458_ 0
C34299 clknet_1_1__leaf__0460_ _0678_/a_68_297# 0
C34300 _0397_ _0396_ 0
C34301 hold74/a_49_47# hold74/a_391_47# 0.00188f
C34302 _0557_/a_240_47# VPWR 0.00219f
C34303 _0705_/a_59_75# _0336_ 0.15543f
C34304 _0734_/a_47_47# _0734_/a_285_47# 0.01755f
C34305 _0705_/a_145_75# _0220_ 0.00127f
C34306 _0459_ _0115_ 0
C34307 _1050_/a_561_413# net11 0
C34308 _0230_ _0602_/a_113_47# 0
C34309 hold32/a_49_47# pp[1] 0
C34310 _1003_/a_381_47# _0487_ 0.00152f
C34311 acc0.A\[12\] _0187_ 0.30735f
C34312 VPWR _0110_ 0.41063f
C34313 _0107_ _0387_ 0
C34314 _0971_/a_299_297# _0181_ 0.05874f
C34315 comp0.B\[12\] net18 0.00548f
C34316 net57 _0354_ 0.0824f
C34317 net88 VPWR 0.44294f
C34318 _0268_ _0219_ 0.02316f
C34319 _1061_/a_891_413# comp0.B\[9\] 0
C34320 _0819_/a_299_297# _0659_/a_68_297# 0
C34321 net61 _0252_ 0.03392f
C34322 _0459_ _0796_/a_297_297# 0
C34323 clkbuf_0_clk/a_110_47# _1063_/a_381_47# 0
C34324 hold59/a_285_47# clkbuf_1_0__f__0461_/a_110_47# 0
C34325 acc0.A\[4\] hold1/a_285_47# 0.01328f
C34326 _0464_ _0182_ 0
C34327 _0389_ _0247_ 0.01893f
C34328 _0198_ net157 0
C34329 hold75/a_391_47# _0082_ 0
C34330 net16 _0350_ 0
C34331 _0983_/a_634_159# _0081_ 0.00555f
C34332 _0983_/a_1059_315# _0455_ 0
C34333 _0983_/a_891_413# _0454_ 0
C34334 _0328_ _0105_ 0
C34335 _1063_/a_634_159# _1063_/a_381_47# 0
C34336 _1046_/a_27_47# net174 0
C34337 _0327_ _0356_ 0.2248f
C34338 net204 _0549_/a_68_297# 0.00171f
C34339 _0555_/a_149_47# net171 0
C34340 net39 net40 0.00224f
C34341 net45 output60/a_27_47# 0.00395f
C34342 hold19/a_391_47# net221 0
C34343 _1037_/a_891_413# _0208_ 0
C34344 _0280_ _0421_ 0
C34345 _0180_ input14/a_75_212# 0
C34346 net231 _0163_ 0
C34347 net67 _0286_ 0
C34348 B[9] input22/a_75_212# 0.00186f
C34349 input32/a_75_212# B[14] 0
C34350 _0462_ _1006_/a_1059_315# 0.00535f
C34351 hold86/a_391_47# net58 0.09467f
C34352 pp[16] _0218_ 0
C34353 _0748_/a_81_21# _0748_/a_299_297# 0.08213f
C34354 _0174_ B[12] 0
C34355 _0119_ acc0.A\[20\] 0
C34356 net125 _0497_/a_150_297# 0.00138f
C34357 hold52/a_49_47# _1025_/a_1059_315# 0
C34358 _0183_ _0507_/a_109_47# 0.00145f
C34359 hold11/a_49_47# net135 0
C34360 _0536_/a_240_47# clknet_0__0464_ 0
C34361 net158 _1049_/a_381_47# 0
C34362 _0343_ _0790_/a_117_297# 0.00209f
C34363 _0216_ control0.sh 0
C34364 _1028_/a_193_47# clknet_1_1__leaf__0462_ 0.05369f
C34365 net70 VPWR 0.37789f
C34366 _0663_/a_27_413# _0345_ 0.00636f
C34367 _0201_ comp0.B\[9\] 0
C34368 net46 _0771_/a_215_297# 0
C34369 _0346_ net206 0
C34370 net96 net98 0.00106f
C34371 _0601_/a_68_297# _0600_/a_103_199# 0.001f
C34372 _0237_ _0345_ 0.0418f
C34373 _0176_ _0545_/a_68_297# 0.13312f
C34374 _0183_ hold82/a_285_47# 0
C34375 _0628_/a_109_297# acc0.A\[3\] 0.00286f
C34376 clkbuf_1_0__f__0464_/a_110_47# net11 0.0011f
C34377 _0663_/a_297_47# _0295_ 0
C34378 net111 net112 0.12329f
C34379 _1011_/a_975_413# acc0.A\[29\] 0
C34380 _0833_/a_79_21# clknet_1_1__leaf__0458_ 0.00346f
C34381 _0570_/a_109_297# net112 0
C34382 _1004_/a_193_47# _1024_/a_381_47# 0
C34383 VPWR _1010_/a_193_47# 0.34083f
C34384 _0369_ _0990_/a_1017_47# 0
C34385 net88 net48 0
C34386 _1000_/a_27_47# _1000_/a_193_47# 0.96285f
C34387 _0394_ _0352_ 0
C34388 _0241_ clknet_1_0__leaf__0457_ 0
C34389 _0080_ _0346_ 0.15478f
C34390 _1060_/a_634_159# _1060_/a_381_47# 0
C34391 _1051_/a_193_47# _0527_/a_109_297# 0
C34392 _0733_/a_544_297# _0319_ 0.00368f
C34393 _0513_/a_299_297# _0513_/a_384_47# 0
C34394 net114 _1008_/a_466_413# 0
C34395 _1028_/a_466_413# net94 0
C34396 clkbuf_0__0457_/a_110_47# hold60/a_285_47# 0.02314f
C34397 net111 acc0.A\[24\] 0
C34398 _1070_/a_193_47# net164 0
C34399 hold49/a_49_47# hold49/a_285_47# 0.22264f
C34400 _1051_/a_193_47# _0346_ 0
C34401 _1053_/a_634_159# net11 0.00577f
C34402 _0143_ _1050_/a_891_413# 0.00255f
C34403 acc0.A\[9\] _0283_ 0
C34404 hold69/a_49_47# clkbuf_0__0460_/a_110_47# 0.00242f
C34405 clknet_1_1__leaf__0463_ comp0.B\[5\] 0.03896f
C34406 hold26/a_49_47# _0176_ 0.00144f
C34407 net203 _1065_/a_634_159# 0
C34408 net163 hold62/a_285_47# 0
C34409 _0988_/a_891_413# net74 0
C34410 _0553_/a_512_297# _0174_ 0
C34411 _1067_/a_1059_315# clknet_1_1__leaf_clk 0
C34412 _0399_ _0986_/a_27_47# 0.03367f
C34413 _0501_/a_27_47# _0924_/a_27_47# 0
C34414 _0973_/a_27_297# _1063_/a_27_47# 0
C34415 _0343_ _0348_ 0.10871f
C34416 _0331_ _1011_/a_193_47# 0
C34417 pp[27] _0568_/a_373_47# 0
C34418 net56 _1011_/a_466_413# 0
C34419 VPWR _1009_/a_634_159# 0.18082f
C34420 _0579_/a_27_297# net187 0.1244f
C34421 _0367_ clknet_0__0460_ 0
C34422 hold19/a_49_47# hold19/a_285_47# 0.22264f
C34423 _0467_ control0.state\[2\] 0.0785f
C34424 hold87/a_285_47# _0345_ 0
C34425 _0280_ _0809_/a_81_21# 0
C34426 _1041_/a_891_413# _0206_ 0.00165f
C34427 _0183_ _0242_ 0.16155f
C34428 _0537_/a_68_297# _0954_/a_32_297# 0.01012f
C34429 _0982_/a_592_47# _0465_ 0
C34430 net120 _0467_ 0
C34431 _0294_ net47 0
C34432 _0118_ clkbuf_0__0457_/a_110_47# 0
C34433 _0234_ _0217_ 0
C34434 _0583_/a_27_297# _0583_/a_109_47# 0.00393f
C34435 VPWR _1014_/a_561_413# 0.00292f
C34436 _1071_/a_1059_315# VPWR 0.42713f
C34437 net15 hold7/a_49_47# 0
C34438 net243 net199 0
C34439 _0470_ _1062_/a_27_47# 0
C34440 net8 comp0.B\[5\] 0
C34441 _0985_/a_27_47# _0179_ 0.06137f
C34442 _0856_/a_215_47# _0452_ 0
C34443 clknet_1_0__leaf__0457_ _0772_/a_510_47# 0.00278f
C34444 _0984_/a_193_47# hold75/a_391_47# 0
C34445 hold39/a_285_47# VPWR 0.28958f
C34446 hold28/a_391_47# clknet_1_0__leaf__0464_ 0
C34447 acc0.A\[15\] _0507_/a_109_47# 0
C34448 _0101_ net240 0
C34449 net85 _0097_ 0.06884f
C34450 _0680_/a_80_21# clknet_0__0460_ 0
C34451 _0316_ _0318_ 0.48372f
C34452 _0500_/a_27_47# _1049_/a_634_159# 0
C34453 hold59/a_391_47# acc0.A\[1\] 0
C34454 _0216_ net157 0.4094f
C34455 _0133_ net27 0.02219f
C34456 _0479_ _0978_/a_109_297# 0.00104f
C34457 _1021_/a_592_47# _0460_ 0
C34458 acc0.A\[15\] hold82/a_285_47# 0.00389f
C34459 net36 hold71/a_391_47# 0
C34460 _0461_ _0347_ 0.02597f
C34461 net157 clknet_1_1__leaf__0464_ 0
C34462 hold20/a_285_47# net35 0.0336f
C34463 clkbuf_0__0462_/a_110_47# _0321_ 0.00993f
C34464 _0258_ _0271_ 0.34642f
C34465 _0309_ _0677_/a_285_47# 0.05006f
C34466 clknet_0__0464_ _1046_/a_27_47# 0.08671f
C34467 clkbuf_0__0464_/a_110_47# _1046_/a_891_413# 0.0036f
C34468 _0997_/a_27_47# output41/a_27_47# 0
C34469 hold35/a_391_47# acc0.A\[9\] 0.01316f
C34470 _1071_/a_27_47# clkbuf_1_0__f_clk/a_110_47# 0.01046f
C34471 clkbuf_0__0462_/a_110_47# clkbuf_0__0460_/a_110_47# 0.01215f
C34472 _0347_ _0318_ 0
C34473 net54 _1027_/a_27_47# 0.03903f
C34474 hold79/a_391_47# control0.count\[0\] 0.00177f
C34475 _1008_/a_466_413# _0365_ 0
C34476 _1008_/a_193_47# _0106_ 0.58445f
C34477 _0959_/a_80_21# _0173_ 0
C34478 output38/a_27_47# net38 0.1886f
C34479 _0558_/a_68_297# net27 0.03262f
C34480 acc0.A\[5\] _0830_/a_79_21# 0
C34481 _0999_/a_1059_315# net43 0
C34482 _0718_/a_47_47# _1030_/a_891_413# 0
C34483 _0626_/a_68_297# _0431_ 0
C34484 net175 _1048_/a_891_413# 0.01047f
C34485 net9 _1048_/a_634_159# 0.01968f
C34486 comp0.B\[11\] _1043_/a_27_47# 0
C34487 _0343_ acc0.A\[31\] 0
C34488 _0958_/a_27_47# _1062_/a_466_413# 0
C34489 net247 control0.sh 0
C34490 _0975_/a_59_75# _1068_/a_27_47# 0
C34491 net44 _0779_/a_510_47# 0
C34492 net149 _1047_/a_466_413# 0.0023f
C34493 clknet_1_0__leaf__0465_ _0527_/a_27_297# 0.00196f
C34494 hold13/a_49_47# _0472_ 0.00458f
C34495 hold13/a_391_47# _0473_ 0.00739f
C34496 pp[8] input2/a_75_212# 0
C34497 clknet_1_0__leaf__0458_ _0399_ 0.06419f
C34498 VPWR _1022_/a_466_413# 0.25404f
C34499 net59 _0568_/a_109_297# 0
C34500 _0946_/a_30_53# clknet_1_0__leaf_clk 0
C34501 _0273_ _0988_/a_27_47# 0
C34502 _0553_/a_512_297# _0208_ 0
C34503 clknet_1_1__leaf__0459_ _0993_/a_634_159# 0
C34504 acc0.A\[29\] _0334_ 0.39795f
C34505 _0993_/a_1059_315# net38 0.09458f
C34506 input22/a_75_212# hold6/a_285_47# 0
C34507 _0999_/a_27_47# _0999_/a_1059_315# 0.04875f
C34508 _0999_/a_193_47# _0999_/a_466_413# 0.07855f
C34509 _0820_/a_215_47# _0290_ 0
C34510 _0820_/a_297_297# _0401_ 0
C34511 net17 _1063_/a_27_47# 0.04311f
C34512 _0992_/a_193_47# net217 0.00155f
C34513 _0992_/a_27_47# _0422_ 0
C34514 VPWR _0771_/a_298_297# 0.19392f
C34515 _0317_ _0319_ 0.10035f
C34516 _1001_/a_27_47# net223 0.00131f
C34517 _0121_ acc0.A\[23\] 0.00684f
C34518 _0341_ _1031_/a_193_47# 0
C34519 _0340_ _1031_/a_27_47# 0
C34520 _0623_/a_109_297# clknet_1_1__leaf__0458_ 0.00295f
C34521 clknet_1_0__leaf__0465_ _0989_/a_634_159# 0
C34522 clknet_1_0__leaf__0465_ hold1/a_391_47# 0.01794f
C34523 _0457_ _0208_ 0.1464f
C34524 net120 _1034_/a_634_159# 0
C34525 _1035_/a_381_47# net25 0
C34526 _0174_ _0475_ 0
C34527 _1062_/a_634_159# _0160_ 0
C34528 input23/a_75_212# net25 0
C34529 net23 input25/a_75_212# 0
C34530 net67 _0673_/a_103_199# 0
C34531 net39 _0647_/a_285_47# 0.07468f
C34532 _0600_/a_253_297# _0345_ 0
C34533 clknet_1_0__leaf__0465_ _1061_/a_27_47# 0.00461f
C34534 hold100/a_49_47# _0635_/a_27_47# 0.00199f
C34535 _1021_/a_634_159# _1021_/a_1017_47# 0
C34536 _1021_/a_466_413# _1021_/a_592_47# 0.00553f
C34537 _1033_/a_891_413# net23 0
C34538 hold24/a_285_47# _1038_/a_1059_315# 0.01349f
C34539 _0455_ _0266_ 0
C34540 _0575_/a_27_297# _0122_ 0.11341f
C34541 _1017_/a_891_413# _0459_ 0.00503f
C34542 _0573_/a_27_47# _0566_/a_27_47# 0.03318f
C34543 net182 acc0.A\[9\] 0.31238f
C34544 _0147_ _1048_/a_381_47# 0
C34545 acc0.A\[16\] _0399_ 0.00126f
C34546 clknet_1_1__leaf__0461_ net42 0
C34547 _0179_ hold82/a_285_47# 0.00429f
C34548 _0744_/a_27_47# _0992_/a_193_47# 0
C34549 VPWR _0540_/a_51_297# 0.54899f
C34550 _0996_/a_27_47# _0302_ 0.00168f
C34551 control0.state\[1\] _0163_ 0.00315f
C34552 _0843_/a_150_297# _0350_ 0
C34553 net69 hold18/a_391_47# 0
C34554 _0459_ net146 0.00102f
C34555 _0733_/a_544_297# _0733_/a_448_47# 0.00203f
C34556 _1056_/a_193_47# acc0.A\[12\] 0.00337f
C34557 net86 _0183_ 0.00434f
C34558 _0963_/a_285_47# clk 0
C34559 _0197_ acc0.A\[15\] 0
C34560 _0481_ control0.count\[0\] 0.04254f
C34561 _1043_/a_27_47# _0202_ 0
C34562 acc0.A\[20\] _0373_ 0.00504f
C34563 net62 _0988_/a_1059_315# 0.0309f
C34564 _1011_/a_466_413# _0345_ 0
C34565 hold11/a_285_47# VPWR 0.28109f
C34566 net48 _1022_/a_466_413# 0.00182f
C34567 _1031_/a_466_413# _1013_/a_466_413# 0
C34568 _1031_/a_193_47# _1013_/a_891_413# 0
C34569 net71 net170 0
C34570 _0375_ _0378_ 0.24599f
C34571 _0216_ _0568_/a_373_47# 0.00413f
C34572 clknet_1_1__leaf__0460_ _0701_/a_80_21# 0.05128f
C34573 clknet_0__0458_ _0435_ 0
C34574 _0461_ comp0.B\[1\] 0.0017f
C34575 net157 net247 0.02616f
C34576 _0782_/a_27_47# net149 0.00275f
C34577 hold57/a_391_47# VPWR 0.18093f
C34578 _0953_/a_304_297# comp0.B\[8\] 0.00124f
C34579 _0953_/a_220_297# _0206_ 0
C34580 comp0.B\[10\] _0547_/a_68_297# 0
C34581 _0424_ _0816_/a_68_297# 0
C34582 net45 _0097_ 0.00636f
C34583 _0260_ VPWR 1.16895f
C34584 _0168_ _0978_/a_27_297# 0.15957f
C34585 net23 net240 0
C34586 VPWR _0795_/a_384_47# 0
C34587 hold26/a_285_47# _0139_ 0
C34588 hold97/a_391_47# net54 0.00509f
C34589 _0742_/a_299_297# clknet_0__0460_ 0
C34590 hold19/a_285_47# _1017_/a_193_47# 0
C34591 hold19/a_49_47# _1017_/a_634_159# 0
C34592 hold19/a_391_47# _1017_/a_27_47# 0
C34593 hold85/a_285_47# hold85/a_391_47# 0.41909f
C34594 _0780_/a_35_297# _0780_/a_285_47# 0.00723f
C34595 clknet_1_0__leaf__0465_ _0538_/a_512_297# 0
C34596 _0349_ clkbuf_1_1__f__0462_/a_110_47# 0
C34597 control0.count\[2\] _1071_/a_27_47# 0.04696f
C34598 _0984_/a_1059_315# _0399_ 0.00303f
C34599 hold78/a_391_47# _0111_ 0.00188f
C34600 _1055_/a_193_47# _0189_ 0
C34601 net160 _0209_ 0
C34602 hold47/a_49_47# _1050_/a_27_47# 0.00196f
C34603 net69 _0195_ 0
C34604 VPWR _1067_/a_891_413# 0.20515f
C34605 _0465_ _0347_ 0.00258f
C34606 net176 _1022_/a_27_47# 0
C34607 _0222_ _1023_/a_27_47# 0.001f
C34608 _1050_/a_466_413# _0186_ 0.0149f
C34609 acc0.A\[14\] _0263_ 0.11938f
C34610 hold31/a_49_47# VPWR 0.28488f
C34611 acc0.A\[14\] clkload4/Y 0
C34612 _0725_/a_80_21# _0707_/a_75_199# 0
C34613 hold28/a_49_47# hold28/a_391_47# 0.00188f
C34614 net17 _1062_/a_1059_315# 0
C34615 hold99/a_285_47# net38 0.10008f
C34616 hold13/a_285_47# _0135_ 0
C34617 _1033_/a_466_413# clknet_1_0__leaf__0461_ 0
C34618 net181 net2 0.00814f
C34619 _0717_/a_209_297# VPWR 0.20087f
C34620 _1019_/a_193_47# _0869_/a_27_47# 0
C34621 _0359_ _1007_/a_193_47# 0
C34622 _0324_ _1007_/a_27_47# 0.00174f
C34623 _0459_ net223 0
C34624 _0475_ _0208_ 0.13588f
C34625 _0346_ _0405_ 0.08979f
C34626 _0390_ _0771_/a_298_297# 0.00138f
C34627 _0243_ _0771_/a_382_47# 0
C34628 acc0.A\[7\] A[4] 0.01051f
C34629 _0780_/a_35_297# _0677_/a_47_47# 0
C34630 _0343_ _0274_ 0
C34631 hold14/a_49_47# net27 0
C34632 _0243_ _0310_ 0
C34633 net243 VPWR 0.23628f
C34634 _1038_/a_27_47# _0554_/a_68_297# 0
C34635 input27/a_75_212# B[4] 0.19633f
C34636 clkbuf_1_0__f__0457_/a_110_47# _0713_/a_27_47# 0
C34637 comp0.B\[15\] _0563_/a_240_47# 0
C34638 hold100/a_49_47# _0850_/a_68_297# 0
C34639 _1047_/a_381_47# _0145_ 0.12489f
C34640 _1000_/a_193_47# acc0.A\[19\] 0
C34641 _0228_ _0765_/a_79_21# 0
C34642 _0338_ _0568_/a_27_297# 0
C34643 _0707_/a_75_199# _0128_ 0
C34644 clknet_1_0__leaf_clk _0487_ 0
C34645 net118 hold40/a_391_47# 0
C34646 _0479_ _0480_ 0.20815f
C34647 hold46/a_285_47# comp0.B\[10\] 0
C34648 _0179_ _0197_ 0.02185f
C34649 net222 _0219_ 0.17453f
C34650 VPWR output60/a_27_47# 0.28045f
C34651 VPWR _0768_/a_109_297# 0.00393f
C34652 _0247_ _0612_/a_59_75# 0
C34653 _0557_/a_51_297# _1036_/a_1059_315# 0.00131f
C34654 clkload3/Y _0309_ 0
C34655 _0587_/a_27_47# _0097_ 0
C34656 hold86/a_285_47# net47 0
C34657 _0546_/a_51_297# _1040_/a_193_47# 0
C34658 net234 acc0.A\[0\] 0
C34659 _0710_/a_109_297# _0219_ 0.01264f
C34660 _0567_/a_109_47# acc0.A\[30\] 0.00125f
C34661 net232 _0959_/a_80_21# 0
C34662 _1004_/a_193_47# _0378_ 0.0013f
C34663 _0620_/a_113_47# acc0.A\[8\] 0
C34664 clkbuf_1_1__f__0462_/a_110_47# _0701_/a_209_297# 0.0016f
C34665 _0513_/a_299_297# net4 0
C34666 acc0.A\[8\] _0989_/a_27_47# 0.03699f
C34667 _0753_/a_79_21# _0374_ 0.01234f
C34668 hold54/a_285_47# _0563_/a_51_297# 0
C34669 hold68/a_49_47# _1022_/a_27_47# 0
C34670 _0328_ _0359_ 0.03204f
C34671 net89 hold3/a_391_47# 0
C34672 _0996_/a_27_47# net6 0
C34673 acc0.A\[12\] clkbuf_1_1__f__0459_/a_110_47# 0.00277f
C34674 _0305_ acc0.A\[17\] 0.42256f
C34675 _0712_/a_297_297# _0341_ 0.04484f
C34676 _0712_/a_79_21# _0340_ 0.01855f
C34677 net168 net15 0.33847f
C34678 net190 net156 0.02805f
C34679 _0119_ net107 0.00102f
C34680 net69 _0852_/a_35_297# 0
C34681 _0387_ _0306_ 0.00347f
C34682 _0544_/a_51_297# _0544_/a_149_47# 0.02487f
C34683 _0733_/a_448_47# _0317_ 0
C34684 _0956_/a_220_297# control0.reset 0.00107f
C34685 _0747_/a_79_21# _0460_ 0.01047f
C34686 VPWR _0524_/a_27_297# 0.1903f
C34687 input28/a_75_212# B[6] 0.00205f
C34688 _1034_/a_634_159# _1034_/a_466_413# 0.23992f
C34689 _1034_/a_193_47# _1034_/a_1059_315# 0.03405f
C34690 _1034_/a_27_47# _1034_/a_891_413# 0.03089f
C34691 _0536_/a_51_297# _0536_/a_240_47# 0.03076f
C34692 _0581_/a_27_297# clknet_1_0__leaf__0461_ 0.0082f
C34693 net162 _1030_/a_1059_315# 0.00184f
C34694 output59/a_27_47# acc0.A\[29\] 0.01112f
C34695 _0497_/a_68_297# _0497_/a_150_297# 0.00477f
C34696 _1021_/a_634_159# acc0.A\[21\] 0
C34697 net168 _1053_/a_1059_315# 0.05664f
C34698 net14 _1053_/a_193_47# 0
C34699 _0430_ _0826_/a_301_297# 0
C34700 net78 _0346_ 0
C34701 _0626_/a_68_297# _0269_ 0
C34702 clknet_0__0465_ _0346_ 0.16377f
C34703 _0427_ net66 0.00223f
C34704 _0982_/a_381_47# clknet_1_0__leaf__0461_ 0.001f
C34705 _0380_ acc0.A\[23\] 0.14263f
C34706 output64/a_27_47# net58 0.09274f
C34707 _0850_/a_150_297# _0446_ 0
C34708 _0217_ _0855_/a_384_47# 0
C34709 _0183_ _0855_/a_81_21# 0.01347f
C34710 _0662_/a_81_21# _0347_ 0
C34711 _0179_ _0153_ 0.02228f
C34712 _1013_/a_27_47# _0219_ 0.02945f
C34713 _0516_/a_109_47# acc0.A\[9\] 0.00185f
C34714 _0397_ net43 0
C34715 net69 _0081_ 0
C34716 control0.state\[0\] _1066_/a_193_47# 0
C34717 _0570_/a_27_297# _0570_/a_109_47# 0.00393f
C34718 clkbuf_0__0464_/a_110_47# _1045_/a_466_413# 0
C34719 net100 net157 0
C34720 _1063_/a_891_413# _0161_ 0.04588f
C34721 _0086_ _0988_/a_27_47# 0.09972f
C34722 net235 _0988_/a_466_413# 0
C34723 _0225_ _0756_/a_377_297# 0.00168f
C34724 _0607_/a_27_297# _0219_ 0
C34725 control0.state\[1\] _1068_/a_27_47# 0
C34726 control0.state\[0\] _1068_/a_193_47# 0
C34727 net65 clknet_0__0465_ 0
C34728 VPWR _1026_/a_634_159# 0.2003f
C34729 net138 hold83/a_391_47# 0.00426f
C34730 hold68/a_391_47# _0216_ 0.00139f
C34731 control0.count\[3\] _1072_/a_466_413# 0.03278f
C34732 _0483_ _1072_/a_193_47# 0
C34733 _0343_ net43 0.03283f
C34734 hold88/a_391_47# clknet_1_1__leaf__0458_ 0
C34735 _0217_ output46/a_27_47# 0
C34736 net78 _0992_/a_466_413# 0
C34737 output43/a_27_47# output41/a_27_47# 0
C34738 _0305_ net5 0.02876f
C34739 VPWR _1024_/a_381_47# 0.07565f
C34740 hold32/a_49_47# hold32/a_285_47# 0.22264f
C34741 _0399_ hold91/a_285_47# 0.03133f
C34742 _0216_ _0462_ 0.04276f
C34743 _0258_ clknet_1_0__leaf__0465_ 0.01677f
C34744 hold13/a_285_47# hold13/a_391_47# 0.41909f
C34745 _0172_ _0498_/a_512_297# 0.0016f
C34746 _0585_/a_373_47# net149 0
C34747 net203 _0563_/a_240_47# 0.04112f
C34748 _0517_/a_81_21# _0517_/a_384_47# 0.00138f
C34749 _0211_ _0175_ 0.09974f
C34750 _0999_/a_27_47# _0397_ 0
C34751 _0361_ _0691_/a_68_297# 0.00791f
C34752 hold97/a_285_47# VPWR 0.29024f
C34753 hold75/a_49_47# _0454_ 0
C34754 clkbuf_0__0465_/a_110_47# _0465_ 0.3209f
C34755 VPWR _1048_/a_975_413# 0.00517f
C34756 clknet_1_0__leaf__0460_ _1005_/a_193_47# 0.01036f
C34757 net198 _0203_ 0.09747f
C34758 control0.state\[0\] _0478_ 0.00132f
C34759 net76 _0428_ 0
C34760 _1017_/a_27_47# _1017_/a_466_413# 0.26005f
C34761 _1017_/a_193_47# _1017_/a_634_159# 0.12262f
C34762 _0195_ net102 0
C34763 _1058_/a_193_47# _0512_/a_27_297# 0
C34764 pp[27] _0725_/a_303_47# 0
C34765 output58/a_27_47# _0831_/a_35_297# 0
C34766 _0473_ _1046_/a_1059_315# 0.01442f
C34767 net248 _0835_/a_215_47# 0
C34768 hold101/a_391_47# _0255_ 0
C34769 net190 acc0.A\[26\] 0.02776f
C34770 _1004_/a_891_413# net110 0
C34771 _1000_/a_634_159# _1000_/a_1017_47# 0
C34772 _1000_/a_466_413# _1000_/a_592_47# 0.00553f
C34773 _0507_/a_27_297# _0507_/a_109_297# 0.17136f
C34774 _0600_/a_337_297# clknet_1_0__leaf__0460_ 0.00148f
C34775 _1060_/a_381_47# net146 0
C34776 _1060_/a_891_413# _0158_ 0.00122f
C34777 _0993_/a_466_413# _0281_ 0
C34778 _1051_/a_561_413# net154 0
C34779 _1051_/a_1059_315# net11 0.02442f
C34780 net64 _0989_/a_27_47# 0
C34781 _0176_ hold51/a_285_47# 0.003f
C34782 net118 comp0.B\[0\] 0
C34783 hold43/a_391_47# acc0.A\[28\] 0.06999f
C34784 _0346_ _0815_/a_199_47# 0
C34785 VPWR net164 0.16578f
C34786 _0427_ _0350_ 0
C34787 _0671_/a_113_297# acc0.A\[15\] 0.06918f
C34788 net230 net14 0.06397f
C34789 _1072_/a_381_47# VPWR 0.07359f
C34790 _0399_ _0288_ 0.00505f
C34791 hold55/a_391_47# clknet_1_0__leaf__0457_ 0.02172f
C34792 clkbuf_0__0463_/a_110_47# _1061_/a_634_159# 0
C34793 _0786_/a_217_297# net228 0.00686f
C34794 acc0.A\[17\] _0675_/a_150_297# 0
C34795 comp0.B\[10\] net127 0
C34796 _0536_/a_51_297# _1046_/a_27_47# 0.00704f
C34797 _0343_ _0368_ 0.05351f
C34798 _0625_/a_145_75# _0218_ 0
C34799 net208 acc0.A\[30\] 0.00818f
C34800 _0174_ _0136_ 0.04431f
C34801 comp0.B\[10\] _0543_/a_150_297# 0
C34802 _0763_/a_193_47# _0345_ 0
C34803 _0287_ _0817_/a_81_21# 0
C34804 _0289_ _0817_/a_266_297# 0
C34805 _0165_ _1063_/a_27_47# 0
C34806 net240 _1063_/a_466_413# 0
C34807 _0346_ _0849_/a_215_47# 0
C34808 _0582_/a_27_297# _0347_ 0.00581f
C34809 _0347_ _1007_/a_27_47# 0.00118f
C34810 net27 _0208_ 0.08811f
C34811 _0234_ _0755_/a_109_297# 0
C34812 _0233_ _0618_/a_79_21# 0
C34813 _0343_ _0618_/a_215_47# 0.00458f
C34814 _0640_/a_215_297# _0824_/a_59_75# 0.00322f
C34815 clkbuf_1_0__f__0457_/a_110_47# _0579_/a_109_297# 0
C34816 hold55/a_49_47# _0457_ 0.01072f
C34817 _0750_/a_27_47# _0750_/a_181_47# 0.00401f
C34818 _1050_/a_634_159# _1050_/a_466_413# 0.23992f
C34819 _1050_/a_193_47# _1050_/a_1059_315# 0.03405f
C34820 _1050_/a_27_47# _1050_/a_891_413# 0.03224f
C34821 _0179_ _0990_/a_27_47# 0
C34822 _0643_/a_103_199# VPWR 0.43893f
C34823 VPWR _0366_ 0.64641f
C34824 _1019_/a_466_413# clknet_1_0__leaf__0457_ 0
C34825 hold50/a_49_47# hold50/a_391_47# 0.00188f
C34826 _0432_ _0826_/a_27_53# 0
C34827 _0294_ _0775_/a_297_297# 0
C34828 _0221_ _1011_/a_1059_315# 0.00463f
C34829 _0958_/a_27_47# _0958_/a_109_47# 0.00578f
C34830 hold21/a_285_47# acc0.A\[7\] 0.07568f
C34831 _0179_ _1049_/a_975_413# 0.00127f
C34832 clknet_1_1__leaf__0463_ _1065_/a_381_47# 0.0013f
C34833 _1051_/a_1059_315# hold7/a_391_47# 0
C34834 _1051_/a_891_413# hold7/a_285_47# 0
C34835 _0157_ _0345_ 0
C34836 _1059_/a_1017_47# _0219_ 0
C34837 net55 _0328_ 0
C34838 _0786_/a_80_21# _0347_ 0
C34839 clknet_1_0__leaf__0462_ hold90/a_49_47# 0.00235f
C34840 _0999_/a_466_413# _1012_/a_466_413# 0
C34841 clkbuf_1_0__f__0460_/a_110_47# _0374_ 0
C34842 net66 net142 0
C34843 _0465_ _0824_/a_59_75# 0
C34844 B[4] net17 0
C34845 _0458_ _0261_ 0.07425f
C34846 _0718_/a_377_297# VPWR 0.00482f
C34847 _0997_/a_975_413# net41 0.00174f
C34848 _0222_ _0345_ 0.04843f
C34849 _0998_/a_193_47# net43 0.00153f
C34850 clknet_0__0463_ net201 0.02881f
C34851 net158 net157 0.06325f
C34852 _0748_/a_81_21# _0246_ 0
C34853 _1071_/a_975_413# clknet_0_clk 0
C34854 _1054_/a_193_47# _1052_/a_193_47# 0
C34855 _1054_/a_27_47# _1052_/a_634_159# 0
C34856 net226 clk 0.00175f
C34857 output54/a_27_47# net156 0
C34858 net224 _1009_/a_466_413# 0
C34859 hold33/a_391_47# VPWR 0.16759f
C34860 clknet_1_1__leaf__0459_ _0788_/a_150_297# 0
C34861 _0982_/a_27_47# net149 0.0026f
C34862 _1039_/a_634_159# clkbuf_0__0463_/a_110_47# 0.00125f
C34863 net9 net134 0
C34864 acc0.A\[27\] net56 0
C34865 _0538_/a_240_47# _1044_/a_193_47# 0
C34866 acc0.A\[17\] _0181_ 0.01885f
C34867 _1056_/a_27_47# _0179_ 0.09661f
C34868 acc0.A\[14\] _1060_/a_891_413# 0.00774f
C34869 hold65/a_49_47# hold65/a_391_47# 0.00188f
C34870 clknet_1_1__leaf__0464_ net13 0
C34871 _1020_/a_1059_315# net187 0.01901f
C34872 _0958_/a_27_47# _0160_ 0
C34873 _0477_ _1062_/a_466_413# 0.00802f
C34874 _1001_/a_27_47# clkbuf_0__0457_/a_110_47# 0
C34875 pp[28] _0725_/a_209_47# 0
C34876 _0486_ _1068_/a_891_413# 0.03867f
C34877 net1 control0.state\[2\] 0.05667f
C34878 hold27/a_391_47# net174 0.13013f
C34879 _0998_/a_1059_315# _0406_ 0
C34880 hold58/a_391_47# _1036_/a_193_47# 0
C34881 _0606_/a_392_297# _0460_ 0
C34882 _0973_/a_27_297# _0973_/a_373_47# 0.01338f
C34883 _0531_/a_109_47# clknet_1_1__leaf__0457_ 0.00121f
C34884 net149 _0145_ 0.07904f
C34885 VPWR net151 0.31096f
C34886 _0257_ acc0.A\[8\] 0
C34887 acc0.A\[12\] clknet_1_1__leaf__0465_ 0.58544f
C34888 hold46/a_49_47# _1046_/a_27_47# 0
C34889 _0946_/a_112_297# clk 0
C34890 _1033_/a_1059_315# _0173_ 0.00163f
C34891 _0343_ _1000_/a_1059_315# 0
C34892 acc0.A\[10\] hold81/a_285_47# 0.00167f
C34893 VPWR _0097_ 0.57632f
C34894 _0136_ _0208_ 0.06925f
C34895 _0999_/a_891_413# _0999_/a_1017_47# 0.00617f
C34896 _0455_ _0399_ 0.31872f
C34897 _0999_/a_634_159# net85 0.00115f
C34898 clkbuf_1_1__f__0459_/a_110_47# net42 0.04988f
C34899 clkbuf_1_0__f__0458_/a_110_47# net69 0
C34900 _0684_/a_59_75# clknet_0__0462_ 0.00136f
C34901 _1001_/a_634_159# _1019_/a_891_413# 0.00167f
C34902 _1001_/a_466_413# _1019_/a_1059_315# 0.00283f
C34903 _1017_/a_592_47# _0115_ 0
C34904 hold76/a_49_47# clkbuf_1_0__f__0461_/a_110_47# 0.02051f
C34905 _0772_/a_79_21# net223 0.10426f
C34906 VPWR _0993_/a_381_47# 0.09733f
C34907 net235 _0186_ 0.03308f
C34908 _1054_/a_1059_315# net148 0
C34909 _1054_/a_193_47# net12 0
C34910 net124 net7 0
C34911 _0752_/a_300_297# _0752_/a_384_47# 0
C34912 net58 _0268_ 0.04405f
C34913 clkbuf_1_1__f__0461_/a_110_47# _0307_ 0.07447f
C34914 _0663_/a_297_47# _0346_ 0.00238f
C34915 hold68/a_391_47# _1024_/a_193_47# 0
C34916 _0298_ hold91/a_391_47# 0
C34917 clknet_1_0__leaf__0462_ _1007_/a_381_47# 0.00496f
C34918 _0322_ _0737_/a_35_297# 0
C34919 _0697_/a_472_297# _0321_ 0.00128f
C34920 _0697_/a_300_47# _0360_ 0
C34921 _0697_/a_80_21# _0364_ 0
C34922 _0270_ _0186_ 0.09663f
C34923 _0207_ _0546_/a_51_297# 0
C34924 _0983_/a_1059_315# _0217_ 0
C34925 _0775_/a_79_21# _0775_/a_215_47# 0.04584f
C34926 _0331_ _0321_ 0
C34927 output66/a_27_47# A[11] 0
C34928 _0186_ _0987_/a_466_413# 0
C34929 _0327_ _0737_/a_35_297# 0
C34930 net57 _0353_ 0.04803f
C34931 clkbuf_1_1__f__0463_/a_110_47# _0564_/a_68_297# 0
C34932 hold74/a_285_47# net45 0.004f
C34933 _0350_ net142 0
C34934 _1043_/a_193_47# _0542_/a_240_47# 0
C34935 _0556_/a_68_297# _1036_/a_634_159# 0
C34936 _0458_ _0509_/a_27_47# 0.02226f
C34937 _1021_/a_592_47# _0119_ 0.00164f
C34938 hold24/a_391_47# net172 0
C34939 net199 acc0.A\[24\] 0.23051f
C34940 _0181_ net5 0.23186f
C34941 _0212_ input25/a_75_212# 0
C34942 _1033_/a_27_47# net17 0
C34943 _0961_/a_113_297# control0.state\[2\] 0
C34944 _0180_ _0087_ 0
C34945 hold34/a_391_47# acc0.A\[11\] 0
C34946 _1016_/a_193_47# _0459_ 0.00442f
C34947 _0648_/a_109_297# _0278_ 0.00379f
C34948 _0255_ _0369_ 0
C34949 clknet_1_1__leaf__0460_ _1012_/a_27_47# 0.0024f
C34950 hold17/a_391_47# _0480_ 0
C34951 hold17/a_285_47# net164 0.00856f
C34952 clknet_1_1__leaf__0460_ _0330_ 0.49956f
C34953 _0996_/a_891_413# _0409_ 0
C34954 hold48/a_391_47# VPWR 0.25874f
C34955 _0237_ hold94/a_391_47# 0
C34956 VPWR _0790_/a_285_47# 0
C34957 _0160_ _0132_ 0
C34958 _0416_ _0402_ 0
C34959 _1002_/a_466_413# clknet_1_0__leaf__0460_ 0.00232f
C34960 net48 net151 0.20758f
C34961 _0401_ _0810_/a_113_47# 0
C34962 output54/a_27_47# acc0.A\[26\] 0.00685f
C34963 _1006_/a_891_413# _0219_ 0
C34964 acc0.A\[9\] _0345_ 0.04574f
C34965 _1003_/a_27_47# _0468_ 0
C34966 _0814_/a_27_47# acc0.A\[9\] 0.09748f
C34967 pp[12] input5/a_75_212# 0.00187f
C34968 _0467_ _1068_/a_561_413# 0
C34969 _0120_ _0225_ 0
C34970 _0510_/a_27_297# acc0.A\[11\] 0
C34971 _0210_ _0175_ 0.00134f
C34972 hold100/a_49_47# hold100/a_285_47# 0.22264f
C34973 hold83/a_285_47# hold83/a_391_47# 0.41909f
C34974 _0985_/a_634_159# _0985_/a_381_47# 0
C34975 _0295_ _0288_ 0.00552f
C34976 comp0.B\[2\] clknet_0__0463_ 0.0205f
C34977 _0650_/a_68_297# clknet_1_1__leaf__0465_ 0
C34978 _0183_ hold29/a_49_47# 0
C34979 _0217_ hold29/a_391_47# 0
C34980 acc0.A\[22\] hold29/a_285_47# 0.00427f
C34981 _0563_/a_51_297# _0562_/a_68_297# 0
C34982 hold19/a_49_47# net103 0.03336f
C34983 _0973_/a_373_47# net17 0
C34984 _1018_/a_634_159# _1018_/a_1059_315# 0
C34985 _1018_/a_27_47# _1018_/a_381_47# 0.05761f
C34986 _1018_/a_193_47# _1018_/a_891_413# 0.19226f
C34987 clknet_1_0__leaf__0465_ _0143_ 0.01623f
C34988 _0794_/a_27_47# net6 0
C34989 _0459_ clkbuf_0__0457_/a_110_47# 0
C34990 _0985_/a_27_47# _1049_/a_891_413# 0
C34991 _0985_/a_193_47# _1049_/a_1059_315# 0
C34992 comp0.B\[14\] _1046_/a_27_47# 0
C34993 net50 _1022_/a_891_413# 0.00182f
C34994 _0642_/a_215_297# _0273_ 0.10053f
C34995 hold28/a_391_47# clkbuf_1_0__f__0464_/a_110_47# 0.00837f
C34996 net213 net46 0
C34997 _0982_/a_193_47# _0982_/a_634_159# 0.11072f
C34998 _0982_/a_27_47# _0982_/a_466_413# 0.27314f
C34999 _0275_ _0990_/a_891_413# 0
C35000 net45 _0583_/a_109_297# 0
C35001 _0343_ _1018_/a_193_47# 0
C35002 _1049_/a_27_47# _1049_/a_634_159# 0.14145f
C35003 _0249_ clkbuf_1_0__f__0460_/a_110_47# 0.01247f
C35004 _0983_/a_634_159# acc0.A\[15\] 0.00213f
C35005 clknet_1_1__leaf__0460_ _0732_/a_209_297# 0.01016f
C35006 clknet_1_1__leaf_clk _0951_/a_368_53# 0
C35007 _0159_ _0913_/a_27_47# 0.11119f
C35008 _0304_ _0670_/a_297_297# 0
C35009 _0131_ clknet_1_0__leaf__0461_ 0.00159f
C35010 net64 _0257_ 0
C35011 _0282_ acc0.A\[10\] 0.01839f
C35012 net221 net206 0
C35013 _0672_/a_79_21# _0302_ 0
C35014 VPWR _0689_/a_68_297# 0.15125f
C35015 _0753_/a_79_21# _0231_ 0
C35016 _0753_/a_297_297# _0233_ 0.04566f
C35017 _0383_ _0754_/a_51_297# 0
C35018 net68 _1047_/a_1059_315# 0
C35019 _0249_ _0250_ 0
C35020 _0530_/a_384_47# _0197_ 0
C35021 hold44/a_391_47# _0216_ 0.0183f
C35022 VPWR _0378_ 0.40471f
C35023 _0644_/a_285_47# _0301_ 0.00568f
C35024 net180 net173 0.00107f
C35025 _1054_/a_27_47# A[8] 0
C35026 _1054_/a_466_413# input15/a_75_212# 0
C35027 hold27/a_391_47# clknet_0__0464_ 0
C35028 _1019_/a_634_159# _0586_/a_27_47# 0
C35029 hold98/a_285_47# hold98/a_391_47# 0.41909f
C35030 VPWR _1027_/a_1017_47# 0
C35031 hold46/a_391_47# net153 0
C35032 hold11/a_49_47# _0172_ 0.00109f
C35033 _0218_ _0391_ 0.27834f
C35034 hold56/a_285_47# net23 0
C35035 acc0.A\[27\] _0345_ 0.02634f
C35036 _1066_/a_27_47# _1066_/a_634_159# 0.14145f
C35037 net101 _0195_ 0.00266f
C35038 net56 _1010_/a_193_47# 0.00253f
C35039 _0837_/a_81_21# acc0.A\[3\] 0
C35040 net45 _0999_/a_634_159# 0.00576f
C35041 _0997_/a_381_47# _0408_ 0
C35042 VPWR _1052_/a_466_413# 0.24072f
C35043 _0328_ _0325_ 0.03972f
C35044 _0833_/a_79_21# _0833_/a_215_47# 0.04584f
C35045 _1031_/a_193_47# acc0.A\[30\] 0.00405f
C35046 _0338_ _0128_ 0.00291f
C35047 _1023_/a_27_47# _1022_/a_466_413# 0
C35048 _0967_/a_215_297# clk 0
C35049 _1056_/a_381_47# acc0.A\[10\] 0.00116f
C35050 _1068_/a_27_47# _1068_/a_634_159# 0.13601f
C35051 net8 _1040_/a_634_159# 0
C35052 _0429_ acc0.A\[8\] 0
C35053 _0176_ _0563_/a_240_47# 0
C35054 _0181_ acc0.A\[11\] 0.16068f
C35055 hold100/a_391_47# _0446_ 0.01551f
C35056 _0677_/a_377_297# acc0.A\[17\] 0.00147f
C35057 _0205_ _1040_/a_891_413# 0
C35058 net152 _1040_/a_466_413# 0
C35059 net32 _1040_/a_634_159# 0
C35060 _0487_ _1063_/a_381_47# 0
C35061 _0218_ _0581_/a_27_297# 0
C35062 clknet_1_0__leaf__0457_ _0352_ 0.07187f
C35063 clkbuf_1_1__f__0464_/a_110_47# _1045_/a_634_159# 0
C35064 _0584_/a_27_297# clknet_1_1__leaf__0457_ 0
C35065 acc0.A\[14\] _0218_ 0.03804f
C35066 hold58/a_285_47# comp0.B\[5\] 0.03331f
C35067 _0649_/a_113_47# _0369_ 0
C35068 net55 _0108_ 0.04186f
C35069 _0720_/a_68_297# _0350_ 0.19023f
C35070 pp[9] _0512_/a_27_297# 0.03736f
C35071 _0804_/a_215_47# _0279_ 0.03739f
C35072 _1032_/a_193_47# net23 0.0358f
C35073 _0449_ _0345_ 0
C35074 net36 hold18/a_285_47# 0
C35075 _0123_ _0105_ 0
C35076 _0222_ net52 0.00267f
C35077 _0346_ _0991_/a_592_47# 0.00131f
C35078 _0478_ _1068_/a_193_47# 0
C35079 _0344_ _0341_ 0.02206f
C35080 clknet_1_0__leaf__0464_ _0987_/a_592_47# 0
C35081 hold78/a_285_47# _0342_ 0
C35082 output55/a_27_47# _0221_ 0.02224f
C35083 hold53/a_49_47# hold53/a_285_47# 0.22264f
C35084 _0544_/a_240_47# net18 0.05798f
C35085 _0544_/a_245_297# _0140_ 0
C35086 _0345_ _0364_ 0.1987f
C35087 net162 VPWR 0.41239f
C35088 input13/a_75_212# A[6] 0.19026f
C35089 _0519_/a_81_21# net65 0
C35090 _0241_ _0246_ 0.09952f
C35091 _0625_/a_59_75# net63 0.16365f
C35092 _0343_ _0708_/a_68_297# 0
C35093 VPWR _0658_/a_113_47# 0
C35094 output66/a_27_47# net66 0.2056f
C35095 VPWR _0194_ 0.42534f
C35096 _1051_/a_27_47# _0186_ 0.00859f
C35097 _0269_ _0631_/a_109_297# 0
C35098 _0536_/a_512_297# _0144_ 0
C35099 _0557_/a_245_297# net26 0
C35100 hold6/a_49_47# net198 0.01442f
C35101 _0116_ clknet_1_0__leaf__0461_ 0.0477f
C35102 net238 _0094_ 0.06746f
C35103 net48 _0378_ 0
C35104 acc0.A\[16\] _0306_ 0.10459f
C35105 B[2] B[4] 0.18737f
C35106 _0341_ _0709_/a_113_47# 0.00995f
C35107 net239 hold95/a_391_47# 0
C35108 _0169_ _0976_/a_76_199# 0
C35109 _0979_/a_27_297# _0488_ 0.13674f
C35110 _0464_ net7 0
C35111 clknet_1_1__leaf__0460_ net190 0
C35112 net43 _0793_/a_51_297# 0.0342f
C35113 _0254_ clkbuf_0__0465_/a_110_47# 0.07929f
C35114 _0243_ control0.add 0.02087f
C35115 hold85/a_391_47# _0477_ 0.00225f
C35116 _0789_/a_201_297# net6 0.04711f
C35117 hold89/a_49_47# control0.count\[0\] 0
C35118 _0787_/a_80_21# net246 0
C35119 clknet_0__0464_ _1045_/a_592_47# 0
C35120 clkbuf_0__0464_/a_110_47# net184 0
C35121 _0534_/a_81_21# _1047_/a_634_159# 0
C35122 _0534_/a_299_297# _1047_/a_193_47# 0.00165f
C35123 _0176_ _1061_/a_193_47# 0
C35124 _0346_ _1006_/a_27_47# 0.09677f
C35125 _0179_ _0293_ 0
C35126 net167 _0468_ 0
C35127 VPWR net112 0.62454f
C35128 net71 _0846_/a_51_297# 0
C35129 _0745_/a_193_47# _0460_ 0
C35130 hold29/a_285_47# _0379_ 0
C35131 _0783_/a_79_21# _0097_ 0
C35132 comp0.B\[8\] _0206_ 0.02907f
C35133 input2/a_75_212# A[10] 0.22679f
C35134 _1001_/a_1059_315# _0352_ 0.0013f
C35135 pp[30] _1031_/a_466_413# 0.00148f
C35136 VPWR acc0.A\[24\] 0.89349f
C35137 net143 _0186_ 0
C35138 _0346_ _0986_/a_27_47# 0
C35139 _0999_/a_27_47# _0793_/a_51_297# 0
C35140 hold89/a_391_47# _0974_/a_79_199# 0.00754f
C35141 hold89/a_285_47# _0974_/a_222_93# 0
C35142 _0172_ _0159_ 0.12527f
C35143 _0805_/a_27_47# _0808_/a_81_21# 0
C35144 _1071_/a_381_47# _0466_ 0.00954f
C35145 _0217_ _0266_ 0.14962f
C35146 _1021_/a_193_47# _0352_ 0
C35147 _0389_ _0248_ 0.02509f
C35148 _0993_/a_891_413# _0286_ 0
C35149 hold38/a_49_47# VPWR 0.30603f
C35150 net81 _0995_/a_891_413# 0
C35151 hold26/a_285_47# _0954_/a_32_297# 0
C35152 hold77/a_285_47# _1009_/a_1059_315# 0.0054f
C35153 _0152_ _0437_ 0
C35154 _0476_ _1062_/a_634_159# 0
C35155 _1017_/a_193_47# net103 0.15496f
C35156 _1017_/a_1059_315# _1017_/a_1017_47# 0
C35157 _0487_ _1062_/a_1017_47# 0.00125f
C35158 _0947_/a_109_297# VPWR 0.00653f
C35159 hold13/a_285_47# _0555_/a_240_47# 0
C35160 _0343_ _0234_ 0.00669f
C35161 net64 _0429_ 0
C35162 _0430_ _0251_ 0.01652f
C35163 clknet_1_0__leaf__0459_ _0790_/a_285_47# 0
C35164 _0429_ _0621_/a_117_297# 0
C35165 clkbuf_1_1__f__0463_/a_110_47# _1015_/a_1059_315# 0
C35166 net70 _0345_ 0
C35167 control0.state\[0\] clkbuf_1_1__f_clk/a_110_47# 0.00168f
C35168 _0126_ hold50/a_391_47# 0
C35169 _0507_/a_373_47# net5 0.00301f
C35170 _0507_/a_109_297# _0185_ 0.00169f
C35171 _1000_/a_381_47# net45 0.00111f
C35172 _0305_ net84 0
C35173 _0514_/a_109_47# _0186_ 0.00271f
C35174 _0804_/a_79_21# _0092_ 0.0499f
C35175 _0804_/a_215_47# _0416_ 0.00549f
C35176 clkbuf_0__0463_/a_110_47# net147 0
C35177 net44 _0780_/a_35_297# 0.00908f
C35178 _0476_ _0561_/a_512_297# 0.00209f
C35179 _1033_/a_634_159# _1033_/a_381_47# 0
C35180 _0521_/a_81_21# _0192_ 0.20787f
C35181 _0200_ _1046_/a_1059_315# 0.06303f
C35182 hold36/a_285_47# _0142_ 0
C35183 _0758_/a_215_47# net51 0.00208f
C35184 _0231_ clkbuf_1_0__f__0460_/a_110_47# 0.00342f
C35185 _0343_ clknet_0__0460_ 0
C35186 _1012_/a_634_159# _1012_/a_381_47# 0
C35187 _1039_/a_193_47# _0176_ 0.01887f
C35188 hold55/a_285_47# _1033_/a_27_47# 0
C35189 _0196_ _0527_/a_373_47# 0
C35190 net240 _0161_ 0.10119f
C35191 _0148_ _0527_/a_27_297# 0.01582f
C35192 hold23/a_49_47# _0186_ 0.01052f
C35193 _0115_ _0347_ 0
C35194 _0216_ _0312_ 0
C35195 net36 hold25/a_49_47# 0.02967f
C35196 _0401_ _0992_/a_592_47# 0
C35197 _0512_/a_373_47# _0186_ 0
C35198 _0285_ _0807_/a_150_297# 0
C35199 _0216_ _1031_/a_561_413# 0
C35200 _0195_ _1031_/a_592_47# 0
C35201 _0107_ _1009_/a_1059_315# 0
C35202 _0231_ _0250_ 0.037f
C35203 net1 net118 0
C35204 _0430_ net58 0
C35205 comp0.B\[8\] _1046_/a_1059_315# 0
C35206 _0476_ _0473_ 0
C35207 acc0.A\[8\] clknet_1_1__leaf__0458_ 0.3491f
C35208 _0254_ _0824_/a_59_75# 0
C35209 net58 _0621_/a_285_47# 0
C35210 _0642_/a_215_297# _0086_ 0
C35211 net116 _0350_ 0
C35212 _0109_ _0332_ 0
C35213 _0343_ net40 0.0237f
C35214 _1002_/a_27_47# hold93/a_391_47# 0.00179f
C35215 _1002_/a_193_47# hold93/a_285_47# 0
C35216 hold86/a_49_47# hold86/a_391_47# 0.00188f
C35217 _0662_/a_81_21# _0991_/a_1059_315# 0
C35218 acc0.A\[17\] clknet_1_1__leaf__0461_ 0.06973f
C35219 _1072_/a_1017_47# clknet_0_clk 0
C35220 clknet_1_0__leaf__0458_ _0346_ 0.10629f
C35221 hold67/a_49_47# VPWR 0.30793f
C35222 net239 net209 0
C35223 net207 clknet_1_0__leaf__0457_ 0.0022f
C35224 _0134_ comp0.B\[5\] 0
C35225 _0343_ _1030_/a_634_159# 0.00823f
C35226 net35 _0760_/a_285_47# 0
C35227 _1055_/a_27_47# acc0.A\[9\] 0
C35228 hold31/a_391_47# _0399_ 0
C35229 net202 control0.reset 0
C35230 hold26/a_391_47# _0540_/a_51_297# 0
C35231 _1041_/a_1059_315# _0546_/a_149_47# 0
C35232 net224 net96 0.00508f
C35233 output53/a_27_47# VPWR 0.32818f
C35234 clknet_1_0__leaf__0464_ _1051_/a_381_47# 0
C35235 _1024_/a_975_413# net50 0
C35236 _0958_/a_109_47# _0477_ 0
C35237 _0946_/a_30_53# _0970_/a_27_297# 0
C35238 clknet_1_1__leaf__0463_ control0.reset 0.04016f
C35239 _0163_ _0564_/a_68_297# 0.00155f
C35240 _0350_ _0988_/a_27_47# 0
C35241 net176 _0122_ 0
C35242 hold26/a_285_47# net173 0.00972f
C35243 net25 _0160_ 0
C35244 _0458_ hold28/a_285_47# 0
C35245 _0730_/a_215_47# _0350_ 0
C35246 hold74/a_285_47# VPWR 0.2722f
C35247 _0180_ net154 1.03167f
C35248 _0517_/a_81_21# _0990_/a_891_413# 0
C35249 _0544_/a_51_297# _1043_/a_466_413# 0
C35250 _0369_ _0830_/a_215_47# 0.05375f
C35251 _0646_/a_47_47# _0797_/a_27_413# 0
C35252 _0129_ _0704_/a_68_297# 0
C35253 _0259_ clknet_0__0465_ 0.07999f
C35254 _0762_/a_215_47# clknet_1_0__leaf__0460_ 0
C35255 _0226_ net51 0.00238f
C35256 net140 _1052_/a_27_47# 0
C35257 net58 net222 0.21239f
C35258 _0163_ clknet_1_1__leaf_clk 0.38767f
C35259 net138 net9 0.1588f
C35260 _0176_ _1040_/a_592_47# 0.00353f
C35261 _0715_/a_27_47# _0986_/a_193_47# 0
C35262 _0179_ _1054_/a_381_47# 0
C35263 net125 clkbuf_0__0463_/a_110_47# 0.00702f
C35264 net21 _1044_/a_381_47# 0
C35265 net60 clknet_1_1__leaf__0461_ 0
C35266 _0403_ VPWR 1.05531f
C35267 net8 control0.reset 0.32996f
C35268 _0143_ net137 0
C35269 _0477_ _0160_ 0.39069f
C35270 clknet_1_0__leaf__0458_ _0629_/a_59_75# 0.00331f
C35271 net235 net62 0.01417f
C35272 _0294_ _0371_ 0
C35273 net45 _1018_/a_466_413# 0
C35274 _0357_ hold95/a_391_47# 0
C35275 clknet_1_1__leaf__0461_ net5 0
C35276 _1031_/a_466_413# _0339_ 0.0172f
C35277 net205 _1036_/a_561_413# 0
C35278 hold58/a_49_47# net161 0
C35279 _0973_/a_373_47# _0165_ 0
C35280 net204 _0173_ 0.32926f
C35281 _0997_/a_1059_315# _1013_/a_193_47# 0
C35282 _1024_/a_381_47# _1023_/a_27_47# 0
C35283 _1024_/a_193_47# _1023_/a_891_413# 0
C35284 _0820_/a_510_47# _0369_ 0.00557f
C35285 _0270_ net62 0.10118f
C35286 comp0.B\[13\] _1046_/a_381_47# 0
C35287 net193 _1046_/a_1059_315# 0
C35288 pp[1] pp[4] 0.18239f
C35289 _0180_ _0465_ 0.07038f
C35290 net8 _1061_/a_891_413# 0
C35291 _0084_ _0840_/a_68_297# 0
C35292 _0432_ _0640_/a_215_297# 0.04864f
C35293 _0443_ _0640_/a_109_53# 0.02935f
C35294 _0779_/a_79_21# _0395_ 0.05762f
C35295 _0465_ net218 0.01484f
C35296 _1012_/a_891_413# net98 0
C35297 _1001_/a_27_47# _0350_ 0
C35298 pp[30] _0712_/a_465_47# 0
C35299 _1046_/a_193_47# _1046_/a_381_47# 0.09799f
C35300 _1046_/a_634_159# _1046_/a_891_413# 0.03684f
C35301 _1046_/a_27_47# _1046_/a_561_413# 0.00163f
C35302 _0991_/a_193_47# _0263_ 0.00174f
C35303 hold86/a_391_47# acc0.A\[14\] 0.01077f
C35304 net233 hold100/a_49_47# 0
C35305 net61 hold100/a_391_47# 0.01077f
C35306 net245 acc0.A\[13\] 0
C35307 _1019_/a_891_413# _0772_/a_215_47# 0
C35308 _0130_ _0208_ 0.06568f
C35309 _0413_ _0409_ 0
C35310 clknet_1_0__leaf__0462_ pp[23] 0
C35311 _0391_ _0099_ 0
C35312 pp[26] _0570_/a_27_297# 0
C35313 _0310_ _0395_ 0
C35314 _0949_/a_59_75# clknet_1_0__leaf_clk 0
C35315 net58 _0182_ 0
C35316 acc0.A\[2\] _0180_ 0
C35317 _0174_ _1045_/a_1059_315# 0.00235f
C35318 _1016_/a_891_413# _0115_ 0
C35319 _1032_/a_891_413# clknet_1_0__leaf__0457_ 0.00252f
C35320 control0.state\[0\] VPWR 1.3441f
C35321 _0234_ _0376_ 0.05636f
C35322 _0221_ _0707_/a_208_47# 0
C35323 VPWR _0698_/a_113_297# 0.16368f
C35324 _0403_ _0654_/a_27_413# 0
C35325 acc0.A\[2\] net218 0
C35326 _0753_/a_79_21# _0225_ 0.01378f
C35327 pp[28] _0219_ 0
C35328 hold68/a_49_47# _0122_ 0
C35329 hold68/a_285_47# net110 0.04513f
C35330 _1051_/a_27_47# _1050_/a_634_159# 0.00348f
C35331 _1051_/a_193_47# _1050_/a_193_47# 0
C35332 _1051_/a_634_159# _1050_/a_27_47# 0.00348f
C35333 VPWR _0583_/a_109_297# 0.20737f
C35334 _0285_ _0422_ 0
C35335 _0985_/a_193_47# net175 0
C35336 VPWR net195 0.96933f
C35337 _0218_ _0823_/a_109_297# 0.002f
C35338 _1050_/a_1059_315# _1045_/a_27_47# 0
C35339 pp[8] _0189_ 0
C35340 hold58/a_49_47# net26 0.00516f
C35341 _0186_ _0085_ 0.00618f
C35342 _0984_/a_1059_315# _0346_ 0
C35343 _0996_/a_381_47# acc0.A\[15\] 0.00319f
C35344 clknet_1_0__leaf__0463_ _1038_/a_1059_315# 0
C35345 _0785_/a_81_21# _0181_ 0.02188f
C35346 net196 _0542_/a_512_297# 0.00345f
C35347 hold33/a_285_47# _0172_ 0.03501f
C35348 _0432_ _0465_ 0.08664f
C35349 _0531_/a_27_297# _1049_/a_1059_315# 0
C35350 pp[28] _0728_/a_59_75# 0
C35351 _0343_ _0828_/a_113_297# 0.00763f
C35352 net64 clknet_1_1__leaf__0458_ 0.19394f
C35353 VPWR _0603_/a_150_297# 0.00193f
C35354 _0621_/a_117_297# clknet_1_1__leaf__0458_ 0.00394f
C35355 _0998_/a_634_159# clknet_1_1__leaf__0461_ 0
C35356 _0662_/a_81_21# _0425_ 0
C35357 _0662_/a_384_47# _0290_ 0.00111f
C35358 _0662_/a_299_297# _0401_ 0.02105f
C35359 _0467_ _0175_ 0
C35360 _0214_ _0560_/a_68_297# 0
C35361 _0457_ _1032_/a_466_413# 0.0076f
C35362 clkbuf_0__0461_/a_110_47# net43 0
C35363 net58 _0443_ 0.06302f
C35364 net44 _0999_/a_381_47# 0
C35365 _0245_ _0393_ 0.12403f
C35366 _0336_ hold62/a_49_47# 0.01349f
C35367 _0220_ hold62/a_285_47# 0
C35368 hold76/a_49_47# _0616_/a_78_199# 0
C35369 pp[30] hold16/a_285_47# 0.00937f
C35370 hold54/a_391_47# net23 0
C35371 _1000_/a_891_413# net46 0
C35372 VPWR _0610_/a_59_75# 0.23514f
C35373 VPWR _0999_/a_634_159# 0.20355f
C35374 hold27/a_391_47# _0536_/a_51_297# 0
C35375 clkload3/Y _0998_/a_27_47# 0.00183f
C35376 _0740_/a_113_47# _0324_ 0
C35377 _1052_/a_193_47# acc0.A\[6\] 0.08243f
C35378 net39 _0399_ 0
C35379 net162 _0567_/a_373_47# 0.00188f
C35380 _0100_ clknet_1_0__leaf__0460_ 0.00426f
C35381 net54 hold50/a_391_47# 0
C35382 _0581_/a_27_297# _0581_/a_109_47# 0.00393f
C35383 _0983_/a_193_47# net165 0
C35384 _0229_ acc0.A\[21\] 0.03231f
C35385 _0179_ _0522_/a_27_297# 0.01124f
C35386 acc0.A\[4\] _0638_/a_109_297# 0.00311f
C35387 net233 _0450_ 0
C35388 _0217_ net50 0.84107f
C35389 _0187_ acc0.A\[11\] 0.10575f
C35390 VPWR _0691_/a_68_297# 0.17236f
C35391 _1039_/a_891_413# net8 0.03002f
C35392 _0687_/a_59_75# _0687_/a_145_75# 0.00658f
C35393 hold78/a_391_47# _0195_ 0.00355f
C35394 _0216_ _0728_/a_145_75# 0
C35395 _0985_/a_891_413# _0083_ 0.04505f
C35396 net186 _0474_ 0
C35397 comp0.B\[0\] _0175_ 0.09388f
C35398 net84 _0181_ 0.00212f
C35399 hold85/a_285_47# _0476_ 0.04083f
C35400 _0682_/a_150_297# VPWR 0.00145f
C35401 _0716_/a_27_47# _0287_ 0
C35402 clkbuf_0__0463_/a_110_47# _0473_ 0.03299f
C35403 hold56/a_49_47# _0173_ 0
C35404 _0343_ _0990_/a_634_159# 0.0017f
C35405 _0260_ _0345_ 0
C35406 _0967_/a_109_93# _0970_/a_27_297# 0
C35407 _0970_/a_285_47# _0484_ 0.00113f
C35408 _0970_/a_114_47# _0485_ 0
C35409 _0970_/a_27_297# _0487_ 0.06308f
C35410 _0795_/a_384_47# _0345_ 0
C35411 _0734_/a_285_47# _0326_ 0
C35412 _1053_/a_27_47# _0191_ 0
C35413 _0982_/a_1059_315# _0982_/a_1017_47# 0
C35414 _0982_/a_193_47# net68 0.00242f
C35415 _0982_/a_27_47# _0080_ 0.09142f
C35416 _1049_/a_891_413# _1049_/a_975_413# 0.00851f
C35417 _1049_/a_27_47# net135 0.22945f
C35418 _1049_/a_381_47# _1049_/a_561_413# 0.00123f
C35419 net106 clknet_1_0__leaf__0457_ 0.00978f
C35420 net69 acc0.A\[15\] 0
C35421 _0459_ _0350_ 0.21651f
C35422 clkbuf_0__0464_/a_110_47# _0176_ 0
C35423 net12 acc0.A\[6\] 0.25855f
C35424 net148 net13 0
C35425 net48 _0603_/a_150_297# 0
C35426 _0291_ net47 0
C35427 clknet_1_0__leaf__0465_ _0174_ 0.0015f
C35428 _0172_ net20 0.64973f
C35429 _0483_ control0.state\[2\] 0
C35430 _0747_/a_215_47# _0747_/a_510_47# 0.00529f
C35431 acc0.A\[12\] _0277_ 0.04269f
C35432 _0383_ _0219_ 0.24883f
C35433 _0985_/a_27_47# _0504_/a_27_47# 0
C35434 _0473_ _1044_/a_193_47# 0
C35435 _1070_/a_27_47# _1070_/a_634_159# 0.14145f
C35436 net40 A[14] 0.10018f
C35437 _0399_ _0444_ 0.1212f
C35438 _1053_/a_634_159# _1053_/a_1059_315# 0
C35439 _1053_/a_27_47# _1053_/a_381_47# 0.06222f
C35440 _1053_/a_193_47# _1053_/a_891_413# 0.19685f
C35441 output44/a_27_47# _1030_/a_27_47# 0
C35442 _1057_/a_27_47# acc0.A\[10\] 0.03886f
C35443 net169 input15/a_75_212# 0.00173f
C35444 hold54/a_49_47# clknet_1_0__leaf__0461_ 0.05109f
C35445 net113 acc0.A\[25\] 0.00388f
C35446 clknet_1_0__leaf__0465_ _1050_/a_27_47# 0.00344f
C35447 _0714_/a_149_47# _0218_ 0.01543f
C35448 _0996_/a_634_159# _0181_ 0
C35449 _0129_ _0216_ 0.00267f
C35450 net163 _0195_ 0.00687f
C35451 _0348_ _0128_ 0
C35452 _1066_/a_891_413# _1066_/a_975_413# 0.00851f
C35453 _1066_/a_27_47# clknet_1_1__leaf_clk 0.22327f
C35454 _1066_/a_381_47# _1066_/a_561_413# 0.00123f
C35455 _0627_/a_369_297# acc0.A\[6\] 0
C35456 _1037_/a_193_47# _0176_ 0.00581f
C35457 _0314_ _1007_/a_27_47# 0.00118f
C35458 hold34/a_391_47# A[12] 0.00192f
C35459 _1034_/a_634_159# _0175_ 0
C35460 _0179_ _1056_/a_1017_47# 0.00106f
C35461 net45 net85 0.02608f
C35462 pp[0] B[5] 0
C35463 net31 _1040_/a_1059_315# 0
C35464 _0833_/a_510_47# _0086_ 0
C35465 _0201_ _1042_/a_1059_315# 0
C35466 net177 _1022_/a_27_47# 0
C35467 net109 _1022_/a_193_47# 0.03312f
C35468 hold56/a_391_47# net185 0
C35469 _1068_/a_891_413# _1068_/a_975_413# 0.00851f
C35470 _1068_/a_381_47# _1068_/a_561_413# 0.00123f
C35471 _0222_ hold94/a_391_47# 0.04094f
C35472 clkbuf_1_1__f__0464_/a_110_47# _1044_/a_193_47# 0.01843f
C35473 _1030_/a_634_159# _1030_/a_381_47# 0
C35474 _1041_/a_1059_315# _0176_ 0
C35475 _0712_/a_465_47# _0339_ 0.01141f
C35476 net152 net174 0
C35477 hold74/a_285_47# clknet_1_0__leaf__0459_ 0
C35478 _0322_ _1009_/a_1059_315# 0
C35479 _0402_ net246 0
C35480 _1017_/a_891_413# _0347_ 0
C35481 _0218_ _0116_ 0
C35482 clkbuf_1_1__f__0464_/a_110_47# net131 0.00171f
C35483 _0461_ _0616_/a_292_297# 0
C35484 _0218_ _0807_/a_150_297# 0
C35485 _0639_/a_109_297# _0271_ 0.01129f
C35486 VPWR net111 0.35043f
C35487 A[12] _0510_/a_27_297# 0
C35488 acc0.A\[12\] _0808_/a_81_21# 0
C35489 VPWR _0570_/a_109_297# 0.17646f
C35490 hold100/a_49_47# _0637_/a_311_297# 0
C35491 net146 _0347_ 0
C35492 _0221_ acc0.A\[30\] 0
C35493 _0258_ _0845_/a_109_47# 0
C35494 _1035_/a_975_413# clknet_1_1__leaf__0463_ 0
C35495 _1035_/a_381_47# net122 0
C35496 _0753_/a_561_47# net46 0.00126f
C35497 hold77/a_49_47# clkbuf_1_1__f__0460_/a_110_47# 0
C35498 _0992_/a_1059_315# net37 0.12233f
C35499 _0343_ _0433_ 0
C35500 control0.count\[1\] control0.state\[2\] 0.0015f
C35501 _0804_/a_510_47# _0347_ 0.00524f
C35502 _0346_ hold91/a_285_47# 0.04442f
C35503 _0786_/a_217_297# _0401_ 0.01578f
C35504 _0786_/a_472_297# _0290_ 0
C35505 hold18/a_49_47# _0346_ 0
C35506 _0201_ net10 0
C35507 net122 input23/a_75_212# 0.00178f
C35508 _0123_ net200 0
C35509 _0679_/a_68_297# _0746_/a_81_21# 0
C35510 _0598_/a_297_47# _0229_ 0.00638f
C35511 _0598_/a_79_21# _0226_ 0.00163f
C35512 _1015_/a_381_47# _0181_ 0
C35513 _0320_ _0737_/a_285_297# 0
C35514 VPWR _0517_/a_299_297# 0.20635f
C35515 _0987_/a_27_47# _0987_/a_891_413# 0.03224f
C35516 _0987_/a_193_47# _0987_/a_1059_315# 0.03405f
C35517 _0987_/a_634_159# _0987_/a_466_413# 0.23992f
C35518 clknet_0__0459_ _0507_/a_109_297# 0
C35519 _0236_ _0218_ 0
C35520 _0183_ net102 0.01047f
C35521 _0152_ _0252_ 0.00425f
C35522 acc0.A\[1\] _0261_ 0
C35523 _0182_ _0262_ 0
C35524 net248 _0437_ 0.00152f
C35525 net194 _1051_/a_193_47# 0.00467f
C35526 _0579_/a_109_297# _0217_ 0.01309f
C35527 output42/a_27_47# net81 0.00776f
C35528 _0695_/a_80_21# _0315_ 0
C35529 _0265_ _0350_ 0.01202f
C35530 _1021_/a_193_47# net106 0
C35531 hold49/a_285_47# _1044_/a_27_47# 0
C35532 _1034_/a_1017_47# comp0.B\[2\] 0
C35533 net168 acc0.A\[5\] 0
C35534 net194 _1045_/a_466_413# 0
C35535 output64/a_27_47# _0833_/a_79_21# 0
C35536 clknet_0__0465_ _0253_ 0
C35537 clknet_0__0459_ hold82/a_49_47# 0
C35538 acc0.A\[27\] _1008_/a_592_47# 0.00112f
C35539 net131 _0186_ 0
C35540 _0992_/a_381_47# net67 0
C35541 clknet_1_0__leaf__0465_ _0518_/a_27_297# 0.00238f
C35542 _0342_ clknet_1_1__leaf__0462_ 0
C35543 hold43/a_285_47# acc0.A\[27\] 0
C35544 _1000_/a_381_47# VPWR 0.07663f
C35545 _1004_/a_27_47# _1004_/a_634_159# 0.14145f
C35546 _0225_ clkbuf_1_0__f__0460_/a_110_47# 0.00149f
C35547 hold16/a_285_47# _0339_ 0.02006f
C35548 _0169_ _0488_ 0.09498f
C35549 clkbuf_0__0464_/a_110_47# net130 0
C35550 _0151_ _1053_/a_466_413# 0
C35551 _0217_ _0399_ 0.07109f
C35552 _0486_ clkbuf_1_0__f_clk/a_110_47# 0
C35553 acc0.A\[14\] net228 0
C35554 _0182_ net23 0
C35555 pp[27] hold61/a_285_47# 0.00675f
C35556 _0476_ _0958_/a_27_47# 0.12267f
C35557 _0718_/a_377_297# net56 0
C35558 input34/a_27_47# _1064_/a_27_47# 0
C35559 _0225_ _0250_ 0.00432f
C35560 net85 _0587_/a_27_47# 0
C35561 _0608_/a_27_47# _0219_ 0.00697f
C35562 hold77/a_391_47# net96 0
C35563 net9 hold83/a_285_47# 0
C35564 _0346_ _0288_ 0.06271f
C35565 net58 _0089_ 0
C35566 _1029_/a_634_159# _1029_/a_466_413# 0.23992f
C35567 _1029_/a_193_47# _1029_/a_1059_315# 0.03405f
C35568 _1029_/a_27_47# _1029_/a_891_413# 0.03224f
C35569 VPWR hold50/a_285_47# 0.29435f
C35570 clknet_1_0__leaf__0459_ _0583_/a_109_297# 0.00529f
C35571 _0629_/a_59_75# hold18/a_49_47# 0
C35572 _0334_ clknet_1_1__leaf__0462_ 0
C35573 hold21/a_285_47# _0186_ 0
C35574 _0482_ hold79/a_391_47# 0
C35575 _0964_/a_109_297# net226 0.00112f
C35576 _0856_/a_297_297# _0346_ 0.00874f
C35577 VPWR _0565_/a_51_297# 0.53714f
C35578 _1001_/a_27_47# _0244_ 0
C35579 _1032_/a_1017_47# clknet_1_0__leaf__0461_ 0
C35580 _0318_ _0360_ 0
C35581 net39 _0299_ 0
C35582 acc0.A\[12\] _0298_ 0.11136f
C35583 A[12] _0181_ 0.0763f
C35584 net61 _0256_ 0.28306f
C35585 net136 _0270_ 0
C35586 _0637_/a_311_297# _0450_ 0
C35587 _0274_ acc0.A\[6\] 0.02992f
C35588 _0343_ _0998_/a_975_413# 0
C35589 _0290_ net47 0
C35590 hold65/a_285_47# VPWR 0.27149f
C35591 _0430_ _0831_/a_285_297# 0.00574f
C35592 comp0.B\[13\] _1045_/a_1059_315# 0.1364f
C35593 _1050_/a_466_413# net73 0
C35594 net136 _0987_/a_466_413# 0
C35595 _0767_/a_59_75# _0294_ 0.0896f
C35596 _0961_/a_113_297# _0961_/a_199_47# 0
C35597 _0369_ acc0.A\[23\] 0
C35598 _1015_/a_193_47# _0565_/a_512_297# 0
C35599 hold97/a_285_47# _0345_ 0.1032f
C35600 acc0.A\[12\] _0296_ 0.10859f
C35601 _1046_/a_891_413# _1045_/a_27_47# 0
C35602 acc0.A\[1\] _0509_/a_27_47# 0.00127f
C35603 _1017_/a_891_413# _1016_/a_891_413# 0
C35604 _1003_/a_1059_315# _0596_/a_59_75# 0
C35605 _0661_/a_27_297# _0292_ 0.05899f
C35606 _0186_ hold71/a_49_47# 0
C35607 _0760_/a_47_47# net51 0
C35608 _0346_ _0247_ 0
C35609 A[10] _0514_/a_27_297# 0
C35610 net187 acc0.A\[20\] 0.73693f
C35611 _1037_/a_891_413# clknet_1_1__leaf__0463_ 0
C35612 net229 _0219_ 0
C35613 clkbuf_1_0__f__0457_/a_110_47# _0346_ 0.01809f
C35614 _1033_/a_466_413# _0956_/a_32_297# 0
C35615 hold96/a_285_47# acc0.A\[23\] 0
C35616 _0960_/a_27_47# _0976_/a_505_21# 0.03113f
C35617 _1028_/a_27_47# _1028_/a_1059_315# 0.04819f
C35618 _1028_/a_193_47# _1028_/a_466_413# 0.07482f
C35619 _0555_/a_149_47# _0555_/a_240_47# 0.06872f
C35620 _0180_ clknet_0__0464_ 0
C35621 hold41/a_391_47# _1057_/a_634_159# 0
C35622 hold41/a_285_47# _1057_/a_466_413# 0
C35623 _0361_ VPWR 0.3592f
C35624 _0465_ _0495_/a_150_297# 0
C35625 net216 _0359_ 0
C35626 _0620_/a_113_47# _0369_ 0
C35627 _0369_ _0989_/a_27_47# 0.00443f
C35628 _0398_ net42 0
C35629 _0924_/a_27_47# clknet_1_1__leaf__0457_ 0.22202f
C35630 _0195_ hold60/a_285_47# 0.03347f
C35631 _0111_ _0220_ 0
C35632 _0999_/a_27_47# _0783_/a_215_47# 0
C35633 _0999_/a_193_47# _0783_/a_297_297# 0
C35634 _0476_ _0132_ 0.25225f
C35635 _0306_ _1009_/a_1059_315# 0
C35636 _0394_ _1009_/a_634_159# 0
C35637 _1033_/a_634_159# comp0.B\[1\] 0
C35638 _1033_/a_891_413# _0131_ 0
C35639 _0369_ _0992_/a_27_47# 0.00832f
C35640 _0985_/a_1059_315# VPWR 0.38668f
C35641 net63 _0987_/a_381_47# 0
C35642 VPWR _1018_/a_466_413# 0.24305f
C35643 input5/a_75_212# pp[14] 0
C35644 _0343_ pp[17] 0
C35645 _0344_ acc0.A\[30\] 0
C35646 _0521_/a_81_21# clknet_1_0__leaf__0465_ 0.00254f
C35647 VPWR _1049_/a_193_47# 0.29722f
C35648 hold55/a_49_47# _0130_ 0.28755f
C35649 _0743_/a_245_297# _0367_ 0.00126f
C35650 clkbuf_0__0463_/a_110_47# _0497_/a_68_297# 0.01186f
C35651 VPWR _0552_/a_68_297# 0.16412f
C35652 net88 hold93/a_49_47# 0
C35653 acc0.A\[1\] net47 0.59762f
C35654 net105 net149 0
C35655 _1009_/a_592_47# _0219_ 0.00169f
C35656 _0482_ _0481_ 0.10024f
C35657 VPWR _1066_/a_193_47# 0.35762f
C35658 _1050_/a_1017_47# acc0.A\[4\] 0.00168f
C35659 net15 _0987_/a_561_413# 0
C35660 _0421_ net37 0
C35661 net242 _0334_ 0.00441f
C35662 net180 clknet_1_1__leaf__0457_ 0.00211f
C35663 VPWR _1068_/a_193_47# 0.28051f
C35664 VPWR input1/a_27_47# 0.26939f
C35665 pp[28] hold61/a_49_47# 0
C35666 _0991_/a_27_47# _0267_ 0
C35667 _1041_/a_891_413# _0139_ 0
C35668 _1041_/a_975_413# net32 0
C35669 clknet_1_0__leaf__0464_ acc0.A\[5\] 0
C35670 _0455_ _0346_ 0.03543f
C35671 _0366_ _0345_ 0
C35672 _0257_ hold101/a_391_47# 0.00283f
C35673 _0258_ hold101/a_49_47# 0
C35674 _0626_/a_68_297# net248 0
C35675 _0277_ net42 0.02822f
C35676 clkbuf_1_1__f__0459_/a_110_47# net5 0
C35677 _0300_ acc0.A\[15\] 0
C35678 _0244_ _0459_ 0.04019f
C35679 _0230_ _0606_/a_109_53# 0
C35680 _0993_/a_193_47# _0417_ 0
C35681 _0993_/a_891_413# net79 0
C35682 VPWR _0204_ 0.22314f
C35683 clknet_0__0457_ hold60/a_49_47# 0
C35684 _0983_/a_891_413# _1018_/a_1059_315# 0
C35685 net243 net52 0
C35686 comp0.B\[13\] clknet_1_0__leaf__0465_ 0
C35687 VPWR _1034_/a_975_413# 0.00418f
C35688 net45 _0587_/a_27_47# 0.01568f
C35689 _0187_ _0281_ 0
C35690 hold66/a_285_47# _0228_ 0.02259f
C35691 hold42/a_391_47# _0179_ 0.05624f
C35692 hold32/a_49_47# input16/a_75_212# 0
C35693 _0179_ _1057_/a_891_413# 0
C35694 _0544_/a_51_297# net196 0
C35695 net198 _1043_/a_891_413# 0.00929f
C35696 _0140_ _1043_/a_193_47# 0.00173f
C35697 _0478_ VPWR 0.57706f
C35698 _1004_/a_193_47# net199 0
C35699 hold34/a_391_47# _0154_ 0.0021f
C35700 _0107_ _0680_/a_80_21# 0
C35701 VPWR hold6/a_391_47# 0.18362f
C35702 clknet_1_0__leaf__0464_ _0528_/a_299_297# 0.01733f
C35703 clknet_1_0__leaf__0465_ _1046_/a_193_47# 0.00705f
C35704 net103 net219 0.00177f
C35705 _0642_/a_27_413# acc0.A\[8\] 0.02098f
C35706 _0697_/a_80_21# _0689_/a_68_297# 0
C35707 _0343_ _0983_/a_1059_315# 0.02921f
C35708 _0531_/a_27_297# net175 0.05897f
C35709 _1057_/a_193_47# _0181_ 0
C35710 _0170_ _1071_/a_27_47# 0
C35711 _0578_/a_109_297# _0460_ 0
C35712 _0578_/a_373_47# clknet_1_0__leaf__0457_ 0
C35713 clknet_0__0458_ _0219_ 0
C35714 _1028_/a_27_47# _0347_ 0.00127f
C35715 hold19/a_285_47# hold72/a_285_47# 0
C35716 acc0.A\[0\] hold2/a_285_47# 0.00906f
C35717 net63 acc0.A\[4\] 0
C35718 acc0.A\[14\] _1016_/a_1059_315# 0
C35719 _1019_/a_27_47# clkbuf_0__0457_/a_110_47# 0.02974f
C35720 _1002_/a_891_413# acc0.A\[20\] 0
C35721 _0998_/a_1059_315# _0998_/a_891_413# 0.31086f
C35722 _0998_/a_193_47# _0998_/a_975_413# 0
C35723 _0998_/a_466_413# _0998_/a_381_47# 0.03733f
C35724 _0551_/a_27_47# _0499_/a_59_75# 0
C35725 _0579_/a_27_297# hold40/a_49_47# 0
C35726 net64 _0988_/a_1017_47# 0.0017f
C35727 _0529_/a_109_297# _0186_ 0.02064f
C35728 _0498_/a_51_297# _0465_ 0.00173f
C35729 _0779_/a_297_297# _0306_ 0
C35730 _0779_/a_215_47# _0308_ 0
C35731 hold10/a_49_47# net247 0
C35732 _1003_/a_891_413# _0369_ 0
C35733 _0267_ _0350_ 0.02866f
C35734 _1024_/a_27_47# acc0.A\[23\] 0.00114f
C35735 net110 _1023_/a_1059_315# 0.00161f
C35736 _0259_ _0986_/a_27_47# 0
C35737 _0386_ clknet_1_0__leaf__0461_ 0
C35738 hold38/a_49_47# comp0.B\[3\] 0.31185f
C35739 _0432_ _0254_ 0.19102f
C35740 _0350_ _0772_/a_79_21# 0.00139f
C35741 VPWR acc0.A\[13\] 1.31622f
C35742 comp0.B\[15\] _0145_ 0.00141f
C35743 _1019_/a_193_47# _1019_/a_381_47# 0.09541f
C35744 _1019_/a_634_159# _1019_/a_891_413# 0.03684f
C35745 _1019_/a_27_47# _1019_/a_561_413# 0.00163f
C35746 _0717_/a_209_47# _0221_ 0
C35747 net44 _1012_/a_975_413# 0
C35748 hold76/a_285_47# _0216_ 0
C35749 _0143_ _0148_ 0
C35750 _1057_/a_27_47# _0188_ 0
C35751 _0837_/a_585_47# _0172_ 0.00114f
C35752 clknet_1_0__leaf__0464_ _0182_ 0
C35753 net72 _0986_/a_193_47# 0.00124f
C35754 clknet_1_1__leaf__0458_ _0986_/a_466_413# 0
C35755 VPWR _1012_/a_1059_315# 0.41387f
C35756 hold54/a_285_47# _0173_ 0
C35757 _0565_/a_149_47# _0215_ 0.00154f
C35758 hold52/a_391_47# _1024_/a_891_413# 0.00274f
C35759 _0548_/a_149_47# _1040_/a_891_413# 0
C35760 _0548_/a_240_47# _1040_/a_1059_315# 0
C35761 _1050_/a_193_47# net184 0
C35762 _1050_/a_634_159# net131 0
C35763 comp0.B\[15\] net17 0.00112f
C35764 output59/a_27_47# clknet_1_1__leaf__0462_ 0.03031f
C35765 _0331_ _0332_ 0.05213f
C35766 _1058_/a_27_47# net67 0.02747f
C35767 net123 net124 0
C35768 _1033_/a_1059_315# _1032_/a_27_47# 0.00468f
C35769 _1033_/a_27_47# _1032_/a_1059_315# 0.00468f
C35770 _1063_/a_27_47# _0468_ 0
C35771 _0211_ comp0.B\[4\] 0.05354f
C35772 net196 _0141_ 0.29847f
C35773 net175 _1049_/a_592_47# 0
C35774 _0389_ _0343_ 0.00206f
C35775 hold8/a_285_47# acc0.A\[25\] 0.0018f
C35776 pp[6] net62 0
C35777 _0786_/a_80_21# hold70/a_285_47# 0.00114f
C35778 B[12] net32 0.00296f
C35779 net84 clknet_1_1__leaf__0461_ 0.03102f
C35780 _0694_/a_113_47# _0324_ 0
C35781 _0287_ _0426_ 0
C35782 _0503_/a_109_297# control0.sh 0
C35783 hold25/a_49_47# _1039_/a_27_47# 0
C35784 hold32/a_285_47# pp[4] 0
C35785 acc0.A\[8\] _0218_ 0
C35786 net1 _0526_/a_27_47# 0.03472f
C35787 _0718_/a_47_47# hold16/a_285_47# 0
C35788 acc0.A\[31\] _1031_/a_1059_315# 0.08415f
C35789 _0502_/a_27_47# acc0.A\[15\] 0.04961f
C35790 net162 _1031_/a_634_159# 0.01053f
C35791 _0457_ net202 0.04456f
C35792 _0974_/a_448_47# _0468_ 0.0017f
C35793 _0342_ hold92/a_49_47# 0
C35794 clknet_1_0__leaf__0465_ _0987_/a_27_47# 0.01588f
C35795 hold99/a_391_47# net79 0
C35796 _0457_ clknet_1_1__leaf__0463_ 0.05227f
C35797 _1021_/a_1059_315# _0578_/a_27_297# 0
C35798 net101 _0183_ 0
C35799 _0294_ net166 0
C35800 net81 _0799_/a_80_21# 0
C35801 _0758_/a_215_47# _0347_ 0.05741f
C35802 _1024_/a_1059_315# pp[24] 0
C35803 _1024_/a_381_47# net52 0
C35804 VPWR net85 0.44503f
C35805 _0236_ _0099_ 0
C35806 _0154_ _0181_ 0
C35807 clknet_0__0458_ _0826_/a_301_297# 0
C35808 _0991_/a_193_47# _0218_ 0
C35809 _0294_ _0991_/a_634_159# 0.00833f
C35810 _0375_ VPWR 0.37087f
C35811 _0984_/a_1017_47# _0465_ 0
C35812 _0246_ _0352_ 0.03135f
C35813 _0350_ net51 0.3228f
C35814 _0990_/a_634_159# _0990_/a_381_47# 0
C35815 _0343_ _0355_ 0.00118f
C35816 _0404_ acc0.A\[15\] 0
C35817 hold81/a_49_47# _0806_/a_199_47# 0
C35818 _0790_/a_285_47# _0345_ 0
C35819 _0179_ _0193_ 0.03781f
C35820 _1002_/a_27_47# _0460_ 0.04892f
C35821 _1002_/a_634_159# clknet_1_0__leaf__0457_ 0.00187f
C35822 _0571_/a_27_297# hold8/a_285_47# 0.00152f
C35823 _0984_/a_592_47# net58 0
C35824 _0747_/a_510_47# _0352_ 0.00378f
C35825 _0174_ _0546_/a_240_47# 0.02494f
C35826 _0362_ _0350_ 0.11299f
C35827 _0296_ net42 0
C35828 hold86/a_49_47# _0268_ 0
C35829 _0183_ _0228_ 0
C35830 _0967_/a_109_93# _0967_/a_487_297# 0
C35831 _0967_/a_215_297# _0967_/a_403_297# 0.00122f
C35832 _0346_ _1014_/a_592_47# 0
C35833 acc0.A\[25\] _1007_/a_891_413# 0
C35834 _0695_/a_217_297# acc0.A\[24\] 0
C35835 hold97/a_391_47# _0329_ 0
C35836 output44/a_27_47# net44 0.17968f
C35837 clkbuf_1_0__f__0465_/a_110_47# _0271_ 0
C35838 clknet_1_0__leaf__0465_ comp0.B\[9\] 0
C35839 output58/a_27_47# pp[2] 0.33656f
C35840 net44 clknet_1_1__leaf__0459_ 0.00388f
C35841 clknet_1_1__leaf__0463_ _1062_/a_891_413# 0
C35842 hold53/a_49_47# _1025_/a_1059_315# 0.00791f
C35843 hold53/a_391_47# _1025_/a_634_159# 0
C35844 _0802_/a_59_75# clknet_1_1__leaf__0459_ 0
C35845 _1049_/a_1017_47# _0147_ 0.00125f
C35846 _1049_/a_561_413# acc0.A\[3\] 0
C35847 net155 clknet_1_1__leaf__0462_ 0.00206f
C35848 _0302_ _0301_ 0
C35849 clknet_1_0__leaf__0459_ _1018_/a_466_413# 0
C35850 _0230_ hold3/a_285_47# 0
C35851 _0226_ hold3/a_391_47# 0
C35852 net248 _0252_ 0
C35853 net243 _0576_/a_109_47# 0
C35854 _0606_/a_109_53# _0236_ 0.11195f
C35855 _0257_ _0369_ 0.00155f
C35856 _0645_/a_47_47# _0399_ 0
C35857 _1045_/a_27_47# _1045_/a_466_413# 0.27314f
C35858 _1045_/a_193_47# _1045_/a_634_159# 0.12729f
C35859 _1070_/a_891_413# _1070_/a_975_413# 0.00851f
C35860 _1070_/a_193_47# VPWR 0.32759f
C35861 _1070_/a_381_47# _1070_/a_561_413# 0.00123f
C35862 _1052_/a_381_47# _0150_ 0.12823f
C35863 _0255_ net75 0
C35864 pp[17] _1030_/a_381_47# 0
C35865 net44 _1030_/a_975_413# 0
C35866 net245 VPWR 0.26302f
C35867 _1015_/a_975_413# net118 0
C35868 control0.reset _0492_/a_27_47# 0.00165f
C35869 _0689_/a_68_297# _0345_ 0.02598f
C35870 net45 _0998_/a_1017_47# 0
C35871 hold26/a_49_47# clknet_0__0463_ 0
C35872 _1014_/a_1059_315# _0465_ 0.00114f
C35873 _1062_/a_1059_315# _0468_ 0
C35874 net203 net17 0
C35875 VPWR _1030_/a_1059_315# 0.37857f
C35876 _0683_/a_113_47# _0105_ 0
C35877 net77 net47 0.13277f
C35878 _0378_ _0345_ 0
C35879 _1043_/a_27_47# _1043_/a_466_413# 0.27314f
C35880 _1043_/a_193_47# _1043_/a_634_159# 0.11072f
C35881 net7 _1040_/a_1059_315# 0
C35882 net234 net104 0
C35883 _0502_/a_27_47# _0179_ 0.00342f
C35884 _0309_ _0395_ 0.0027f
C35885 _1017_/a_466_413# hold72/a_49_47# 0
C35886 _0749_/a_81_21# _0219_ 0
C35887 B[12] net10 0
C35888 _0997_/a_381_47# net83 0.00161f
C35889 _0366_ net52 0.00371f
C35890 _1038_/a_634_159# _0209_ 0.00124f
C35891 _0678_/a_68_297# _0219_ 0.00963f
C35892 net236 _0975_/a_145_75# 0
C35893 clknet_1_1__leaf__0463_ _0475_ 0
C35894 net103 _0352_ 0
C35895 control0.state\[0\] comp0.B\[3\] 0
C35896 hold67/a_391_47# _0399_ 0
C35897 net46 net104 0
C35898 _1021_/a_466_413# _1002_/a_27_47# 0
C35899 _1021_/a_27_47# _1002_/a_466_413# 0.00138f
C35900 _1021_/a_634_159# _1002_/a_193_47# 0.01021f
C35901 _1021_/a_193_47# _1002_/a_634_159# 0
C35902 _1004_/a_193_47# VPWR 0.31772f
C35903 net242 _0724_/a_113_297# 0
C35904 clknet_1_0__leaf__0458_ _1047_/a_466_413# 0
C35905 _0785_/a_299_297# _0990_/a_27_47# 0
C35906 VPWR _0493_/a_27_47# 0.00145f
C35907 A[12] _0187_ 0
C35908 acc0.A\[14\] _0268_ 0.07562f
C35909 hold100/a_391_47# _0269_ 0
C35910 net182 _0517_/a_299_297# 0
C35911 _0125_ net113 0
C35912 _0645_/a_377_297# _0277_ 0.00272f
C35913 _1056_/a_634_159# _1056_/a_381_47# 0
C35914 _1032_/a_561_413# net17 0
C35915 _0671_/a_199_47# _0303_ 0.00181f
C35916 hold28/a_49_47# _0182_ 0
C35917 comp0.B\[10\] _1042_/a_27_47# 0
C35918 _0423_ _0218_ 0
C35919 _0294_ _0290_ 0.17132f
C35920 _0256_ _0431_ 0
C35921 pp[27] _0730_/a_79_21# 0
C35922 net194 _1044_/a_634_159# 0
C35923 _0987_/a_634_159# _0085_ 0.04557f
C35924 _0987_/a_466_413# net73 0
C35925 _0476_ net25 0.03424f
C35926 _0282_ _0806_/a_113_297# 0
C35927 input11/a_75_212# A[5] 0.03292f
C35928 A[4] input12/a_75_212# 0.00451f
C35929 _0245_ _0773_/a_35_297# 0.02339f
C35930 _0315_ clknet_1_0__leaf__0460_ 0.00427f
C35931 _0335_ _0703_/a_109_297# 0.01294f
C35932 hold87/a_391_47# _0241_ 0
C35933 _0327_ _0367_ 0.00371f
C35934 _0833_/a_215_47# acc0.A\[8\] 0.00542f
C35935 _1007_/a_27_47# _0360_ 0
C35936 _0855_/a_81_21# _0456_ 0.12757f
C35937 _0799_/a_80_21# _0797_/a_207_413# 0.00121f
C35938 acc0.A\[1\] _1047_/a_1017_47# 0
C35939 _0199_ _1047_/a_891_413# 0
C35940 _0182_ _1047_/a_592_47# 0.00129f
C35941 net194 net184 0
C35942 net162 _0345_ 0
C35943 _0145_ hold71/a_285_47# 0
C35944 net54 pp[26] 0.01118f
C35945 net71 clknet_1_1__leaf__0457_ 0.00112f
C35946 clknet_1_0__leaf__0465_ _0191_ 0.00136f
C35947 _1004_/a_381_47# _1004_/a_561_413# 0.00123f
C35948 _1004_/a_891_413# _1004_/a_975_413# 0.00851f
C35949 net45 VPWR 2.3717f
C35950 net47 _0986_/a_1059_315# 0.00348f
C35951 clknet_1_0__leaf__0459_ acc0.A\[13\] 0.10956f
C35952 _1027_/a_466_413# _1008_/a_891_413# 0
C35953 _1027_/a_891_413# _1008_/a_466_413# 0
C35954 acc0.A\[31\] _0712_/a_561_47# 0
C35955 net162 _0712_/a_381_47# 0
C35956 net170 _0186_ 0.23445f
C35957 pp[8] net67 0
C35958 _1067_/a_466_413# hold93/a_391_47# 0
C35959 _0983_/a_27_47# _0983_/a_193_47# 0.96544f
C35960 _0476_ _0477_ 0.08255f
C35961 _0181_ acc0.A\[18\] 0
C35962 _0735_/a_109_297# clknet_1_1__leaf__0460_ 0
C35963 hold69/a_49_47# clknet_0__0460_ 0
C35964 _1029_/a_634_159# net191 0
C35965 acc0.A\[16\] net221 0.50435f
C35966 _0301_ net6 0
C35967 _1019_/a_1059_315# _0352_ 0
C35968 _0625_/a_145_75# acc0.A\[5\] 0
C35969 B[1] B[5] 0.42071f
C35970 net150 clknet_1_0__leaf__0460_ 0.0399f
C35971 _0244_ _0772_/a_79_21# 0
C35972 VPWR _0531_/a_373_47# 0
C35973 _0535_/a_150_297# _0176_ 0
C35974 clknet_1_0__leaf__0462_ _0574_/a_27_297# 0.02767f
C35975 acc0.A\[24\] _0345_ 0
C35976 clknet_1_0__leaf__0458_ _0782_/a_27_47# 0
C35977 acc0.A\[4\] _0987_/a_1017_47# 0
C35978 _0514_/a_109_297# net143 0
C35979 _1000_/a_466_413# acc0.A\[18\] 0
C35980 _0113_ _0565_/a_51_297# 0
C35981 hold47/a_285_47# _0180_ 0.0086f
C35982 _1020_/a_466_413# _0183_ 0.019f
C35983 _1020_/a_891_413# _0217_ 0
C35984 net216 _0325_ 0
C35985 net103 _1016_/a_975_413# 0
C35986 net162 hold16/a_49_47# 0.13713f
C35987 hold15/a_391_47# _0129_ 0.01869f
C35988 _0289_ _0287_ 0.51647f
C35989 _0292_ _0293_ 0.00234f
C35990 _0210_ comp0.B\[4\] 0.0076f
C35991 _1016_/a_634_159# _1016_/a_1059_315# 0
C35992 _1016_/a_27_47# _1016_/a_381_47# 0.05761f
C35993 _1016_/a_193_47# _1016_/a_891_413# 0.19226f
C35994 _0172_ B[9] 0
C35995 _0854_/a_79_21# clknet_1_0__leaf__0461_ 0.01458f
C35996 A[10] _0189_ 0.05117f
C35997 hold101/a_391_47# clknet_1_1__leaf__0458_ 0
C35998 hold57/a_49_47# control0.reset 0
C35999 hold13/a_49_47# _0176_ 0
C36000 VPWR _0726_/a_51_297# 0.52474f
C36001 net60 _0567_/a_27_297# 0
C36002 _0429_ _0369_ 0.00452f
C36003 output59/a_27_47# hold92/a_49_47# 0.02157f
C36004 hold11/a_391_47# _1061_/a_634_159# 0
C36005 hold11/a_285_47# _1061_/a_466_413# 0
C36006 hold11/a_49_47# _1061_/a_1059_315# 0
C36007 acc0.A\[11\] clknet_1_1__leaf__0465_ 0.02153f
C36008 VPWR _0587_/a_27_47# 0.43165f
C36009 _0566_/a_27_47# _0171_ 0
C36010 _0131_ _0956_/a_32_297# 0.00282f
C36011 _0960_/a_27_47# _0466_ 0
C36012 _0960_/a_109_47# _0488_ 0.00144f
C36013 _1028_/a_634_159# net114 0
C36014 _1028_/a_891_413# _1028_/a_1017_47# 0.00617f
C36015 hold25/a_285_47# _1041_/a_634_159# 0
C36016 hold89/a_285_47# _0477_ 0
C36017 hold41/a_285_47# net189 0.00329f
C36018 hold17/a_285_47# _1070_/a_193_47# 0
C36019 hold17/a_391_47# _1070_/a_27_47# 0
C36020 _0343_ _0996_/a_975_413# 0
C36021 hold87/a_391_47# _0982_/a_193_47# 0
C36022 _0232_ _0460_ 0
C36023 _0723_/a_27_413# _0723_/a_207_413# 0.18542f
C36024 hold42/a_49_47# net4 0.00442f
C36025 _1067_/a_466_413# control0.reset 0
C36026 _1057_/a_193_47# _0187_ 0.01912f
C36027 _1057_/a_466_413# net4 0
C36028 _0442_ _0255_ 0.02461f
C36029 _0303_ clkbuf_1_1__f__0459_/a_110_47# 0.00871f
C36030 _0462_ clkbuf_1_0__f__0460_/a_110_47# 0
C36031 clkbuf_0__0462_/a_110_47# clknet_0__0460_ 0
C36032 _0736_/a_311_297# _0361_ 0
C36033 VPWR _0990_/a_1059_315# 0.42957f
C36034 _0812_/a_79_21# net217 0.05853f
C36035 net220 clknet_1_0__leaf__0457_ 0.00205f
C36036 _0542_/a_51_297# hold51/a_285_47# 0.00175f
C36037 _0999_/a_466_413# _0096_ 0
C36038 net85 _0783_/a_79_21# 0
C36039 hold57/a_391_47# net171 0
C36040 hold57/a_285_47# _0207_ 0
C36041 _0514_/a_27_297# _0514_/a_373_47# 0.01338f
C36042 _0462_ _0250_ 0.00295f
C36043 _0557_/a_149_47# _1037_/a_1059_315# 0
C36044 _0584_/a_27_297# _0584_/a_109_47# 0.00393f
C36045 _0195_ net116 0
C36046 _0179_ net16 0.01156f
C36047 _0472_ _0560_/a_68_297# 0.01458f
C36048 net219 _0774_/a_68_297# 0.05089f
C36049 _0238_ net216 0
C36050 hold59/a_49_47# _0181_ 0
C36051 _0788_/a_68_297# _0417_ 0
C36052 hold4/a_49_47# _1022_/a_27_47# 0.01435f
C36053 _0422_ net228 0.20196f
C36054 _0800_/a_51_297# net5 0
C36055 _1017_/a_466_413# clknet_0__0461_ 0
C36056 _0460_ _1006_/a_561_413# 0
C36057 net199 VPWR 0.44765f
C36058 _0186_ _0525_/a_81_21# 0.00389f
C36059 net21 clknet_1_1__leaf__0464_ 0.23091f
C36060 _0532_/a_81_21# _1047_/a_1059_315# 0
C36061 comp0.B\[1\] clkbuf_0__0457_/a_110_47# 0
C36062 net120 _0474_ 0
C36063 net167 _0480_ 0
C36064 net53 _0743_/a_51_297# 0
C36065 clknet_1_0__leaf__0462_ _0757_/a_150_297# 0
C36066 _0170_ _1072_/a_634_159# 0
C36067 _0370_ _0359_ 0.3894f
C36068 hold57/a_391_47# net24 0
C36069 _0562_/a_68_297# _0173_ 0.01939f
C36070 net34 _0466_ 0.07048f
C36071 net81 _0997_/a_1059_315# 0.00124f
C36072 net61 clknet_0__0465_ 0
C36073 clknet_1_0__leaf__0462_ _0326_ 0
C36074 clkload0/X _0217_ 0
C36075 _0305_ _0776_/a_109_297# 0
C36076 _0357_ net97 0.00193f
C36077 net236 _0960_/a_27_47# 0
C36078 net137 _0987_/a_27_47# 0
C36079 _1051_/a_27_47# net73 0
C36080 clknet_1_0__leaf__0462_ _1025_/a_634_159# 0.00356f
C36081 _1056_/a_1059_315# VPWR 0.39673f
C36082 clkbuf_1_0__f__0459_/a_110_47# _0983_/a_1059_315# 0
C36083 clknet_1_1__leaf__0459_ _0655_/a_369_297# 0
C36084 net15 acc0.A\[8\] 0
C36085 hold87/a_391_47# _0450_ 0
C36086 clknet_1_1__leaf__0463_ net27 0.03424f
C36087 acc0.A\[12\] _0652_/a_109_297# 0
C36088 _1041_/a_193_47# input7/a_75_212# 0
C36089 clknet_1_0__leaf__0460_ control0.add 0.13729f
C36090 _0388_ _0294_ 0.01987f
C36091 _0386_ _0218_ 0
C36092 _0742_/a_81_21# clknet_1_0__leaf__0460_ 0.00207f
C36093 _0695_/a_300_47# _0368_ 0
C36094 _1018_/a_27_47# acc0.A\[18\] 0.04661f
C36095 _0217_ _0576_/a_27_297# 0.16956f
C36096 _1028_/a_27_47# _0106_ 0
C36097 _0271_ _0824_/a_145_75# 0.00146f
C36098 _0387_ _0245_ 0.0016f
C36099 hold57/a_285_47# _1039_/a_1059_315# 0
C36100 clknet_0_clk _1068_/a_891_413# 0.00541f
C36101 acc0.A\[21\] _0382_ 0.02463f
C36102 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# 1.78756f
C36103 VPWR clkbuf_1_1__f_clk/a_110_47# 1.26537f
C36104 _1021_/a_27_47# _0385_ 0
C36105 _1021_/a_193_47# net220 0
C36106 net178 _1055_/a_1059_315# 0
C36107 _0415_ net80 0
C36108 _0374_ _0754_/a_512_297# 0.00102f
C36109 hold47/a_49_47# net10 0
C36110 _0101_ _0383_ 0
C36111 _0961_/a_199_47# control0.count\[1\] 0.01066f
C36112 hold30/a_49_47# hold30/a_285_47# 0.22264f
C36113 _0159_ _1061_/a_1059_315# 0
C36114 hold56/a_285_47# _0131_ 0.01838f
C36115 hold56/a_391_47# net119 0.02001f
C36116 _0403_ _0345_ 0.00488f
C36117 _1001_/a_27_47# _0195_ 0
C36118 _0346_ _0448_ 0
C36119 _1019_/a_27_47# _0350_ 0
C36120 net197 acc0.A\[29\] 0
C36121 clkbuf_1_0__f__0461_/a_110_47# _0391_ 0
C36122 net34 net236 0.01947f
C36123 net231 _1065_/a_466_413# 0
C36124 net39 _0346_ 0
C36125 _1019_/a_891_413# net105 0
C36126 _1019_/a_1059_315# net207 0
C36127 _0792_/a_209_297# net41 0.00274f
C36128 net35 _1071_/a_27_47# 0.00164f
C36129 _1008_/a_27_47# _0738_/a_68_297# 0.00156f
C36130 _0965_/a_377_297# control0.count\[3\] 0.00142f
C36131 net51 _1005_/a_1059_315# 0.09846f
C36132 hold21/a_285_47# input12/a_75_212# 0
C36133 _0539_/a_68_297# comp0.B\[11\] 0
C36134 net45 clknet_1_0__leaf__0459_ 0.09022f
C36135 hold98/a_391_47# _0297_ 0
C36136 _0256_ _0269_ 0.00368f
C36137 _0195_ hold8/a_49_47# 0.00379f
C36138 clknet_1_1__leaf__0460_ _0699_/a_150_297# 0
C36139 _0725_/a_303_47# _0333_ 0
C36140 VPWR _0584_/a_109_297# 0.18898f
C36141 _0343_ net50 0
C36142 _0760_/a_47_47# hold3/a_391_47# 0.006f
C36143 hold52/a_285_47# acc0.A\[24\] 0.11264f
C36144 hold83/a_391_47# net13 0.00363f
C36145 _0343_ _0995_/a_27_47# 0.0347f
C36146 _1014_/a_193_47# clknet_1_0__leaf__0461_ 0.04585f
C36147 _0726_/a_512_297# _0355_ 0.00103f
C36148 _0726_/a_245_297# net227 0
C36149 _0726_/a_149_47# _0354_ 0.0224f
C36150 acc0.A\[4\] _1045_/a_592_47# 0
C36151 _0324_ _0350_ 0
C36152 _0172_ hold6/a_285_47# 0.04652f
C36153 clkbuf_1_0__f__0461_/a_110_47# _0581_/a_27_297# 0.00614f
C36154 comp0.B\[14\] net152 0
C36155 net242 _1010_/a_381_47# 0
C36156 _0287_ _0655_/a_109_93# 0.00267f
C36157 net45 _0783_/a_79_21# 0.01012f
C36158 net9 acc0.A\[3\] 0
C36159 control0.state\[0\] _1064_/a_466_413# 0
C36160 net34 _1064_/a_193_47# 0.05531f
C36161 control0.state\[1\] _1064_/a_634_159# 0
C36162 _0274_ _0826_/a_219_297# 0.00378f
C36163 _0402_ hold70/a_391_47# 0
C36164 _0272_ _0826_/a_27_53# 0
C36165 clknet_1_0__leaf__0465_ input11/a_75_212# 0
C36166 _1033_/a_193_47# clknet_1_1__leaf__0463_ 0.00228f
C36167 _0130_ _1032_/a_466_413# 0
C36168 _1015_/a_466_413# _0584_/a_109_297# 0
C36169 _1015_/a_1059_315# _0584_/a_27_297# 0.01145f
C36170 _0692_/a_113_47# _0219_ 0
C36171 _0223_ net93 0
C36172 _1050_/a_27_47# _0148_ 0.09093f
C36173 net187 _0772_/a_297_297# 0
C36174 _1001_/a_634_159# _0247_ 0
C36175 clkbuf_0__0460_/a_110_47# _0460_ 0.32366f
C36176 _0369_ clknet_1_1__leaf__0458_ 0.90161f
C36177 _0951_/a_209_311# hold84/a_285_47# 0
C36178 net245 _0800_/a_149_47# 0.00446f
C36179 net58 _0844_/a_297_47# 0.04057f
C36180 _0739_/a_215_47# _0739_/a_510_47# 0.00529f
C36181 _0186_ net37 0
C36182 _0119_ _0578_/a_109_297# 0.00357f
C36183 _0843_/a_150_297# acc0.A\[15\] 0
C36184 _0195_ _1047_/a_193_47# 0
C36185 _0596_/a_145_75# net35 0
C36186 _1014_/a_27_47# _0265_ 0
C36187 _0352_ _0102_ 0.06376f
C36188 _0465_ _1048_/a_891_413# 0.0026f
C36189 acc0.A\[24\] net52 0.66981f
C36190 hold59/a_49_47# _1018_/a_27_47# 0.00693f
C36191 hold100/a_49_47# _0264_ 0.00784f
C36192 _0623_/a_109_297# acc0.A\[5\] 0.002f
C36193 _0294_ net77 0
C36194 _0990_/a_891_413# _0088_ 0.04061f
C36195 _0537_/a_150_297# VPWR 0.00237f
C36196 net125 _0498_/a_240_47# 0.00278f
C36197 _0546_/a_240_47# comp0.B\[9\] 0
C36198 comp0.B\[3\] _1066_/a_193_47# 0
C36199 _0174_ input31/a_75_212# 0
C36200 _0982_/a_193_47# _0264_ 0.00135f
C36201 _0610_/a_59_75# _0345_ 0.01129f
C36202 net88 clknet_1_0__leaf__0457_ 0.02488f
C36203 _0172_ _1041_/a_1017_47# 0
C36204 _0999_/a_634_159# _0345_ 0
C36205 acc0.A\[2\] _1048_/a_891_413# 0.00302f
C36206 _0136_ net8 0.07061f
C36207 _0793_/a_149_47# _0793_/a_240_47# 0.06872f
C36208 _0644_/a_47_47# acc0.A\[14\] 0.00111f
C36209 net152 _0543_/a_68_297# 0.17384f
C36210 _0343_ _0516_/a_27_297# 0
C36211 _0607_/a_109_297# _1017_/a_891_413# 0
C36212 acc0.A\[16\] _1017_/a_27_47# 0.00641f
C36213 _0482_ hold89/a_49_47# 0
C36214 pp[30] net239 0.001f
C36215 _0229_ _0381_ 0.06916f
C36216 _0211_ _1035_/a_193_47# 0
C36217 _0314_ _0740_/a_113_47# 0
C36218 net187 _0208_ 0
C36219 hold86/a_285_47# acc0.A\[1\] 0
C36220 hold86/a_49_47# _0182_ 0
C36221 _0539_/a_68_297# _0202_ 0.11423f
C36222 _0958_/a_197_47# _0468_ 0
C36223 _0243_ net46 0.07808f
C36224 comp0.B\[7\] _1039_/a_891_413# 0.0211f
C36225 pp[15] net42 0.0075f
C36226 _0123_ _1025_/a_1017_47# 0
C36227 _0195_ _0459_ 0.00846f
C36228 _0965_/a_47_47# clkbuf_1_0__f_clk/a_110_47# 0.0072f
C36229 _1051_/a_27_47# _1044_/a_27_47# 0.00214f
C36230 _0995_/a_634_159# acc0.A\[13\] 0
C36231 clkload4/Y _0369_ 0.02721f
C36232 _1037_/a_193_47# net28 0.02956f
C36233 _1034_/a_891_413# comp0.B\[6\] 0.01053f
C36234 _0777_/a_129_47# clknet_1_1__leaf__0461_ 0
C36235 net57 hold80/a_391_47# 0.08023f
C36236 _1051_/a_193_47# _1051_/a_592_47# 0
C36237 _1051_/a_466_413# _1051_/a_561_413# 0.00772f
C36238 _1051_/a_634_159# _1051_/a_975_413# 0
C36239 control0.sh _0175_ 0.35767f
C36240 _1045_/a_27_47# _1044_/a_634_159# 0
C36241 _1045_/a_193_47# _1044_/a_193_47# 0
C36242 _1045_/a_634_159# _1044_/a_27_47# 0.00897f
C36243 _1056_/a_561_413# clknet_1_1__leaf__0465_ 0
C36244 comp0.B\[14\] _1042_/a_466_413# 0
C36245 acc0.A\[21\] _1005_/a_634_159# 0
C36246 _0227_ _1005_/a_193_47# 0.00607f
C36247 net58 _0841_/a_297_297# 0.00327f
C36248 hold15/a_391_47# hold61/a_285_47# 0
C36249 VPWR _0439_ 0.66925f
C36250 _0992_/a_193_47# _0650_/a_150_297# 0
C36251 _0661_/a_27_297# clkbuf_1_1__f__0465_/a_110_47# 0
C36252 _0294_ _0656_/a_59_75# 0
C36253 acc0.A\[14\] net222 0.08543f
C36254 _0236_ _0238_ 0
C36255 net106 _1033_/a_1017_47# 0
C36256 _1070_/a_1017_47# _0168_ 0
C36257 _1045_/a_27_47# net184 0.21176f
C36258 _1045_/a_193_47# net131 0.01514f
C36259 _1045_/a_1059_315# _1045_/a_1017_47# 0
C36260 clkbuf_1_0__f__0464_/a_110_47# _0528_/a_299_297# 0
C36261 hold56/a_49_47# _1032_/a_27_47# 0
C36262 net23 _1067_/a_193_47# 0.12385f
C36263 net157 _0526_/a_27_47# 0.00699f
C36264 _0979_/a_109_297# clknet_1_0__leaf_clk 0
C36265 _1003_/a_27_47# net213 0
C36266 _0680_/a_80_21# _0346_ 0
C36267 _0251_ clknet_0__0458_ 0
C36268 clknet_0__0458_ _0640_/a_109_53# 0
C36269 VPWR _1043_/a_561_413# 0.00309f
C36270 _0852_/a_285_297# _0261_ 0
C36271 _0618_/a_79_21# _0219_ 0.02077f
C36272 hold63/a_49_47# hold63/a_391_47# 0.00188f
C36273 _0294_ _0986_/a_1059_315# 0
C36274 _0399_ _0397_ 0.04337f
C36275 _1018_/a_891_413# _0399_ 0
C36276 _0361_ _0697_/a_80_21# 0
C36277 _1043_/a_27_47# net196 0.10241f
C36278 _1043_/a_193_47# net129 0.0034f
C36279 _1043_/a_1059_315# _1043_/a_1017_47# 0
C36280 net9 net157 0
C36281 hold18/a_391_47# _0265_ 0.00137f
C36282 _0450_ _0264_ 0.0149f
C36283 VPWR _1015_/a_466_413# 0.25513f
C36284 net103 hold72/a_285_47# 0
C36285 _0217_ _0346_ 0.71882f
C36286 net160 input24/a_75_212# 0
C36287 _1034_/a_27_47# _1065_/a_193_47# 0
C36288 _0734_/a_129_47# acc0.A\[27\] 0
C36289 _0343_ _0399_ 0.11246f
C36290 A[7] hold83/a_285_47# 0
C36291 net124 _0209_ 0.00211f
C36292 clknet_1_1__leaf__0465_ _0281_ 0
C36293 _1030_/a_891_413# net208 0
C36294 VPWR _0654_/a_27_413# 0.2561f
C36295 _0275_ _0819_/a_299_297# 0.00596f
C36296 _1038_/a_1059_315# control0.sh 0
C36297 _0476_ hold89/a_49_47# 0
C36298 _0119_ _1002_/a_27_47# 0
C36299 _1021_/a_193_47# net88 0.02438f
C36300 _1021_/a_27_47# _0100_ 0.0058f
C36301 _0276_ _0218_ 0
C36302 output53/a_27_47# net52 0
C36303 net53 output52/a_27_47# 0
C36304 _1054_/a_1059_315# _1054_/a_891_413# 0.31086f
C36305 _1054_/a_193_47# _1054_/a_975_413# 0
C36306 _1054_/a_466_413# _1054_/a_381_47# 0.03733f
C36307 _1071_/a_1059_315# control0.count\[0\] 0
C36308 _1015_/a_634_159# _1015_/a_1059_315# 0
C36309 _1015_/a_27_47# _1015_/a_381_47# 0.06222f
C36310 _1015_/a_193_47# _1015_/a_891_413# 0.19489f
C36311 clknet_1_0__leaf__0458_ _0145_ 0.00179f
C36312 _0983_/a_381_47# VPWR 0.07234f
C36313 _0376_ net50 0
C36314 _0182_ clkbuf_1_0__f__0464_/a_110_47# 0
C36315 _0676_/a_113_47# _0308_ 0.00963f
C36316 _0991_/a_27_47# _0347_ 0
C36317 _0398_ acc0.A\[17\] 0
C36318 _0357_ _1010_/a_27_47# 0.00821f
C36319 _0439_ output62/a_27_47# 0
C36320 net247 _0261_ 0.25918f
C36321 net113 _1027_/a_634_159# 0
C36322 clknet_1_1__leaf__0462_ _1027_/a_1059_315# 0.01192f
C36323 clknet_0__0458_ net58 0.07815f
C36324 _0347_ _0773_/a_285_297# 0
C36325 VPWR output62/a_27_47# 0.43775f
C36326 net194 net130 0.08784f
C36327 _0752_/a_27_413# _0228_ 0
C36328 _0989_/a_193_47# output63/a_27_47# 0.00145f
C36329 net73 _0085_ 0
C36330 _0792_/a_209_47# _0400_ 0
C36331 _0343_ _1031_/a_27_47# 0.0231f
C36332 _0216_ net47 0
C36333 _0195_ _0265_ 0.00309f
C36334 _1038_/a_193_47# _1038_/a_381_47# 0.09784f
C36335 _1038_/a_634_159# _1038_/a_891_413# 0.03684f
C36336 _1038_/a_27_47# _1038_/a_561_413# 0.0027f
C36337 _1053_/a_193_47# _0180_ 0
C36338 _0246_ _0392_ 0
C36339 net62 net170 0
C36340 _0829_/a_109_297# _0435_ 0.00993f
C36341 _0319_ _1008_/a_466_413# 0
C36342 net48 VPWR 2.26407f
C36343 _0240_ clknet_1_0__leaf__0461_ 0
C36344 _0655_/a_109_93# _0655_/a_297_297# 0
C36345 _0655_/a_215_53# _0655_/a_369_297# 0.00854f
C36346 _0316_ _0350_ 0
C36347 VPWR input4/a_75_212# 0.24955f
C36348 clknet_0__0457_ clknet_1_0__leaf__0461_ 0.39266f
C36349 clknet_0__0461_ _0393_ 0.02465f
C36350 _0342_ _0218_ 0.04458f
C36351 _0446_ _0845_/a_193_297# 0.01408f
C36352 net61 _0529_/a_109_47# 0.00101f
C36353 clknet_1_0__leaf__0458_ _0446_ 0.05985f
C36354 _1050_/a_891_413# net10 0
C36355 _0157_ _1060_/a_1017_47# 0
C36356 _0536_/a_51_297# _0498_/a_51_297# 0
C36357 _0983_/a_634_159# _0983_/a_1017_47# 0
C36358 _0983_/a_466_413# _0983_/a_592_47# 0.00553f
C36359 net214 hold67/a_285_47# 0.02055f
C36360 _0981_/a_27_297# _0486_ 0
C36361 clknet_1_0__leaf__0465_ _1051_/a_975_413# 0
C36362 _0527_/a_109_297# _0142_ 0
C36363 hold59/a_285_47# _0242_ 0
C36364 _0183_ hold60/a_285_47# 0
C36365 _0081_ _0459_ 0
C36366 clknet_1_0__leaf__0465_ _1045_/a_1017_47# 0
C36367 _0261_ _0844_/a_382_297# 0
C36368 _0347_ _0350_ 0.58569f
C36369 _0262_ _0844_/a_297_47# 0
C36370 _0263_ _0844_/a_79_21# 0
C36371 net40 _0995_/a_1059_315# 0.16076f
C36372 net245 _0995_/a_634_159# 0.00221f
C36373 _0212_ _0557_/a_51_297# 0.00387f
C36374 _0423_ net228 0
C36375 net115 net191 0.02469f
C36376 _0965_/a_47_47# control0.count\[2\] 0.02193f
C36377 _0574_/a_27_297# _0574_/a_373_47# 0.01338f
C36378 hold89/a_49_47# hold89/a_285_47# 0.22264f
C36379 _0245_ _1006_/a_27_47# 0
C36380 _0985_/a_891_413# net71 0
C36381 _0286_ _0806_/a_199_47# 0
C36382 _0200_ _0139_ 0
C36383 _0854_/a_79_21# _0218_ 0
C36384 _0339_ net239 0
C36385 _0390_ VPWR 0.75539f
C36386 net31 _0547_/a_68_297# 0
C36387 hold50/a_285_47# _0345_ 0
C36388 hold44/a_285_47# net190 0
C36389 output64/a_27_47# acc0.A\[8\] 0
C36390 net71 _1049_/a_634_159# 0
C36391 hold77/a_285_47# _0397_ 0
C36392 _0747_/a_79_21# _1006_/a_193_47# 0
C36393 net219 hold72/a_391_47# 0.1417f
C36394 _0592_/a_68_297# net51 0.01488f
C36395 _0104_ _0350_ 0.21437f
C36396 _0466_ _1068_/a_466_413# 0.02422f
C36397 _1056_/a_193_47# _0154_ 0
C36398 _0459_ _0505_/a_373_47# 0
C36399 _0098_ acc0.A\[18\] 0
C36400 _0637_/a_139_47# _0269_ 0.00138f
C36401 _0118_ _0183_ 0.05317f
C36402 _1048_/a_634_159# _1047_/a_27_47# 0
C36403 _1048_/a_27_47# _1047_/a_634_159# 0
C36404 _1048_/a_193_47# _1047_/a_193_47# 0
C36405 _1003_/a_975_413# _0217_ 0
C36406 _0852_/a_35_297# _0265_ 0.01445f
C36407 _0852_/a_285_297# net47 0.00442f
C36408 net80 _0347_ 0
C36409 hold10/a_391_47# acc0.A\[15\] 0.06388f
C36410 _1016_/a_466_413# net166 0.00503f
C36411 _0244_ _0581_/a_373_47# 0.00182f
C36412 _0179_ _1056_/a_592_47# 0.00164f
C36413 net56 _1012_/a_1059_315# 0
C36414 _0719_/a_27_47# _0771_/a_27_413# 0
C36415 _0251_ net178 0
C36416 hold87/a_49_47# net206 0.00445f
C36417 control0.state\[1\] clknet_1_0__leaf__0460_ 0
C36418 net230 _0180_ 0.06275f
C36419 clknet_0__0459_ _0996_/a_891_413# 0
C36420 clknet_0__0465_ _0431_ 0.02314f
C36421 _0361_ _0743_/a_149_47# 0
C36422 net113 _1026_/a_891_413# 0
C36423 _0998_/a_27_47# _0096_ 0.11047f
C36424 _0998_/a_193_47# _0399_ 0.02409f
C36425 _0195_ _0220_ 0.21922f
C36426 _0414_ clknet_1_1__leaf__0459_ 0.00437f
C36427 _0277_ net5 0.00444f
C36428 hold17/a_285_47# VPWR 0.27452f
C36429 _0337_ hold61/a_285_47# 0.0048f
C36430 net189 net4 0.02338f
C36431 _0555_/a_512_297# _0176_ 0
C36432 _0354_ _0568_/a_109_297# 0
C36433 _0422_ _0090_ 0.02863f
C36434 clknet_0__0465_ _0659_/a_68_297# 0.00168f
C36435 hold37/a_49_47# _0180_ 0.00257f
C36436 net19 hold51/a_391_47# 0
C36437 _0433_ acc0.A\[6\] 0
C36438 _0361_ _0345_ 0
C36439 _0559_/a_245_297# VPWR 0.00631f
C36440 _0248_ _0346_ 0.64616f
C36441 _0258_ _0445_ 0
C36442 _0577_/a_109_297# hold4/a_285_47# 0
C36443 _0577_/a_27_297# hold4/a_391_47# 0.01653f
C36444 _0514_/a_373_47# _0189_ 0.00104f
C36445 net39 _0994_/a_592_47# 0.00257f
C36446 _1052_/a_27_47# net154 0
C36447 hold28/a_285_47# _0198_ 0
C36448 _0195_ _0585_/a_109_297# 0.00815f
C36449 _1032_/a_381_47# _0352_ 0
C36450 _1059_/a_1017_47# acc0.A\[14\] 0.00109f
C36451 _0985_/a_27_47# _0219_ 0
C36452 _0985_/a_1059_315# _0345_ 0
C36453 hold54/a_391_47# _0131_ 0
C36454 clknet_1_1__leaf__0459_ _1057_/a_891_413# 0
C36455 net160 _1035_/a_634_159# 0
C36456 _1057_/a_381_47# acc0.A\[11\] 0
C36457 hold48/a_49_47# _0201_ 0
C36458 net120 _0563_/a_51_297# 0
C36459 _0224_ net50 0.00151f
C36460 acc0.A\[0\] _0631_/a_109_297# 0
C36461 _1002_/a_1059_315# acc0.A\[21\] 0
C36462 net178 net58 0.02566f
C36463 _0677_/a_47_47# _0776_/a_27_47# 0
C36464 comp0.B\[4\] _1034_/a_634_159# 0
C36465 clknet_1_0__leaf__0459_ VPWR 3.7296f
C36466 net193 _0139_ 0
C36467 acc0.A\[20\] _0764_/a_81_21# 0
C36468 _0343_ _0299_ 0.02678f
C36469 _0753_/a_297_297# _0219_ 0
C36470 _0356_ hold95/a_391_47# 0
C36471 pp[7] pp[3] 0.18239f
C36472 _1056_/a_1059_315# net182 0.00113f
C36473 hold29/a_285_47# net176 0.0097f
C36474 _0107_ net95 0.00192f
C36475 hold18/a_391_47# _0267_ 0
C36476 _1054_/a_1017_47# VPWR 0
C36477 _0179_ _0989_/a_193_47# 0
C36478 _0179_ hold1/a_285_47# 0
C36479 _0275_ _0626_/a_68_297# 0.00419f
C36480 net2 _0744_/a_27_47# 0
C36481 VPWR _0569_/a_109_47# 0
C36482 net63 _0519_/a_384_47# 0
C36483 hold39/a_49_47# _0472_ 0
C36484 _0343_ _0712_/a_79_21# 0.18832f
C36485 clknet_1_0__leaf__0459_ _1015_/a_466_413# 0
C36486 hold34/a_391_47# net181 0.13119f
C36487 _0179_ _0992_/a_193_47# 0
C36488 _0174_ _0548_/a_51_297# 0.10856f
C36489 _0163_ _1065_/a_891_413# 0.00526f
C36490 VPWR _0783_/a_79_21# 0.47289f
C36491 _1038_/a_592_47# VPWR 0
C36492 _0338_ _0705_/a_59_75# 0.00941f
C36493 net64 output64/a_27_47# 0.24031f
C36494 hold11/a_391_47# net125 0.00207f
C36495 hold45/a_391_47# _0188_ 0.00178f
C36496 _0270_ _0196_ 0
C36497 VPWR _0283_ 1.40758f
C36498 _0989_/a_27_47# net75 0.21845f
C36499 hold1/a_49_47# net75 0
C36500 net35 _1072_/a_634_159# 0.00515f
C36501 net114 _0365_ 0.004f
C36502 _0731_/a_384_47# _0359_ 0
C36503 hold57/a_391_47# _0553_/a_51_297# 0
C36504 _1067_/a_466_413# _0460_ 0.00112f
C36505 A[12] clknet_1_1__leaf__0465_ 0.08199f
C36506 _1067_/a_891_413# clknet_1_0__leaf__0457_ 0.01246f
C36507 _0484_ _0468_ 0
C36508 _0148_ _0987_/a_27_47# 0
C36509 clkbuf_0__0465_/a_110_47# _0350_ 0.02989f
C36510 _0519_/a_299_297# _0191_ 0.00863f
C36511 net120 _1065_/a_592_47# 0
C36512 net188 _0515_/a_384_47# 0
C36513 _0473_ _0954_/a_32_297# 0.37176f
C36514 _0312_ _0250_ 0.95046f
C36515 _1059_/a_27_47# net41 0.00112f
C36516 comp0.B\[5\] net201 0
C36517 clkbuf_1_1__f__0463_/a_110_47# _0214_ 0.00741f
C36518 clknet_0__0463_ _0563_/a_240_47# 0.0049f
C36519 _1020_/a_193_47# net118 0.01042f
C36520 _0557_/a_512_297# net27 0
C36521 VPWR _0453_ 0.36068f
C36522 hold101/a_391_47# _0218_ 0.01852f
C36523 _0982_/a_27_47# hold18/a_49_47# 0
C36524 clknet_1_1__leaf__0459_ _0300_ 0.29646f
C36525 _1031_/a_193_47# _1030_/a_891_413# 0
C36526 _1031_/a_466_413# _1030_/a_466_413# 0
C36527 clknet_1_0__leaf__0464_ net7 0
C36528 _0424_ _0346_ 0.20392f
C36529 _0457_ _1067_/a_466_413# 0
C36530 VPWR _0794_/a_110_297# 0.00527f
C36531 clkbuf_1_1__f__0464_/a_110_47# _0954_/a_32_297# 0
C36532 hold68/a_49_47# hold29/a_285_47# 0
C36533 _0176_ _1045_/a_27_47# 0
C36534 _0298_ net5 0.13909f
C36535 acc0.A\[13\] _0345_ 0.02273f
C36536 _0507_/a_109_47# _0219_ 0.00239f
C36537 _1032_/a_1059_315# comp0.B\[15\] 0
C36538 _0180_ _0987_/a_381_47# 0
C36539 clknet_1_1__leaf__0460_ _0323_ 0.00107f
C36540 hold7/a_285_47# net148 0.06151f
C36541 _0554_/a_68_297# _1037_/a_891_413# 0.00287f
C36542 _0458_ acc0.A\[1\] 0.00139f
C36543 _0350_ hold95/a_49_47# 0
C36544 _1025_/a_193_47# _1025_/a_381_47# 0.09799f
C36545 _1025_/a_634_159# _1025_/a_891_413# 0.03684f
C36546 _1025_/a_27_47# _1025_/a_561_413# 0.0027f
C36547 _0355_ _0109_ 0.11475f
C36548 _1012_/a_1059_315# _0345_ 0
C36549 _1012_/a_27_47# _0219_ 0
C36550 clkbuf_1_0__f__0461_/a_110_47# _0116_ 0.00391f
C36551 hold35/a_391_47# VPWR 0.18432f
C36552 hold82/a_285_47# _0219_ 0
C36553 _0330_ _0219_ 0
C36554 net58 _0627_/a_109_93# 0.00137f
C36555 hold25/a_49_47# _0174_ 0.01278f
C36556 B[11] _0541_/a_68_297# 0.00173f
C36557 _0130_ net202 0
C36558 _0113_ _0584_/a_109_297# 0.00169f
C36559 _1015_/a_592_47# net157 0
C36560 _1055_/a_466_413# _0181_ 0
C36561 net205 net121 0
C36562 net238 hold91/a_285_47# 0.00948f
C36563 _0410_ hold91/a_49_47# 0.08826f
C36564 _0616_/a_78_199# _0391_ 0
C36565 _1070_/a_466_413# _0466_ 0
C36566 _1070_/a_1059_315# _0488_ 0
C36567 VPWR _0976_/a_535_374# 0
C36568 _0800_/a_149_47# VPWR 0.00398f
C36569 _0390_ clknet_1_0__leaf__0459_ 0
C36570 _0130_ clknet_1_1__leaf__0463_ 0.00148f
C36571 _0352_ hold72/a_391_47# 0
C36572 _0330_ _0728_/a_59_75# 0
C36573 _0157_ _0508_/a_81_21# 0.14641f
C36574 hold54/a_49_47# _1032_/a_193_47# 0
C36575 hold49/a_49_47# _0954_/a_32_297# 0
C36576 clkbuf_1_0__f__0457_/a_110_47# _0772_/a_215_47# 0
C36577 _1046_/a_381_47# net10 0.01664f
C36578 clknet_0__0457_ _1001_/a_1017_47# 0
C36579 _0955_/a_32_297# _0175_ 0.0011f
C36580 _0118_ hold40/a_285_47# 0.00152f
C36581 acc0.A\[11\] _0808_/a_81_21# 0
C36582 _0982_/a_193_47# _0856_/a_79_21# 0.00587f
C36583 net181 _0181_ 0.00372f
C36584 clknet_0__0463_ _0935_/a_27_47# 0
C36585 _1021_/a_193_47# _1067_/a_891_413# 0
C36586 hold17/a_49_47# hold17/a_391_47# 0.00188f
C36587 _0403_ _0994_/a_27_47# 0.00647f
C36588 _0645_/a_47_47# _0346_ 0
C36589 clknet_0__0463_ _1061_/a_193_47# 0
C36590 _0516_/a_109_297# _0990_/a_891_413# 0
C36591 net61 _0845_/a_193_297# 0
C36592 A[10] net67 0
C36593 net61 clknet_1_0__leaf__0458_ 0
C36594 B[8] net153 0
C36595 net31 net127 0.13882f
C36596 hold18/a_49_47# _0446_ 0.00111f
C36597 _1003_/a_1059_315# control0.state\[2\] 0
C36598 _0996_/a_1059_315# _0996_/a_891_413# 0.31086f
C36599 _0996_/a_193_47# _0996_/a_975_413# 0
C36600 _0996_/a_466_413# _0996_/a_381_47# 0.03733f
C36601 _1055_/a_193_47# _0517_/a_81_21# 0
C36602 _1055_/a_27_47# _0517_/a_299_297# 0
C36603 _0852_/a_35_297# _0267_ 0
C36604 _0769_/a_384_47# _0352_ 0
C36605 _0244_ _0347_ 0.02839f
C36606 net92 net51 0
C36607 net45 _1031_/a_634_159# 0
C36608 VPWR _0835_/a_493_297# 0.00248f
C36609 clknet_0__0464_ comp0.B\[12\] 0
C36610 _0728_/a_145_75# _0333_ 0.00192f
C36611 net2 net66 0.10535f
C36612 _0473_ net173 0
C36613 _0216_ net93 0
C36614 hold64/a_49_47# clknet_1_0__leaf__0461_ 0.0176f
C36615 clknet_1_0__leaf__0464_ _1048_/a_1059_315# 0
C36616 _0329_ hold50/a_391_47# 0
C36617 clknet_1_1__leaf__0457_ _1061_/a_634_159# 0.00221f
C36618 _0343_ _0190_ 0
C36619 _0375_ _0345_ 0
C36620 _0234_ _0377_ 0.04919f
C36621 _1060_/a_27_47# net6 0.00587f
C36622 _0732_/a_209_297# _0219_ 0.00256f
C36623 _0559_/a_51_297# _0559_/a_512_297# 0.0116f
C36624 hold57/a_49_47# _0475_ 0
C36625 _0317_ _0686_/a_219_297# 0.00642f
C36626 _0642_/a_27_413# _0369_ 0.00498f
C36627 acc0.A\[4\] _0180_ 0.02927f
C36628 _1057_/a_193_47# clknet_1_1__leaf__0465_ 0.10166f
C36629 VPWR _0996_/a_1017_47# 0
C36630 VPWR _1036_/a_27_47# 0.67056f
C36631 _0621_/a_285_297# clkbuf_1_1__f__0458_/a_110_47# 0
C36632 _1065_/a_1017_47# comp0.B\[0\] 0
C36633 _0330_ _1008_/a_634_159# 0
C36634 _1044_/a_27_47# _1044_/a_193_47# 0.96851f
C36635 _0774_/a_68_297# hold72/a_285_47# 0
C36636 _0672_/a_215_47# clkbuf_1_1__f__0459_/a_110_47# 0
C36637 _0272_ _0640_/a_215_297# 0.10602f
C36638 VPWR _0523_/a_81_21# 0.21422f
C36639 comp0.B\[2\] comp0.B\[5\] 0.0056f
C36640 hold24/a_285_47# comp0.B\[10\] 0
C36641 clknet_0__0465_ _0269_ 0.00483f
C36642 _1051_/a_1059_315# acc0.A\[5\] 0.08398f
C36643 hold65/a_285_47# net212 0.00769f
C36644 net182 VPWR 0.34399f
C36645 hold22/a_285_47# _1054_/a_891_413# 0.00163f
C36646 hold65/a_49_47# _0437_ 0
C36647 hold22/a_391_47# _1054_/a_1059_315# 0.00124f
C36648 hold64/a_285_47# net47 0
C36649 net131 _1044_/a_27_47# 0.00302f
C36650 _1045_/a_27_47# net130 0.00992f
C36651 acc0.A\[21\] net91 0
C36652 hold59/a_285_47# _0855_/a_81_21# 0
C36653 _0992_/a_561_413# acc0.A\[10\] 0
C36654 _1030_/a_561_413# _0353_ 0
C36655 _0293_ clkbuf_1_1__f__0465_/a_110_47# 0
C36656 net62 _0986_/a_1017_47# 0.00175f
C36657 _0374_ acc0.A\[23\] 0
C36658 clknet_1_1__leaf__0459_ _0404_ 0.15426f
C36659 net164 control0.count\[0\] 0.0104f
C36660 _0736_/a_311_297# VPWR 0.0046f
C36661 _0399_ _0990_/a_381_47# 0.01646f
C36662 _0432_ acc0.A\[4\] 0
C36663 _0179_ net142 0.15987f
C36664 net56 _0726_/a_51_297# 0
C36665 control0.state\[0\] hold93/a_49_47# 0
C36666 _0299_ A[14] 0
C36667 _1051_/a_1059_315# _0528_/a_299_297# 0
C36668 _0399_ _0793_/a_51_297# 0
C36669 _0789_/a_75_199# VPWR 0.16547f
C36670 _0442_ hold1/a_49_47# 0.00263f
C36671 _0272_ _0465_ 0.0266f
C36672 hold100/a_285_47# _0449_ 0.00111f
C36673 _0537_/a_68_297# _0172_ 0
C36674 clkbuf_1_0__f__0459_/a_110_47# _0399_ 0.11388f
C36675 _1002_/a_561_413# net240 0
C36676 net245 _0345_ 0
C36677 _1039_/a_193_47# clknet_0__0463_ 0.02521f
C36678 _1060_/a_466_413# net229 0
C36679 _0714_/a_51_297# _1013_/a_466_413# 0.0044f
C36680 _0714_/a_149_47# _1013_/a_27_47# 0
C36681 VPWR _0113_ 0.2369f
C36682 _1003_/a_891_413# _0467_ 0
C36683 _0644_/a_377_297# net41 0.0012f
C36684 clknet_1_1__leaf__0460_ net237 0
C36685 clkbuf_0__0464_/a_110_47# _0142_ 0.09969f
C36686 _1030_/a_27_47# _0219_ 0.00891f
C36687 _1072_/a_193_47# net159 0
C36688 _0972_/a_250_297# _1062_/a_193_47# 0
C36689 _0972_/a_93_21# _1062_/a_634_159# 0
C36690 hold76/a_391_47# _1000_/a_27_47# 0
C36691 hold76/a_285_47# _1000_/a_193_47# 0
C36692 _0662_/a_81_21# _0817_/a_266_47# 0
C36693 _0849_/a_79_21# _0849_/a_297_297# 0.01735f
C36694 clknet_1_0__leaf__0463_ _1040_/a_381_47# 0
C36695 _0502_/a_27_47# _0171_ 0
C36696 acc0.A\[12\] output67/a_27_47# 0
C36697 hold101/a_49_47# _0987_/a_27_47# 0
C36698 _0218_ _0240_ 0
C36699 _1032_/a_634_159# _1032_/a_592_47# 0
C36700 _1054_/a_381_47# net169 0.12476f
C36701 net9 net13 0.02166f
C36702 _1015_/a_466_413# _0113_ 0.0209f
C36703 net247 _0173_ 0
C36704 _0369_ _0218_ 0.06772f
C36705 _1038_/a_381_47# net29 0
C36706 hold5/a_391_47# _0176_ 0
C36707 clknet_0__0457_ _0218_ 0
C36708 _0235_ _0346_ 0.03972f
C36709 hold31/a_285_47# _0186_ 0
C36710 hold14/a_285_47# net28 0
C36711 _0343_ _0327_ 0
C36712 _1051_/a_466_413# _0180_ 0.01719f
C36713 _0435_ _0827_/a_27_47# 0.05426f
C36714 _0820_/a_297_297# _0990_/a_27_47# 0
C36715 _1014_/a_193_47# _0112_ 0.18441f
C36716 _1014_/a_381_47# net149 0.02661f
C36717 _0769_/a_81_21# _0773_/a_35_297# 0.00217f
C36718 VPWR net30 0.57383f
C36719 _1038_/a_1059_315# net172 0
C36720 _1038_/a_891_413# net124 0
C36721 init _1066_/a_891_413# 0
C36722 net33 _1066_/a_1059_315# 0.04302f
C36723 hold21/a_49_47# hold21/a_285_47# 0.22264f
C36724 _0472_ _0159_ 0.08868f
C36725 hold8/a_391_47# _1026_/a_1059_315# 0
C36726 _1067_/a_1017_47# clknet_1_0__leaf__0461_ 0
C36727 _0551_/a_27_47# _0533_/a_109_297# 0
C36728 hold75/a_285_47# VPWR 0.27988f
C36729 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk 0.31698f
C36730 _0401_ _0422_ 0.00128f
C36731 _0960_/a_27_47# _1069_/a_1059_315# 0
C36732 _0750_/a_27_47# _0383_ 0.04662f
C36733 net54 _0697_/a_217_297# 0
C36734 clknet_1_0__leaf__0465_ _1044_/a_592_47# 0
C36735 net45 _0345_ 0.0645f
C36736 _0170_ _0486_ 0.00402f
C36737 hold16/a_391_47# _1030_/a_634_159# 0.00982f
C36738 hold16/a_285_47# _1030_/a_466_413# 0.01371f
C36739 hold16/a_49_47# _1030_/a_1059_315# 0.00923f
C36740 _1020_/a_634_159# net1 0.0185f
C36741 hold12/a_391_47# _1068_/a_1059_315# 0
C36742 _0350_ _0106_ 0
C36743 _0234_ net109 0
C36744 _0997_/a_466_413# net43 0.02503f
C36745 _0227_ _0762_/a_215_47# 0
C36746 net198 hold51/a_285_47# 0.01718f
C36747 VPWR pp[22] 0.21099f
C36748 VPWR _0995_/a_634_159# 0.1842f
C36749 _0285_ _0993_/a_27_47# 0
C36750 _0454_ _0450_ 0.0024f
C36751 _0461_ _0181_ 0.00113f
C36752 _0304_ hold81/a_49_47# 0
C36753 clknet_1_1__leaf__0458_ _0084_ 0
C36754 net72 _0445_ 0.08068f
C36755 net247 _0848_/a_109_297# 0
C36756 net7 _0547_/a_68_297# 0
C36757 hold13/a_49_47# net28 0
C36758 _0511_/a_81_21# _0187_ 0.20733f
C36759 _0347_ _0986_/a_634_159# 0.00127f
C36760 acc0.A\[26\] _0320_ 0.11469f
C36761 _0280_ _0670_/a_79_21# 0
C36762 net90 net51 0
C36763 _0550_/a_51_297# net180 0.12933f
C36764 _0240_ _0775_/a_215_47# 0.00237f
C36765 net190 _1008_/a_634_159# 0
C36766 _0371_ _1006_/a_1059_315# 0
C36767 net216 _1006_/a_891_413# 0.00134f
C36768 _0104_ _1006_/a_634_159# 0.00367f
C36769 _0533_/a_27_297# _0533_/a_109_297# 0.17136f
C36770 _0354_ _0725_/a_209_297# 0
C36771 _0726_/a_149_47# _0353_ 0
C36772 _0355_ _0725_/a_80_21# 0.08183f
C36773 net106 _1032_/a_381_47# 0
C36774 _0466_ _0166_ 0.13317f
C36775 hold32/a_285_47# _1055_/a_891_413# 0
C36776 hold31/a_391_47# _0253_ 0.03293f
C36777 _1000_/a_466_413# _0461_ 0.00375f
C36778 _0186_ _0524_/a_109_297# 0.01564f
C36779 _0684_/a_59_75# acc0.A\[27\] 0.09f
C36780 clknet_1_0__leaf__0462_ _1005_/a_1017_47# 0
C36781 VPWR comp0.B\[3\] 0.7455f
C36782 _1061_/a_1017_47# acc0.A\[15\] 0
C36783 _0247_ _0245_ 0
C36784 _0249_ acc0.A\[23\] 0
C36785 _0546_/a_51_297# _0546_/a_149_47# 0.02487f
C36786 VPWR _1023_/a_27_47# 0.68903f
C36787 hold100/a_49_47# _0846_/a_51_297# 0
C36788 _1036_/a_891_413# _0175_ 0.01807f
C36789 _0163_ hold93/a_285_47# 0
C36790 hold101/a_285_47# net63 0.00475f
C36791 _0534_/a_384_47# _0182_ 0
C36792 _0991_/a_27_47# _0991_/a_1059_315# 0.04875f
C36793 _0991_/a_193_47# _0991_/a_466_413# 0.07911f
C36794 _0534_/a_299_297# net218 0.01949f
C36795 VPWR _0516_/a_109_47# 0
C36796 net84 _0398_ 0.04342f
C36797 _0726_/a_51_297# _0345_ 0.10768f
C36798 _0315_ hold90/a_285_47# 0.01164f
C36799 _1054_/a_1059_315# _0255_ 0
C36800 _0263_ _0084_ 0
C36801 clkbuf_1_0__f__0458_/a_110_47# _0267_ 0.03141f
C36802 _0587_/a_27_47# _0345_ 0.02048f
C36803 _0397_ _0306_ 0.01988f
C36804 net23 clkbuf_1_1__f__0457_/a_110_47# 0
C36805 _0241_ _0771_/a_382_47# 0.0011f
C36806 _0195_ _0178_ 0.02122f
C36807 _1041_/a_193_47# net22 0
C36808 _0120_ hold4/a_391_47# 0.04366f
C36809 acc0.A\[19\] hold60/a_49_47# 0
C36810 _0210_ _0957_/a_220_297# 0
C36811 _0554_/a_68_297# _0475_ 0
C36812 net160 _0957_/a_304_297# 0
C36813 acc0.A\[20\] _0372_ 0
C36814 _0343_ _0576_/a_27_297# 0
C36815 net61 hold18/a_49_47# 0
C36816 _1052_/a_975_413# net11 0
C36817 hold46/a_285_47# net7 0
C36818 _0833_/a_215_47# _0369_ 0.05716f
C36819 net236 _0166_ 0.05065f
C36820 net160 net121 0
C36821 _1001_/a_634_159# _0217_ 0
C36822 _1001_/a_27_47# _0183_ 0.15246f
C36823 hold6/a_49_47# _1040_/a_634_159# 0
C36824 hold6/a_285_47# _1040_/a_193_47# 0
C36825 net186 _0173_ 0.01698f
C36826 hold39/a_391_47# _0132_ 0.00138f
C36827 net55 _0334_ 0.10423f
C36828 _0399_ _0996_/a_193_47# 0.03343f
C36829 acc0.A\[17\] _0308_ 0.02025f
C36830 control0.count\[2\] clknet_0_clk 0
C36831 net23 _0951_/a_109_93# 0
C36832 _0808_/a_81_21# _0281_ 0.03456f
C36833 _0229_ _0762_/a_79_21# 0
C36834 _1021_/a_27_47# net150 0
C36835 hold54/a_49_47# hold54/a_391_47# 0.00188f
C36836 _0579_/a_373_47# VPWR 0
C36837 _0548_/a_51_297# comp0.B\[9\] 0.11449f
C36838 _1041_/a_193_47# clknet_1_0__leaf__0463_ 0.03905f
C36839 _0125_ hold9/a_49_47# 0.29201f
C36840 _0174_ _0540_/a_149_47# 0.02112f
C36841 acc0.A\[20\] hold40/a_49_47# 0.32351f
C36842 net11 net75 0
C36843 _0348_ _0705_/a_59_75# 0.00214f
C36844 clknet_0__0461_ _0773_/a_35_297# 0
C36845 _1058_/a_193_47# acc0.A\[10\] 0.01008f
C36846 net48 _1023_/a_27_47# 0.00191f
C36847 _1067_/a_193_47# _0161_ 0
C36848 clknet_1_0__leaf__0459_ _0113_ 0
C36849 _0366_ _1007_/a_975_413# 0
C36850 _0430_ acc0.A\[8\] 0.01721f
C36851 _0446_ _0846_/a_245_297# 0.00131f
C36852 _0713_/a_27_47# net87 0
C36853 _0476_ _0469_ 0
C36854 comp0.B\[10\] _0138_ 0
C36855 hold65/a_391_47# _0434_ 0
C36856 _0258_ _0440_ 0
C36857 _0722_/a_79_21# _0352_ 0.14517f
C36858 _0522_/a_109_47# acc0.A\[6\] 0
C36859 _0257_ _0442_ 0.00338f
C36860 _1050_/a_975_413# clknet_1_1__leaf__0464_ 0
C36861 output66/a_27_47# _0179_ 0.01247f
C36862 clknet_0__0457_ _0112_ 0.00465f
C36863 _0181_ _0465_ 0.03007f
C36864 _0196_ _0085_ 0
C36865 _0663_/a_27_413# _0663_/a_207_413# 0.18542f
C36866 _0463_ _0496_/a_27_47# 0
C36867 VPWR _0697_/a_80_21# 0.23899f
C36868 _0290_ _0291_ 0.25302f
C36869 acc0.A\[5\] acc0.A\[8\] 0.00647f
C36870 _0401_ acc0.A\[8\] 0.00854f
C36871 _1017_/a_975_413# _0369_ 0
C36872 _0399_ clkbuf_0__0461_/a_110_47# 0
C36873 _1002_/a_466_413# _0352_ 0
C36874 pp[17] _1031_/a_1059_315# 0.01686f
C36875 net167 _1068_/a_27_47# 0.01281f
C36876 _0490_ _1068_/a_193_47# 0
C36877 clknet_1_0__leaf__0462_ _0762_/a_79_21# 0
C36878 VPWR net56 0.97019f
C36879 _0296_ _0303_ 0.0441f
C36880 VPWR _0695_/a_217_297# 0.20378f
C36881 net168 input15/a_75_212# 0.04132f
C36882 _1011_/a_27_47# _0350_ 0
C36883 hold29/a_49_47# _1023_/a_1059_315# 0.00336f
C36884 acc0.A\[2\] _0181_ 0
C36885 control0.count\[3\] _0488_ 0.01599f
C36886 _0627_/a_297_297# _0254_ 0.00247f
C36887 _1033_/a_1059_315# _1067_/a_27_47# 0
C36888 _1004_/a_193_47# net52 0.0178f
C36889 VPWR _1031_/a_634_159# 0.18231f
C36890 clkbuf_0__0465_/a_110_47# _0986_/a_634_159# 0.00581f
C36891 _0381_ _0382_ 0.07184f
C36892 _0134_ net27 0.00728f
C36893 _0195_ _1019_/a_27_47# 0
C36894 net178 _0988_/a_975_413# 0
C36895 hold31/a_391_47# net74 0.02312f
C36896 _0217_ net221 0.24502f
C36897 _0290_ _0991_/a_634_159# 0
C36898 _0401_ _0991_/a_193_47# 0
C36899 _0425_ _0991_/a_27_47# 0
C36900 _0983_/a_975_413# _0399_ 0
C36901 _0749_/a_384_47# _0460_ 0
C36902 pp[23] _1022_/a_891_413# 0
C36903 _0200_ _0954_/a_32_297# 0
C36904 _0490_ _0478_ 0
C36905 hold26/a_391_47# VPWR 0.1873f
C36906 _0515_/a_81_21# acc0.A\[11\] 0
C36907 _1031_/a_27_47# _0568_/a_27_297# 0
C36908 net36 net175 0
C36909 clknet_1_0__leaf__0465_ net10 0.01245f
C36910 _0955_/a_32_297# _0955_/a_114_297# 0.01439f
C36911 hold76/a_49_47# _0242_ 0.02128f
C36912 hold76/a_391_47# acc0.A\[19\] 0.02137f
C36913 hold35/a_391_47# net182 0.13432f
C36914 hold23/a_391_47# net10 0.039f
C36915 _1004_/a_634_159# clknet_1_0__leaf__0460_ 0.01495f
C36916 _0216_ _0581_/a_109_297# 0
C36917 _1025_/a_193_47# acc0.A\[25\] 0.0875f
C36918 net49 _0103_ 0
C36919 _0296_ _0281_ 0.02207f
C36920 net207 _0264_ 0
C36921 _1030_/a_891_413# _0221_ 0
C36922 _0183_ _0459_ 1.26847f
C36923 pp[15] net60 0
C36924 hold72/a_285_47# hold72/a_391_47# 0.41909f
C36925 hold36/a_391_47# _0172_ 0.00802f
C36926 hold89/a_391_47# _0468_ 0.00312f
C36927 _0369_ net240 0.0341f
C36928 hold65/a_49_47# _0252_ 0
C36929 hold64/a_49_47# _0218_ 0
C36930 net179 _0181_ 0
C36931 hold65/a_285_47# _0989_/a_891_413# 0.00677f
C36932 hold65/a_391_47# _0989_/a_1059_315# 0.00126f
C36933 _0168_ _0466_ 0.02425f
C36934 _0179_ _0988_/a_27_47# 0
C36935 _1001_/a_466_413# control0.add 0
C36936 hold20/a_285_47# _1072_/a_27_47# 0.00123f
C36937 _0369_ _0099_ 0.00129f
C36938 _0425_ _0350_ 0
C36939 clknet_0__0457_ _0099_ 0.01437f
C36940 _0474_ _0175_ 0.02254f
C36941 comp0.B\[6\] _0215_ 0
C36942 clknet_1_1__leaf__0459_ _0419_ 0.02253f
C36943 net38 _0091_ 0
C36944 net7 net127 0.04867f
C36945 _1021_/a_27_47# control0.add 0
C36946 hold22/a_285_47# hold22/a_391_47# 0.41909f
C36947 net233 _0449_ 0.18319f
C36948 _0260_ hold100/a_285_47# 0
C36949 _0101_ _0486_ 0
C36950 VPWR _0808_/a_266_47# 0.00238f
C36951 _1055_/a_1059_315# _0153_ 0.02743f
C36952 net217 hold70/a_285_47# 0.0078f
C36953 _0422_ hold70/a_49_47# 0.00806f
C36954 _0315_ clknet_0__0462_ 0.0402f
C36955 _0358_ _0332_ 0.00233f
C36956 _1047_/a_193_47# acc0.A\[15\] 0
C36957 net64 _0430_ 0.1709f
C36958 _0769_/a_299_297# _0769_/a_384_47# 0
C36959 net64 _0621_/a_285_47# 0.00124f
C36960 _0317_ clknet_1_1__leaf__0462_ 0.00126f
C36961 pp[1] net47 0.01614f
C36962 clkload2/Y clknet_1_0__leaf__0465_ 0.00374f
C36963 _0217_ _0782_/a_27_47# 0
C36964 _0231_ acc0.A\[23\] 0.23609f
C36965 clknet_0__0458_ _0625_/a_145_75# 0
C36966 _0369_ _0359_ 0
C36967 _0993_/a_27_47# _0218_ 0
C36968 _0994_/a_27_47# acc0.A\[13\] 0
C36969 net133 net134 0
C36970 _0358_ _0685_/a_68_297# 0
C36971 hold87/a_285_47# hold87/a_391_47# 0.41909f
C36972 clknet_1_1__leaf__0457_ net147 0.00103f
C36973 net15 _0369_ 0
C36974 hold30/a_285_47# _0222_ 0
C36975 _0525_/a_81_21# net73 0.00209f
C36976 _0662_/a_81_21# _0181_ 0.0082f
C36977 _1060_/a_592_47# _0184_ 0
C36978 _0274_ _0831_/a_35_297# 0.01509f
C36979 hold101/a_49_47# clkbuf_1_0__f__0465_/a_110_47# 0.02088f
C36980 net45 _0791_/a_113_297# 0
C36981 hold24/a_49_47# _0555_/a_51_297# 0
C36982 _0433_ _0826_/a_219_297# 0
C36983 _0343_ _0346_ 1.0508f
C36984 _1041_/a_634_159# _0544_/a_51_297# 0
C36985 _0176_ _0546_/a_51_297# 0.00128f
C36986 hold8/a_49_47# net156 0.01412f
C36987 clknet_1_0__leaf__0463_ _1039_/a_592_47# 0
C36988 clkbuf_1_1__f__0459_/a_110_47# _0669_/a_29_53# 0.01151f
C36989 _1050_/a_466_413# _0524_/a_27_297# 0
C36990 comp0.B\[7\] _0136_ 0
C36991 _0330_ net94 0
C36992 _0437_ _0828_/a_199_47# 0.00144f
C36993 _0144_ clknet_1_1__leaf__0464_ 0
C36994 _0200_ net173 0
C36995 _1059_/a_193_47# clkbuf_0__0459_/a_110_47# 0.00812f
C36996 net44 _0776_/a_27_47# 0
C36997 _1065_/a_466_413# _0564_/a_68_297# 0
C36998 _1044_/a_466_413# _1044_/a_592_47# 0.00553f
C36999 _1044_/a_634_159# _1044_/a_1017_47# 0
C37000 _0654_/a_27_413# _0808_/a_266_47# 0
C37001 _0178_ _1048_/a_193_47# 0
C37002 _0554_/a_68_297# net27 0.00242f
C37003 comp0.B\[13\] _0954_/a_220_297# 0.00703f
C37004 _0272_ _0254_ 0.02571f
C37005 net193 _0954_/a_32_297# 0.0113f
C37006 net158 _0536_/a_512_297# 0
C37007 _0529_/a_27_297# _0529_/a_109_297# 0.17136f
C37008 _1038_/a_381_47# comp0.B\[6\] 0
C37009 _0343_ net65 0.0015f
C37010 hold52/a_285_47# net199 0.02264f
C37011 hold41/a_391_47# _1058_/a_466_413# 0.0056f
C37012 hold41/a_285_47# _1058_/a_1059_315# 0.002f
C37013 hold41/a_49_47# _1058_/a_891_413# 0.00283f
C37014 _0328_ _0692_/a_113_47# 0
C37015 _0423_ _0401_ 0.2596f
C37016 _0985_/a_193_47# _0465_ 0
C37017 _0971_/a_299_297# _1062_/a_27_47# 0
C37018 _0971_/a_81_21# _1062_/a_193_47# 0
C37019 _0459_ acc0.A\[15\] 0.13722f
C37020 VPWR _0743_/a_149_47# 0.00162f
C37021 _0183_ _0265_ 0
C37022 _0958_/a_27_47# _0972_/a_93_21# 0
C37023 net180 _0913_/a_27_47# 0
C37024 _0140_ _0541_/a_68_297# 0
C37025 clknet_1_1__leaf__0458_ net75 0.13644f
C37026 net173 comp0.B\[8\] 0.00359f
C37027 net55 output59/a_27_47# 0
C37028 net36 _1038_/a_193_47# 0.16387f
C37029 clknet_1_1__leaf_clk _1065_/a_466_413# 0.01483f
C37030 _0180_ _0350_ 0
C37031 _0278_ pp[13] 0
C37032 _0387_ clknet_0__0461_ 0
C37033 _0329_ _0726_/a_245_297# 0
C37034 _0624_/a_59_75# _0835_/a_78_199# 0
C37035 net44 _0219_ 0.09781f
C37036 _0985_/a_27_47# net58 0.00838f
C37037 _0985_/a_193_47# acc0.A\[2\] 0.00613f
C37038 _0237_ _1005_/a_193_47# 0.00145f
C37039 pp[19] _1023_/a_975_413# 0
C37040 net46 _1023_/a_1017_47# 0
C37041 _0216_ _1028_/a_634_159# 0
C37042 _0195_ _1028_/a_1059_315# 0.05104f
C37043 _1067_/a_561_413# net17 0
C37044 hold42/a_49_47# hold42/a_285_47# 0.22264f
C37045 hold42/a_49_47# _1057_/a_1059_315# 0
C37046 _1051_/a_975_413# _0148_ 0
C37047 hold49/a_391_47# net20 0.04223f
C37048 _1057_/a_193_47# _1057_/a_381_47# 0.09503f
C37049 _1057_/a_634_159# _1057_/a_891_413# 0.03684f
C37050 _1057_/a_27_47# _1057_/a_561_413# 0.0027f
C37051 VPWR _0814_/a_27_47# 0.20818f
C37052 VPWR _0345_ 9.97101f
C37053 hold48/a_391_47# hold49/a_285_47# 0.00113f
C37054 B[13] _1042_/a_27_47# 0.00105f
C37055 _0269_ _0986_/a_27_47# 0
C37056 _0579_/a_109_297# net87 0
C37057 pp[17] _0712_/a_561_47# 0
C37058 net21 B[11] 0.07647f
C37059 _0111_ _1013_/a_193_47# 0.37815f
C37060 _0158_ net229 0
C37061 net225 _1013_/a_466_413# 0
C37062 VPWR _1064_/a_466_413# 0.25507f
C37063 _0854_/a_215_47# _0116_ 0
C37064 _0552_/a_68_297# net171 0.00163f
C37065 _0199_ clkbuf_0__0463_/a_110_47# 0
C37066 _1059_/a_27_47# _1059_/a_561_413# 0.0027f
C37067 _1059_/a_634_159# _1059_/a_891_413# 0.03684f
C37068 _1059_/a_193_47# _1059_/a_381_47# 0.09972f
C37069 net199 net52 0.17557f
C37070 net248 _0256_ 0
C37071 net231 _1062_/a_634_159# 0.00199f
C37072 _0164_ _1062_/a_193_47# 0.0011f
C37073 _0458_ _0198_ 0
C37074 _0849_/a_215_47# _0082_ 0
C37075 _0259_ _0424_ 0
C37076 _1015_/a_466_413# _0345_ 0
C37077 net55 _0724_/a_113_297# 0
C37078 net248 _0987_/a_1059_315# 0
C37079 _0179_ _1047_/a_193_47# 0
C37080 net125 clknet_1_1__leaf__0457_ 0.02505f
C37081 hold37/a_391_47# clknet_1_1__leaf__0464_ 0.00752f
C37082 VPWR hold2/a_49_47# 0.28381f
C37083 _0654_/a_27_413# _0345_ 0.00385f
C37084 _0820_/a_79_21# clknet_1_1__leaf__0465_ 0.02454f
C37085 _1065_/a_1059_315# clkbuf_1_1__f_clk/a_110_47# 0.0152f
C37086 _0552_/a_68_297# net24 0
C37087 _0181_ _0582_/a_27_297# 0
C37088 _0573_/a_27_47# _0178_ 0.26095f
C37089 _0481_ _0978_/a_373_47# 0.00186f
C37090 _0149_ _0180_ 0.07102f
C37091 net193 _0540_/a_245_297# 0
C37092 comp0.B\[13\] _0540_/a_149_47# 0.00184f
C37093 hold46/a_285_47# _0202_ 0.01274f
C37094 acc0.A\[0\] net149 0.03954f
C37095 clknet_1_0__leaf__0460_ clknet_1_1__leaf_clk 0
C37096 _0783_/a_510_47# _0398_ 0.00378f
C37097 _0783_/a_215_47# _0399_ 0.02844f
C37098 net45 _0394_ 0
C37099 hold8/a_49_47# acc0.A\[26\] 0.32737f
C37100 _1046_/a_1059_315# _0540_/a_51_297# 0
C37101 _0349_ _0705_/a_145_75# 0
C37102 _0385_ _0352_ 0.12452f
C37103 _0265_ acc0.A\[15\] 0
C37104 net61 _0846_/a_245_297# 0
C37105 acc0.A\[27\] _1028_/a_975_413# 0
C37106 _0328_ _0618_/a_79_21# 0
C37107 comp0.B\[14\] comp0.B\[12\] 0.07922f
C37108 net40 _0994_/a_634_159# 0
C37109 hold38/a_391_47# _1062_/a_193_47# 0
C37110 _0960_/a_181_47# clknet_1_0__leaf_clk 0
C37111 hold16/a_49_47# VPWR 0.26425f
C37112 _0179_ _0459_ 0
C37113 net48 _0345_ 0
C37114 _0144_ net247 0
C37115 _0369_ net228 0.11628f
C37116 _0218_ pp[31] 0
C37117 _1052_/a_1059_315# _0186_ 0
C37118 _0195_ _0347_ 0.02159f
C37119 _0352_ _1006_/a_1017_47# 0
C37120 net197 clknet_1_1__leaf__0462_ 0.07945f
C37121 net186 _1033_/a_1059_315# 0
C37122 _1058_/a_193_47# _0188_ 0.00153f
C37123 clknet_1_0__leaf__0458_ _0269_ 0.00333f
C37124 _0386_ clkbuf_1_0__f__0461_/a_110_47# 0
C37125 _1056_/a_27_47# _1055_/a_1059_315# 0.00914f
C37126 net14 _0179_ 0.00945f
C37127 clkload1/a_268_47# VPWR 0
C37128 _0972_/a_250_297# net17 0
C37129 clkbuf_1_0__f__0464_/a_110_47# _1048_/a_1059_315# 0.0015f
C37130 net46 clknet_1_0__leaf__0460_ 0.03724f
C37131 _0217_ _0585_/a_373_47# 0
C37132 acc0.A\[11\] _0652_/a_109_297# 0
C37133 clknet_0__0465_ clkbuf_0__0458_/a_110_47# 0
C37134 _0094_ net6 0
C37135 _0399_ _0794_/a_326_47# 0.00105f
C37136 acc0.A\[14\] net229 0.04156f
C37137 _1014_/a_1059_315# clkbuf_0__0457_/a_110_47# 0.00129f
C37138 _0340_ net209 0
C37139 hold28/a_391_47# net134 0
C37140 _0216_ _0371_ 0
C37141 _0107_ hold69/a_49_47# 0
C37142 pp[9] acc0.A\[10\] 0
C37143 net180 _0172_ 0.02758f
C37144 net190 net94 0
C37145 _0390_ _0345_ 0
C37146 _0104_ net92 0
C37147 _0533_/a_109_297# _0199_ 0.00191f
C37148 _0533_/a_373_47# net8 0.00194f
C37149 hold43/a_391_47# _0126_ 0
C37150 _0951_/a_209_311# _1062_/a_381_47# 0
C37151 net35 _0486_ 0.05554f
C37152 hold66/a_285_47# net51 0.00364f
C37153 control0.state\[0\] control0.count\[0\] 0
C37154 _0282_ _0091_ 0
C37155 _0183_ _1060_/a_381_47# 0.01149f
C37156 clkbuf_1_1__f__0463_/a_110_47# _0472_ 0
C37157 clknet_0__0458_ hold86/a_49_47# 0
C37158 _0555_/a_512_297# net28 0
C37159 net169 _0193_ 0
C37160 B[12] _0203_ 0
C37161 hold87/a_285_47# _0264_ 0.00439f
C37162 _0098_ _0461_ 0.00325f
C37163 clknet_1_0__leaf__0462_ _1022_/a_634_159# 0.00591f
C37164 _0123_ _1024_/a_634_159# 0
C37165 net108 _1022_/a_27_47# 0.22551f
C37166 hold23/a_49_47# _0449_ 0
C37167 _1005_/a_27_47# _1005_/a_193_47# 0.9705f
C37168 net11 hold83/a_285_47# 0
C37169 _0978_/a_109_297# _0484_ 0
C37170 _0978_/a_27_297# _0485_ 0
C37171 _0369_ hold3/a_285_47# 0
C37172 _0376_ hold94/a_49_47# 0
C37173 _0375_ hold94/a_391_47# 0
C37174 _0546_/a_240_47# net32 0.05893f
C37175 hold75/a_49_47# hold75/a_391_47# 0.00188f
C37176 _0399_ acc0.A\[6\] 0.79747f
C37177 _0546_/a_245_297# _0139_ 0
C37178 _1047_/a_1059_315# clknet_1_1__leaf__0457_ 0.00936f
C37179 _0473_ clknet_1_1__leaf__0457_ 0
C37180 hold45/a_49_47# VPWR 0.36432f
C37181 _0446_ _0448_ 0.21078f
C37182 net149 _0580_/a_109_297# 0.00203f
C37183 _0991_/a_891_413# _0991_/a_1017_47# 0.00617f
C37184 _0991_/a_193_47# _0089_ 0.31328f
C37185 _0346_ net38 0
C37186 _0991_/a_634_159# net77 0
C37187 control0.state\[0\] clknet_1_0__leaf__0457_ 0
C37188 _0442_ clknet_1_1__leaf__0458_ 0.01648f
C37189 _0536_/a_149_47# net134 0
C37190 _0236_ _0384_ 0.19028f
C37191 _0370_ _1006_/a_891_413# 0
C37192 _0356_ net97 0
C37193 net82 _0305_ 0
C37194 _0817_/a_81_21# _0218_ 0
C37195 _0817_/a_266_297# _0294_ 0
C37196 comp0.B\[4\] control0.sh 0.04732f
C37197 net205 _0555_/a_51_297# 0
C37198 _0260_ _0270_ 0
C37199 _0985_/a_27_47# _0262_ 0.0016f
C37200 _0583_/a_27_297# _1060_/a_27_47# 0
C37201 _0216_ _1029_/a_975_413# 0
C37202 hold52/a_285_47# VPWR 0.29612f
C37203 clknet_1_1__leaf__0459_ _0992_/a_193_47# 0.04301f
C37204 _0217_ _0973_/a_27_297# 0
C37205 _0183_ _0267_ 0
C37206 _0460_ hold73/a_285_47# 0.00741f
C37207 _0411_ acc0.A\[13\] 0
C37208 net178 _0833_/a_79_21# 0
C37209 _0982_/a_466_413# acc0.A\[0\] 0.00506f
C37210 _0982_/a_561_413# net100 0
C37211 VPWR _1065_/a_1059_315# 0.40631f
C37212 _0174_ _0542_/a_245_297# 0.00206f
C37213 _0107_ clkbuf_0__0462_/a_110_47# 0
C37214 _0363_ _0462_ 0
C37215 _0600_/a_103_199# _0600_/a_253_47# 0.06061f
C37216 net78 net67 0.02414f
C37217 net140 _0150_ 0
C37218 _0195_ _1016_/a_891_413# 0
C37219 _0725_/a_303_47# acc0.A\[29\] 0
C37220 _0995_/a_27_47# _0995_/a_1059_315# 0.04875f
C37221 _0995_/a_193_47# _0995_/a_466_413# 0.08183f
C37222 _0529_/a_27_297# net170 0.12233f
C37223 _0413_ _0297_ 0
C37224 clknet_1_0__leaf__0457_ _0610_/a_59_75# 0
C37225 _0357_ _0701_/a_303_47# 0.00402f
C37226 _0230_ _0383_ 0.00146f
C37227 _0543_/a_150_297# _0202_ 0
C37228 _1021_/a_975_413# _0183_ 0.00176f
C37229 clknet_0__0458_ acc0.A\[14\] 0
C37230 hold87/a_49_47# clknet_1_0__leaf__0458_ 0.00242f
C37231 _1060_/a_381_47# acc0.A\[15\] 0.00209f
C37232 _1002_/a_1059_315# _0381_ 0
C37233 _0081_ _0347_ 0.09691f
C37234 _0501_/a_27_47# _0533_/a_27_297# 0
C37235 clknet_1_0__leaf__0459_ _0345_ 0.06341f
C37236 VPWR net52 1.53041f
C37237 _0529_/a_27_297# _0845_/a_109_297# 0
C37238 hold9/a_285_47# _1027_/a_193_47# 0.00369f
C37239 hold9/a_391_47# _1027_/a_27_47# 0
C37240 hold9/a_49_47# _1027_/a_634_159# 0.00169f
C37241 VPWR _0819_/a_81_21# 0.21012f
C37242 _0218_ _0084_ 0.00422f
C37243 hold101/a_285_47# _0824_/a_59_75# 0
C37244 _1050_/a_193_47# _0142_ 0.00372f
C37245 _0398_ _0777_/a_129_47# 0
C37246 _0467_ clknet_1_0__leaf__0461_ 0
C37247 net53 _1007_/a_891_413# 0.02753f
C37248 _0976_/a_439_47# _0466_ 0.00508f
C37249 _0723_/a_27_413# acc0.A\[30\] 0
C37250 net34 _1062_/a_193_47# 0
C37251 control0.state\[0\] _1062_/a_466_413# 0.00328f
C37252 control0.state\[1\] _1062_/a_634_159# 0.02569f
C37253 net46 _0576_/a_109_297# 0.00114f
C37254 _0412_ _0413_ 0.20307f
C37255 _0800_/a_240_47# _0093_ 0.00121f
C37256 _0982_/a_27_47# _0217_ 0
C37257 acc0.A\[16\] hold72/a_49_47# 0
C37258 VPWR _0836_/a_68_297# 0.15908f
C37259 _1034_/a_1059_315# _0957_/a_32_297# 0
C37260 output64/a_27_47# _0369_ 0.00155f
C37261 acc0.A\[27\] net191 0
C37262 _0368_ _0460_ 0
C37263 _0346_ hold81/a_285_47# 0
C37264 _0305_ _0115_ 0
C37265 _0225_ acc0.A\[23\] 0
C37266 _0100_ _0352_ 0.14961f
C37267 _0283_ _0345_ 0.06371f
C37268 _1011_/a_193_47# _1011_/a_381_47# 0.09799f
C37269 _1011_/a_634_159# _1011_/a_891_413# 0.03684f
C37270 _1011_/a_27_47# _1011_/a_561_413# 0.00163f
C37271 _0814_/a_27_47# _0283_ 0
C37272 _1016_/a_1059_315# _0369_ 0.027f
C37273 VPWR net212 0.14896f
C37274 _0402_ acc0.A\[10\] 0
C37275 hold10/a_391_47# _0171_ 0.04014f
C37276 _0133_ _1034_/a_27_47# 0.01651f
C37277 net233 _0260_ 0
C37278 output47/a_27_47# net62 0.05158f
C37279 _0217_ _0145_ 0
C37280 _1034_/a_1059_315# net23 0
C37281 _0241_ control0.add 0
C37282 hold85/a_49_47# _0164_ 0.36819f
C37283 _0350_ _1006_/a_381_47# 0.0232f
C37284 _0304_ _0286_ 0
C37285 clknet_0__0465_ _0986_/a_975_413# 0
C37286 _0183_ net51 0.01785f
C37287 _0289_ _0992_/a_27_47# 0
C37288 net45 _0997_/a_193_47# 0.00118f
C37289 _0714_/a_240_47# _0216_ 0
C37290 acc0.A\[12\] _0279_ 0.33098f
C37291 net39 _0278_ 0.11884f
C37292 _0267_ acc0.A\[15\] 0.04809f
C37293 _0130_ _1067_/a_466_413# 0
C37294 _0423_ _0089_ 0.08701f
C37295 _0179_ _1056_/a_975_413# 0
C37296 clkbuf_0_clk/a_110_47# _0181_ 0
C37297 comp0.B\[0\] clknet_1_0__leaf__0461_ 0.00274f
C37298 net210 _1025_/a_193_47# 0
C37299 _0195_ _1025_/a_27_47# 0
C37300 _1055_/a_27_47# VPWR 0.72287f
C37301 hold67/a_285_47# _0186_ 0
C37302 _0347_ net90 0.28448f
C37303 _1020_/a_561_413# VPWR 0.00332f
C37304 _0453_ _0345_ 0.0189f
C37305 VPWR _0791_/a_113_297# 0.25295f
C37306 _0217_ net17 0
C37307 _0803_/a_68_297# _0277_ 0
C37308 _0982_/a_1059_315# _0580_/a_27_297# 0
C37309 _0181_ _1063_/a_634_159# 0.01044f
C37310 _0163_ _1063_/a_27_47# 0
C37311 _0534_/a_81_21# _0146_ 0
C37312 _0955_/a_304_297# comp0.B\[6\] 0.00104f
C37313 _0458_ net247 0
C37314 net57 hold95/a_285_47# 0.00459f
C37315 _0195_ hold95/a_49_47# 0.05309f
C37316 hold44/a_391_47# acc0.A\[29\] 0.05122f
C37317 clknet_1_0__leaf__0463_ net133 0
C37318 _0311_ _0748_/a_384_47# 0
C37319 _0292_ _0427_ 0.2433f
C37320 _0966_/a_109_297# _0488_ 0.00122f
C37321 control0.reset net201 0.37661f
C37322 _0217_ _0446_ 0
C37323 net240 _1067_/a_1017_47# 0
C37324 _0165_ _1067_/a_561_413# 0.0016f
C37325 clknet_1_0__leaf__0465_ _0492_/a_27_47# 0
C37326 _1042_/a_27_47# _1042_/a_634_159# 0.13601f
C37327 net245 _0411_ 0
C37328 _0511_/a_81_21# clknet_1_1__leaf__0465_ 0
C37329 _0181_ _1060_/a_634_159# 0.04563f
C37330 net54 _1008_/a_1017_47# 0
C37331 control0.state\[2\] net159 0.19016f
C37332 net44 hold61/a_49_47# 0.00832f
C37333 _0172_ _0545_/a_150_297# 0
C37334 _0175_ _0563_/a_51_297# 0.03802f
C37335 clkbuf_1_0__f__0457_/a_110_47# net105 0
C37336 _0290_ _0656_/a_59_75# 0
C37337 _1010_/a_634_159# _0352_ 0.01546f
C37338 acc0.A\[30\] _0352_ 0
C37339 _0531_/a_27_297# _0465_ 0.00771f
C37340 clknet_1_1__leaf__0460_ _0730_/a_215_47# 0
C37341 _1051_/a_891_413# clknet_1_1__leaf__0464_ 0
C37342 hold63/a_285_47# _0216_ 0.01301f
C37343 hold63/a_391_47# net155 0.00245f
C37344 _0800_/a_149_47# _0345_ 0.00164f
C37345 net22 comp0.B\[10\] 0.0229f
C37346 _0458_ _0844_/a_382_297# 0
C37347 _1036_/a_634_159# _1036_/a_592_47# 0
C37348 _0714_/a_51_297# _0339_ 0.00925f
C37349 clkbuf_1_1__f__0464_/a_110_47# net19 0
C37350 _0290_ _0986_/a_1059_315# 0
C37351 _0313_ acc0.A\[25\] 0.31825f
C37352 acc0.A\[2\] _0531_/a_27_297# 0
C37353 _0346_ _0793_/a_51_297# 0
C37354 hold26/a_285_47# _0172_ 0.00515f
C37355 _0480_ _0484_ 0.05337f
C37356 _0517_/a_299_297# _0988_/a_1059_315# 0
C37357 _0578_/a_109_297# net187 0.0015f
C37358 _0644_/a_47_47# _0276_ 0.1453f
C37359 VPWR _1040_/a_27_47# 0.42359f
C37360 _0725_/a_209_297# _0353_ 0.02819f
C37361 _0646_/a_47_47# _0300_ 0
C37362 _0179_ _0267_ 0.02128f
C37363 A[7] net13 0.00202f
C37364 _1050_/a_891_413# net12 0
C37365 _0227_ net150 0.02033f
C37366 acc0.A\[21\] _0217_ 0.07384f
C37367 _0238_ _0240_ 0
C37368 clknet_1_0__leaf__0463_ comp0.B\[10\] 0.02584f
C37369 clkbuf_1_1__f_clk/a_110_47# hold93/a_49_47# 0.00189f
C37370 net36 net29 0
C37371 pp[28] hold62/a_391_47# 0
C37372 output56/a_27_47# net209 0.0033f
C37373 _0467_ clk 0
C37374 _0529_/a_373_47# net10 0
C37375 net158 _0144_ 0.22311f
C37376 net82 _0181_ 0.00381f
C37377 clknet_1_0__leaf__0462_ _1026_/a_193_47# 0
C37378 _0236_ _0383_ 0
C37379 _0238_ _0369_ 0.02616f
C37380 hold13/a_49_47# clknet_0__0463_ 0.00102f
C37381 _0483_ _0981_/a_109_47# 0
C37382 _0965_/a_47_47# _0170_ 0.0035f
C37383 hold49/a_49_47# net19 0
C37384 hold49/a_285_47# net195 0
C37385 _0497_/a_68_297# clknet_1_1__leaf__0457_ 0
C37386 VPWR _0394_ 0.5889f
C37387 _0576_/a_109_47# VPWR 0
C37388 _0163_ _1062_/a_1059_315# 0.00612f
C37389 clknet_1_0__leaf__0462_ _1024_/a_891_413# 0.00358f
C37390 _0467_ _1063_/a_891_413# 0.00352f
C37391 _1058_/a_1059_315# net4 0.0564f
C37392 _1058_/a_634_159# _0187_ 0
C37393 _0477_ _0972_/a_93_21# 0.01668f
C37394 _0416_ acc0.A\[12\] 0
C37395 hold32/a_285_47# net47 0.001f
C37396 _0467_ _0959_/a_217_297# 0.04895f
C37397 net58 _0990_/a_27_47# 0
C37398 hold19/a_391_47# _0583_/a_27_297# 0.01653f
C37399 hold19/a_285_47# _0583_/a_109_297# 0
C37400 _1032_/a_27_47# _1067_/a_27_47# 0
C37401 _0777_/a_47_47# _0395_ 0.14353f
C37402 _1049_/a_592_47# _0465_ 0
C37403 net165 clknet_1_0__leaf__0461_ 0
C37404 net187 net202 0.00181f
C37405 net194 _0142_ 0.11706f
C37406 _0476_ hold39/a_285_47# 0
C37407 clkload0/a_27_47# clknet_0_clk 0.02356f
C37408 _0582_/a_27_297# clknet_1_1__leaf__0461_ 0.01184f
C37409 clkbuf_0__0461_/a_110_47# _0306_ 0
C37410 clkbuf_1_0__f__0458_/a_110_47# _0347_ 0.01887f
C37411 net61 _0448_ 0.07839f
C37412 _1012_/a_466_413# net239 0
C37413 _0381_ net91 0
C37414 _1054_/a_27_47# acc0.A\[7\] 0
C37415 _0216_ net114 0
C37416 _1054_/a_1059_315# _0989_/a_27_47# 0
C37417 hold42/a_285_47# net189 0.0104f
C37418 pp[9] _0188_ 0.08341f
C37419 clkbuf_1_1__f__0463_/a_110_47# _1033_/a_27_47# 0.01577f
C37420 _0803_/a_150_297# _0404_ 0.00135f
C37421 hold10/a_285_47# control0.sh 0
C37422 clkbuf_0__0463_/a_110_47# _0498_/a_149_47# 0
C37423 _0463_ _0498_/a_51_297# 0
C37424 _0648_/a_27_297# _0403_ 0
C37425 acc0.A\[16\] clknet_0__0461_ 0.1119f
C37426 _1053_/a_193_47# _1052_/a_27_47# 0.00148f
C37427 _1053_/a_27_47# _1052_/a_193_47# 0.00114f
C37428 _0579_/a_27_297# net211 0.05719f
C37429 _0093_ _0995_/a_466_413# 0
C37430 _0789_/a_208_47# _0298_ 0.00102f
C37431 _1059_/a_891_413# net145 0
C37432 _0789_/a_75_199# _0345_ 0
C37433 _0732_/a_209_297# _0328_ 0.00656f
C37434 _0754_/a_51_297# _0754_/a_149_47# 0.02487f
C37435 _0643_/a_103_199# _0270_ 0
C37436 comp0.B\[2\] control0.reset 0.73874f
C37437 _0951_/a_109_93# _0161_ 0.09586f
C37438 input14/a_75_212# _0150_ 0
C37439 _0217_ _0245_ 0
C37440 net188 _0186_ 0
C37441 VPWR input10/a_75_212# 0.26637f
C37442 _0196_ net170 0.08672f
C37443 _0113_ _0345_ 0
C37444 clknet_1_0__leaf__0461_ acc0.A\[19\] 0.16776f
C37445 _0322_ clkbuf_0__0462_/a_110_47# 0.01572f
C37446 _0313_ _0737_/a_117_297# 0
C37447 _0642_/a_27_413# net75 0
C37448 _0490_ VPWR 0.287f
C37449 _0619_/a_68_297# acc0.A\[6\] 0
C37450 _1055_/a_466_413# clknet_1_1__leaf__0465_ 0.00919f
C37451 _0855_/a_299_297# _0465_ 0
C37452 net120 _0173_ 0.00552f
C37453 _0779_/a_79_21# _0352_ 0.13456f
C37454 _0710_/a_109_297# _0342_ 0.23298f
C37455 _0176_ _1042_/a_891_413# 0.00229f
C37456 _0779_/a_510_47# _0347_ 0
C37457 _0327_ clkbuf_0__0462_/a_110_47# 0.13474f
C37458 _0767_/a_145_75# _0369_ 0
C37459 _0673_/a_103_199# _0304_ 0.12614f
C37460 _0673_/a_253_297# _0295_ 0
C37461 clknet_1_0__leaf__0458_ _0082_ 0.13125f
C37462 _0555_/a_51_297# net160 0.10201f
C37463 _0352_ _0771_/a_382_47# 0.00271f
C37464 _0181_ _0115_ 0
C37465 net14 hold83/a_49_47# 0
C37466 _1038_/a_1059_315# _0549_/a_68_297# 0.00603f
C37467 net181 clknet_1_1__leaf__0465_ 0
C37468 net46 hold94/a_285_47# 0
C37469 _0304_ _0672_/a_79_21# 0.05051f
C37470 _0310_ _0352_ 0.00132f
C37471 net69 _0219_ 0
C37472 _1002_/a_891_413# _0578_/a_109_297# 0
C37473 clknet_0__0457_ _0721_/a_27_47# 0
C37474 _0407_ _0791_/a_199_47# 0.00151f
C37475 _1051_/a_27_47# _0524_/a_27_297# 0
C37476 _0672_/a_215_47# _0296_ 0.05773f
C37477 clkload3/a_110_47# _0459_ 0
C37478 _0454_ _0849_/a_79_21# 0
C37479 _0992_/a_634_159# _0281_ 0
C37480 hold23/a_49_47# _0260_ 0
C37481 _1030_/a_592_47# clknet_1_1__leaf__0462_ 0
C37482 net61 _0444_ 0
C37483 _0369_ _0090_ 0.15869f
C37484 _1046_/a_891_413# net20 0
C37485 net231 _0132_ 0
C37486 _0971_/a_81_21# net17 0
C37487 _1053_/a_27_47# net12 0.03887f
C37488 net83 _0408_ 0
C37489 _0536_/a_149_47# net22 0
C37490 control0.state\[1\] hold85/a_285_47# 0
C37491 control0.state\[0\] hold85/a_391_47# 0.01355f
C37492 net34 hold85/a_49_47# 0
C37493 net81 net41 0
C37494 VPWR _0994_/a_27_47# 0.69234f
C37495 _0974_/a_448_47# _1068_/a_27_47# 0
C37496 VPWR _1008_/a_592_47# 0
C37497 _0478_ control0.count\[0\] 0.15346f
C37498 _0981_/a_27_297# clknet_0_clk 0.00293f
C37499 hold43/a_285_47# VPWR 0.27991f
C37500 output60/a_27_47# output41/a_27_47# 0.02615f
C37501 _0461_ _1015_/a_27_47# 0.056f
C37502 _0216_ _0365_ 0
C37503 _0195_ _0106_ 0
C37504 clkload2/a_110_47# clkload2/Y 0.00568f
C37505 clkbuf_1_1__f__0458_/a_110_47# _0825_/a_68_297# 0.01503f
C37506 _0338_ hold62/a_49_47# 0.00225f
C37507 _0222_ _1005_/a_193_47# 0
C37508 net239 net98 0
C37509 _0785_/a_81_21# _0428_ 0.00199f
C37510 _0785_/a_299_297# _0427_ 0
C37511 _0305_ _1017_/a_891_413# 0.01206f
C37512 _0341_ _1013_/a_1059_315# 0.00188f
C37513 _0340_ _1013_/a_466_413# 0
C37514 _0342_ _1013_/a_27_47# 0
C37515 hold10/a_285_47# net157 0.05866f
C37516 net14 input13/a_75_212# 0.04425f
C37517 clknet_1_0__leaf__0463_ _0536_/a_149_47# 0.0011f
C37518 _0218_ hold40/a_391_47# 0
C37519 _0164_ net17 0.07737f
C37520 _0369_ _0760_/a_285_47# 0.00494f
C37521 _0305_ net146 0
C37522 net50 _0377_ 0
C37523 VPWR hold93/a_49_47# 0.28273f
C37524 comp0.B\[4\] _0955_/a_32_297# 0.12629f
C37525 _0343_ _0259_ 0.03067f
C37526 _0695_/a_80_21# _0695_/a_472_297# 0.01636f
C37527 _1010_/a_1059_315# hold95/a_285_47# 0.0054f
C37528 _0361_ hold90/a_391_47# 0
C37529 net248 clknet_0__0465_ 0
C37530 comp0.B\[10\] _0544_/a_245_297# 0.00322f
C37531 _1031_/a_27_47# _1031_/a_1059_315# 0.04875f
C37532 _1031_/a_193_47# _1031_/a_466_413# 0.07855f
C37533 _0292_ _0818_/a_193_47# 0
C37534 _0517_/a_384_47# _0186_ 0
C37535 input31/a_75_212# net32 0
C37536 _0996_/a_193_47# _0346_ 0
C37537 _0804_/a_79_21# _0403_ 0.0967f
C37538 _0457_ _1034_/a_381_47# 0
C37539 hold30/a_285_47# net243 0
C37540 _0476_ hold57/a_391_47# 0
C37541 _1000_/a_27_47# _0218_ 0
C37542 _1000_/a_193_47# _0294_ 0.00163f
C37543 _0123_ net110 0.00123f
C37544 hold53/a_285_47# acc0.A\[24\] 0
C37545 _1005_/a_634_159# _1005_/a_1017_47# 0
C37546 _1005_/a_466_413# _1005_/a_592_47# 0.00553f
C37547 clkbuf_0__0458_/a_110_47# _0986_/a_27_47# 0
C37548 net178 hold88/a_391_47# 0
C37549 _0769_/a_81_21# _0247_ 0.01404f
C37550 _0244_ _0616_/a_292_297# 0
C37551 hold66/a_49_47# net49 0.32126f
C37552 VPWR _0156_ 0.22728f
C37553 _0519_/a_81_21# _0152_ 0.13864f
C37554 _0984_/a_1059_315# _0082_ 0
C37555 _0984_/a_561_413# net222 0
C37556 _0192_ net12 0
C37557 _1060_/a_1059_315# _0507_/a_109_297# 0
C37558 _0646_/a_47_47# _0646_/a_285_47# 0.01755f
C37559 _1013_/a_1059_315# _1013_/a_891_413# 0.31086f
C37560 _1013_/a_193_47# _1013_/a_975_413# 0
C37561 _1013_/a_466_413# _1013_/a_381_47# 0.03733f
C37562 _0991_/a_592_47# net67 0
C37563 _1002_/a_27_47# _1002_/a_891_413# 0.03224f
C37564 _1002_/a_193_47# _1002_/a_1059_315# 0.03405f
C37565 _1002_/a_634_159# _1002_/a_466_413# 0.23992f
C37566 VPWR _0527_/a_373_47# 0
C37567 _1027_/a_634_159# _0739_/a_79_21# 0
C37568 _0821_/a_113_47# VPWR 0
C37569 _0985_/a_27_47# hold28/a_49_47# 0.00377f
C37570 clknet_1_1__leaf__0460_ clkbuf_1_0__f__0462_/a_110_47# 0.0011f
C37571 _0984_/a_193_47# clknet_1_0__leaf__0458_ 0.02395f
C37572 _1027_/a_27_47# _0352_ 0
C37573 _1027_/a_466_413# _0347_ 0
C37574 net243 _0102_ 0.04105f
C37575 _1017_/a_1059_315# net43 0.00435f
C37576 _0985_/a_1017_47# _0261_ 0
C37577 clknet_1_1__leaf__0459_ _0997_/a_975_413# 0
C37578 net165 _1060_/a_891_413# 0
C37579 clknet_0_clk hold84/a_391_47# 0
C37580 _0178_ acc0.A\[15\] 0.00552f
C37581 net59 _0350_ 0
C37582 _0612_/a_59_75# _0611_/a_68_297# 0.0083f
C37583 _0108_ _1012_/a_27_47# 0
C37584 hold35/a_391_47# _1055_/a_27_47# 0
C37585 hold35/a_285_47# _1055_/a_193_47# 0
C37586 VPWR _0989_/a_891_413# 0.17143f
C37587 _0248_ _0245_ 0
C37588 _0217_ _0165_ 0
C37589 VPWR _0997_/a_193_47# 0.32253f
C37590 _0080_ acc0.A\[0\] 0.23193f
C37591 _0795_/a_299_297# _0405_ 0.07411f
C37592 _0795_/a_81_21# _0400_ 0
C37593 _1038_/a_466_413# _1040_/a_381_47# 0
C37594 _0217_ _1019_/a_634_159# 0.0092f
C37595 _0183_ _1019_/a_27_47# 0.024f
C37596 _0690_/a_68_297# _0319_ 0.04293f
C37597 VPWR _0992_/a_891_413# 0.19396f
C37598 _0362_ _0733_/a_222_93# 0
C37599 _0734_/a_129_47# _0361_ 0.00412f
C37600 _0438_ _0465_ 0
C37601 _1018_/a_891_413# net221 0.00319f
C37602 _1018_/a_27_47# _0115_ 0
C37603 control0.state\[0\] _0958_/a_109_47# 0
C37604 control0.state\[1\] _0958_/a_27_47# 0.24463f
C37605 _0154_ _0515_/a_81_21# 0.13864f
C37606 VPWR hold94/a_391_47# 0.17182f
C37607 _0768_/a_27_47# _0352_ 0.00223f
C37608 _0995_/a_891_413# _0995_/a_1017_47# 0.00617f
C37609 hold65/a_391_47# _0186_ 0.00176f
C37610 _1035_/a_27_47# _0175_ 0.03658f
C37611 net10 _0148_ 0
C37612 output56/a_27_47# _1011_/a_634_159# 0
C37613 VPWR _1061_/a_466_413# 0.25819f
C37614 clknet_1_1__leaf__0459_ _0668_/a_297_47# 0.00214f
C37615 hold23/a_285_47# _0447_ 0
C37616 _0343_ net221 0.0492f
C37617 _0234_ _0460_ 0.00172f
C37618 _0636_/a_59_75# _0465_ 0.00137f
C37619 _0501_/a_27_47# _0199_ 0.1085f
C37620 _0783_/a_79_21# _0394_ 0
C37621 VPWR net171 0.36744f
C37622 net63 output63/a_27_47# 0.2402f
C37623 _0534_/a_299_297# _1048_/a_891_413# 0
C37624 net36 acc0.A\[18\] 0
C37625 _1034_/a_466_413# _0173_ 0.00926f
C37626 _1034_/a_27_47# _0208_ 0
C37627 _1034_/a_1059_315# _0213_ 0.00401f
C37628 acc0.A\[12\] _0512_/a_27_297# 0
C37629 clknet_1_0__leaf__0464_ _0197_ 0.00188f
C37630 _0529_/a_109_297# _0449_ 0
C37631 hold87/a_285_47# _0454_ 0.00169f
C37632 _1035_/a_193_47# control0.sh 0.00425f
C37633 _0183_ _0581_/a_373_47# 0.00162f
C37634 net36 _0137_ 0.13045f
C37635 net77 _0986_/a_1059_315# 0
C37636 _0736_/a_311_297# net52 0
C37637 net117 _0704_/a_68_297# 0
C37638 _1000_/a_27_47# _0775_/a_215_47# 0
C37639 _0800_/a_51_297# _0799_/a_80_21# 0
C37640 hold54/a_285_47# _0216_ 0.0011f
C37641 net232 control0.state\[2\] 0
C37642 clknet_1_0__leaf__0458_ clkbuf_0__0458_/a_110_47# 0
C37643 _1018_/a_561_413# _0459_ 0
C37644 _1019_/a_891_413# _0580_/a_109_297# 0
C37645 _0327_ _0725_/a_80_21# 0
C37646 _0168_ _1069_/a_1059_315# 0.00454f
C37647 _1070_/a_193_47# control0.count\[0\] 0.00118f
C37648 control0.count\[1\] _1069_/a_193_47# 0.07856f
C37649 _1070_/a_891_413# clknet_1_0__leaf_clk 0
C37650 VPWR _1069_/a_381_47# 0.07969f
C37651 control0.state\[0\] _0160_ 0.0012f
C37652 _0982_/a_592_47# _0183_ 0
C37653 output53/a_27_47# hold53/a_285_47# 0
C37654 hold27/a_285_47# _0138_ 0.07166f
C37655 _0269_ _0846_/a_245_297# 0.00111f
C37656 comp0.B\[12\] _1045_/a_891_413# 0
C37657 _0695_/a_80_21# _0743_/a_240_47# 0
C37658 _1052_/a_891_413# _0987_/a_193_47# 0
C37659 clknet_0__0460_ _0460_ 0.16022f
C37660 _1011_/a_891_413# net97 0
C37661 VPWR net24 0.68706f
C37662 _1011_/a_193_47# net57 0.00471f
C37663 _0239_ _0352_ 0.10112f
C37664 _1000_/a_1059_315# _0614_/a_29_53# 0
C37665 net50 net109 0.00298f
C37666 _0195_ _1011_/a_27_47# 0
C37667 _0985_/a_891_413# _0186_ 0.00213f
C37668 _0728_/a_145_75# acc0.A\[29\] 0.00112f
C37669 _1055_/a_634_159# A[9] 0
C37670 net243 _0574_/a_109_47# 0
C37671 rst _0162_ 0.00166f
C37672 _1006_/a_634_159# _1006_/a_381_47# 0
C37673 pp[10] net4 0.0805f
C37674 clkload2/Y _0148_ 0.01634f
C37675 _0993_/a_466_413# _0807_/a_68_297# 0.01106f
C37676 net182 _1055_/a_27_47# 0
C37677 acc0.A\[1\] _1014_/a_634_159# 0
C37678 net206 _0580_/a_109_297# 0.0015f
C37679 _0891_/a_27_47# net87 0
C37680 net56 _0345_ 0.03012f
C37681 _1052_/a_193_47# A[5] 0
C37682 output59/a_27_47# _0710_/a_109_297# 0
C37683 _0984_/a_27_47# _0984_/a_891_413# 0.03206f
C37684 _0984_/a_193_47# _0984_/a_1059_315# 0.03405f
C37685 _0984_/a_634_159# _0984_/a_466_413# 0.23992f
C37686 _0352_ _1026_/a_466_413# 0
C37687 _0179_ _0178_ 0.13699f
C37688 net185 _1034_/a_891_413# 0
C37689 hold66/a_391_47# hold3/a_285_47# 0.00309f
C37690 hold66/a_285_47# hold3/a_391_47# 0.00309f
C37691 acc0.A\[22\] net49 0
C37692 _1003_/a_1017_47# VPWR 0
C37693 _0429_ _0436_ 0.2353f
C37694 _0442_ _0218_ 0.3677f
C37695 hold69/a_49_47# _0346_ 0.0388f
C37696 _1039_/a_466_413# VPWR 0.24035f
C37697 _0986_/a_634_159# _0986_/a_381_47# 0
C37698 net148 _0987_/a_975_413# 0
C37699 _0524_/a_27_297# _0085_ 0
C37700 _0524_/a_109_297# net73 0
C37701 _0300_ _0219_ 0
C37702 _0486_ _0161_ 0
C37703 _1017_/a_891_413# _0181_ 0.05134f
C37704 _1023_/a_634_159# _1023_/a_592_47# 0
C37705 clknet_0__0461_ _0247_ 0.01728f
C37706 clkbuf_1_0__f__0461_/a_110_47# _0240_ 0
C37707 _0616_/a_215_47# _1006_/a_27_47# 0
C37708 net1 clknet_1_0__leaf__0461_ 0.07429f
C37709 VPWR _0411_ 0.29397f
C37710 net36 comp0.B\[6\] 0.00848f
C37711 _0277_ _0669_/a_29_53# 0.14033f
C37712 hold101/a_285_47# _0432_ 0
C37713 _0405_ net6 0.02f
C37714 clknet_1_0__leaf__0463_ _0177_ 0
C37715 _1042_/a_891_413# _1042_/a_975_413# 0.00851f
C37716 _1042_/a_27_47# net128 0.22701f
C37717 _1042_/a_381_47# _1042_/a_561_413# 0.00123f
C37718 clknet_1_0__leaf__0458_ net67 0.0013f
C37719 _1019_/a_466_413# control0.add 0
C37720 _0181_ net146 0.20411f
C37721 A[5] net12 0.13075f
C37722 output67/a_27_47# acc0.A\[11\] 0
C37723 net34 net17 0
C37724 _1033_/a_27_47# _0163_ 0
C37725 net96 _0352_ 0
C37726 net50 pp[24] 0
C37727 _0731_/a_81_21# clkbuf_0__0460_/a_110_47# 0.00898f
C37728 _1011_/a_891_413# _0707_/a_201_297# 0
C37729 clknet_1_1__leaf__0464_ _1044_/a_381_47# 0.01548f
C37730 _1045_/a_27_47# _0142_ 0
C37731 _0832_/a_113_47# clknet_1_1__leaf__0458_ 0
C37732 hold68/a_391_47# acc0.A\[23\] 0.00151f
C37733 hold89/a_49_47# _0972_/a_93_21# 0
C37734 _1021_/a_381_47# net118 0
C37735 net225 _0339_ 0.00667f
C37736 _1036_/a_891_413# comp0.B\[4\] 0.00527f
C37737 _0466_ _1064_/a_891_413# 0
C37738 _0399_ _0826_/a_219_297# 0
C37739 _0254_ _0990_/a_193_47# 0
C37740 net10 _1042_/a_592_47# 0
C37741 hold16/a_285_47# _1031_/a_193_47# 0
C37742 hold16/a_49_47# _1031_/a_634_159# 0
C37743 hold16/a_391_47# _1031_/a_27_47# 0
C37744 net45 clknet_1_0__leaf__0457_ 0
C37745 _0229_ net213 0
C37746 _0153_ _0988_/a_975_413# 0
C37747 _0710_/a_109_47# _0195_ 0
C37748 net9 hold7/a_285_47# 0.02544f
C37749 _0343_ _0253_ 0.20847f
C37750 _0430_ _0369_ 0.02416f
C37751 _0808_/a_266_47# _0345_ 0
C37752 net165 _0848_/a_27_47# 0.00171f
C37753 _0621_/a_285_47# _0369_ 0
C37754 _0752_/a_27_413# net51 0.0136f
C37755 _0746_/a_384_47# _0462_ 0
C37756 pp[29] _1011_/a_1059_315# 0.00158f
C37757 _1057_/a_27_47# net192 0
C37758 _1038_/a_27_47# _1037_/a_193_47# 0
C37759 _1038_/a_193_47# _1037_/a_27_47# 0
C37760 _0399_ _0611_/a_68_297# 0
C37761 hold52/a_391_47# net215 0.00804f
C37762 _0975_/a_59_75# _0477_ 0
C37763 _0218_ net165 0.02622f
C37764 net101 _1020_/a_27_47# 0
C37765 _0997_/a_634_159# _0407_ 0
C37766 _0732_/a_80_21# net93 0
C37767 _0784_/a_113_47# _0369_ 0
C37768 _0401_ _0369_ 0.02455f
C37769 acc0.A\[5\] _0369_ 0
C37770 net87 _0346_ 0.02729f
C37771 _0315_ _0352_ 0
C37772 _0366_ _0102_ 0
C37773 _0179_ net63 0.01924f
C37774 _0790_/a_35_297# net41 0
C37775 _1002_/a_466_413# net220 0
C37776 _0777_/a_129_47# _0308_ 0
C37777 _0311_ _0393_ 0
C37778 hold85/a_391_47# _1066_/a_193_47# 0
C37779 net21 net9 0
C37780 net144 _0187_ 0
C37781 hold28/a_49_47# _0197_ 0.01794f
C37782 _0099_ hold40/a_391_47# 0
C37783 _0477_ net231 0.02163f
C37784 _0216_ acc0.A\[1\] 0
C37785 _0195_ _0180_ 0.2526f
C37786 _0662_/a_299_297# _0293_ 0.00863f
C37787 _0195_ net218 0.258f
C37788 hold19/a_391_47# _0114_ 0.0556f
C37789 acc0.A\[25\] _0321_ 0.01093f
C37790 clkload4/a_110_47# VPWR 0
C37791 net117 _0216_ 0.1053f
C37792 _0743_/a_149_47# _0345_ 0.00154f
C37793 _0115_ clknet_1_1__leaf__0461_ 0.1352f
C37794 _0218_ acc0.A\[19\] 0.22822f
C37795 hold30/a_285_47# net151 0
C37796 _0444_ _0431_ 0
C37797 _0195_ _1013_/a_193_47# 0.02837f
C37798 net33 comp0.B\[6\] 0
C37799 _0236_ _0749_/a_81_21# 0.23535f
C37800 _1058_/a_561_413# acc0.A\[11\] 0
C37801 _0457_ net201 0.00581f
C37802 _0280_ _0403_ 0
C37803 clknet_1_1__leaf__0459_ _0420_ 0.00189f
C37804 VPWR _1035_/a_381_47# 0.07736f
C37805 _1001_/a_1059_315# net45 0
C37806 net180 _1040_/a_193_47# 0.00181f
C37807 net30 _1040_/a_27_47# 0
C37808 _0183_ _0347_ 0.02275f
C37809 net150 _0352_ 0.25577f
C37810 VPWR input23/a_75_212# 0.27912f
C37811 _0274_ _0271_ 0.2182f
C37812 _0275_ _0256_ 0.00571f
C37813 _0404_ _0219_ 0
C37814 _0982_/a_891_413# _0181_ 0.05866f
C37815 _0754_/a_149_47# _0219_ 0.00242f
C37816 _0754_/a_240_47# net241 0.06201f
C37817 _0814_/a_27_47# _0345_ 0.00282f
C37818 VPWR _0809_/a_299_297# 0.28386f
C37819 net15 net75 0
C37820 _0179_ _1053_/a_891_413# 0
C37821 _0992_/a_1059_315# _0286_ 0
C37822 _0992_/a_891_413# _0283_ 0
C37823 _0207_ input29/a_75_212# 0
C37824 _0298_ _0669_/a_29_53# 0
C37825 _1055_/a_634_159# _0516_/a_27_297# 0
C37826 _1064_/a_634_159# _1064_/a_1059_315# 0
C37827 _1064_/a_27_47# _1064_/a_381_47# 0.05761f
C37828 _1064_/a_193_47# _1064_/a_891_413# 0.19421f
C37829 net179 clknet_1_1__leaf__0465_ 0.0858f
C37830 _0643_/a_337_297# _0431_ 0
C37831 _1018_/a_634_159# net149 0
C37832 _0837_/a_266_47# _0271_ 0
C37833 clknet_1_1__leaf__0460_ net51 0.00211f
C37834 clknet_0__0457_ _0182_ 0
C37835 clk _1068_/a_381_47# 0
C37836 clk net1 0
C37837 _1018_/a_891_413# _1017_/a_27_47# 0
C37838 _1018_/a_1059_315# _1017_/a_193_47# 0
C37839 net170 _0449_ 0
C37840 net45 _0588_/a_113_47# 0
C37841 _1047_/a_193_47# _0171_ 0
C37842 _0440_ _0987_/a_27_47# 0
C37843 _1026_/a_381_47# _1025_/a_27_47# 0
C37844 _1026_/a_27_47# _1025_/a_381_47# 0
C37845 _0712_/a_297_297# _0712_/a_465_47# 0
C37846 _0712_/a_79_21# _0712_/a_561_47# 0
C37847 clkload1/Y _0255_ 0
C37848 _0294_ _0250_ 0.0024f
C37849 _1051_/a_891_413# net148 0
C37850 _1051_/a_27_47# _0194_ 0
C37851 _0343_ _1017_/a_27_47# 0.00308f
C37852 _0607_/a_27_297# _0240_ 0
C37853 hold98/a_285_47# _0218_ 0
C37854 _1033_/a_891_413# comp0.B\[0\] 0.00438f
C37855 net132 _0142_ 0.17245f
C37856 _0845_/a_109_297# _0449_ 0
C37857 _0362_ clknet_1_1__leaf__0460_ 0.00562f
C37858 _0467_ net240 0
C37859 net1 _0585_/a_27_297# 0.17617f
C37860 _0852_/a_285_297# acc0.A\[1\] 0
C37861 hold53/a_285_47# net111 0
C37862 _0343_ _1060_/a_975_413# 0
C37863 _0324_ acc0.A\[26\] 0.00275f
C37864 _0974_/a_79_199# _0166_ 0.11939f
C37865 _0452_ _0465_ 0.00258f
C37866 _0170_ clknet_0_clk 0.06667f
C37867 _0348_ hold62/a_49_47# 0.00105f
C37868 _0373_ hold73/a_285_47# 0
C37869 _0946_/a_184_297# control0.state\[2\] 0
C37870 _0343_ net74 0.15445f
C37871 net114 _1027_/a_891_413# 0.00274f
C37872 _0627_/a_215_53# clkbuf_1_1__f__0458_/a_110_47# 0
C37873 _0553_/a_240_47# _0209_ 0
C37874 hold25/a_49_47# net8 0.05319f
C37875 _0346_ acc0.A\[6\] 0
C37876 _1010_/a_592_47# _0350_ 0.00164f
C37877 clknet_0__0458_ acc0.A\[8\] 0
C37878 _0737_/a_117_297# _0321_ 0.00183f
C37879 _0737_/a_285_297# _0360_ 0.06712f
C37880 hold16/a_49_47# _0345_ 0
C37881 _0854_/a_79_21# _0854_/a_215_47# 0.04584f
C37882 clknet_1_1__leaf__0464_ _1042_/a_193_47# 0
C37883 hold74/a_285_47# net103 0.00271f
C37884 _0697_/a_472_297# _0322_ 0
C37885 _0697_/a_217_297# _0329_ 0.00405f
C37886 _0601_/a_68_297# clknet_1_0__leaf__0460_ 0.00669f
C37887 hold39/a_49_47# _0176_ 0
C37888 _0961_/a_113_297# clk 0
C37889 _0347_ acc0.A\[15\] 0.03457f
C37890 net65 acc0.A\[6\] 0.00732f
C37891 net157 _1061_/a_592_47# 0
C37892 _0331_ _0322_ 0
C37893 _0217_ _0574_/a_27_297# 0.12214f
C37894 _0989_/a_466_413# acc0.A\[6\] 0
C37895 _0305_ _1016_/a_193_47# 0
C37896 _0800_/a_51_297# _0997_/a_1059_315# 0
C37897 _0800_/a_240_47# _0997_/a_27_47# 0
C37898 hold36/a_285_47# _0201_ 0
C37899 _0830_/a_79_21# _0830_/a_510_47# 0.00844f
C37900 _0830_/a_297_297# _0830_/a_215_47# 0
C37901 _0331_ _0327_ 0
C37902 _0179_ _0812_/a_79_21# 0.02154f
C37903 comp0.B\[4\] _0474_ 0.04649f
C37904 _0695_/a_300_47# _0327_ 0
C37905 clkbuf_1_1__f__0465_/a_110_47# _0992_/a_193_47# 0
C37906 _0174_ net18 0.5203f
C37907 acc0.A\[1\] net247 0.34684f
C37908 _0343_ output61/a_27_47# 0.00377f
C37909 clknet_1_0__leaf__0465_ _1052_/a_193_47# 0.00631f
C37910 _0251_ _0829_/a_109_297# 0
C37911 _0475_ net201 0
C37912 input33/a_75_212# init 0.20079f
C37913 _1037_/a_466_413# VPWR 0.25751f
C37914 _0837_/a_368_297# acc0.A\[4\] 0
C37915 _0183_ _1016_/a_891_413# 0
C37916 _0228_ _0219_ 0.12029f
C37917 clkbuf_1_1__f_clk/a_110_47# clknet_1_0__leaf__0457_ 0.06584f
C37918 _1031_/a_891_413# _1031_/a_1017_47# 0.00617f
C37919 net175 _1047_/a_634_159# 0
C37920 _0289_ _0786_/a_300_47# 0
C37921 hold30/a_285_47# _0378_ 0.01284f
C37922 net23 _0566_/a_27_47# 0
C37923 _0733_/a_222_93# _0324_ 0.00268f
C37924 _1041_/a_381_47# VPWR 0.07133f
C37925 _0457_ comp0.B\[2\] 0
C37926 _1022_/a_27_47# _1005_/a_1059_315# 0
C37927 pp[15] _0995_/a_891_413# 0.00232f
C37928 _0722_/a_215_47# _0351_ 0.01166f
C37929 _0722_/a_79_21# _0110_ 0.05051f
C37930 _1005_/a_592_47# _0103_ 0.00188f
C37931 _0983_/a_27_47# clknet_1_0__leaf__0461_ 0
C37932 _0229_ _0603_/a_68_297# 0
C37933 net17 _0565_/a_512_297# 0
C37934 control0.add _0352_ 0.07687f
C37935 _0260_ _0529_/a_109_297# 0
C37936 _0742_/a_81_21# _0352_ 0.01772f
C37937 _0438_ _0831_/a_117_297# 0
C37938 _0326_ _0367_ 0
C37939 clkbuf_1_1__f__0465_/a_110_47# _0427_ 0.00423f
C37940 _1066_/a_193_47# _0160_ 0
C37941 clknet_1_1__leaf_clk _1062_/a_634_159# 0.01165f
C37942 _1056_/a_634_159# pp[9] 0
C37943 _0082_ _0506_/a_299_297# 0
C37944 _1060_/a_891_413# _0185_ 0.01331f
C37945 _0158_ _0507_/a_109_47# 0
C37946 _1021_/a_27_47# clknet_1_1__leaf_clk 0
C37947 _1054_/a_1059_315# clknet_1_1__leaf__0458_ 0.07873f
C37948 _0254_ _0438_ 0.03659f
C37949 _1002_/a_466_413# net88 0.00992f
C37950 _1020_/a_193_47# _1020_/a_634_159# 0.11897f
C37951 _1020_/a_27_47# _1020_/a_466_413# 0.27314f
C37952 _1002_/a_634_159# _0100_ 0.04448f
C37953 _0792_/a_209_47# net42 0
C37954 _0405_ _0790_/a_285_297# 0.00134f
C37955 _0182_ _0844_/a_79_21# 0
C37956 _1027_/a_466_413# _0106_ 0
C37957 clknet_1_0__leaf__0465_ net12 0.12378f
C37958 _0269_ _0448_ 0.0183f
C37959 net156 _0347_ 0
C37960 net63 _0441_ 0
C37961 net45 hold19/a_285_47# 0
C37962 _0363_ _0746_/a_299_297# 0
C37963 _0598_/a_79_21# _0752_/a_27_413# 0
C37964 _0820_/a_215_47# _0820_/a_510_47# 0.00529f
C37965 _0310_ _0392_ 0.04077f
C37966 _0680_/a_80_21# _0326_ 0
C37967 _0983_/a_193_47# net47 0.05484f
C37968 _1016_/a_27_47# net43 0
C37969 acc0.A\[22\] _0757_/a_68_297# 0
C37970 _1058_/a_634_159# clknet_1_1__leaf__0465_ 0
C37971 _0309_ _0352_ 0.00138f
C37972 _1059_/a_1017_47# _0369_ 0
C37973 _0217_ net105 0.01325f
C37974 _0180_ _1048_/a_193_47# 0.02678f
C37975 _0182_ _1048_/a_634_159# 0
C37976 _0998_/a_193_47# _1017_/a_27_47# 0
C37977 _0998_/a_27_47# _1017_/a_193_47# 0
C37978 clkbuf_1_0__f__0459_/a_110_47# net221 0
C37979 _1001_/a_466_413# net46 0
C37980 _0179_ _0347_ 0.0491f
C37981 control0.state\[1\] _0477_ 0.12076f
C37982 _0440_ _0191_ 0
C37983 _0284_ clknet_1_1__leaf__0459_ 0.14397f
C37984 _0222_ _0762_/a_215_47# 0
C37985 net220 _0385_ 0.29589f
C37986 hold88/a_285_47# _0181_ 0
C37987 _1003_/a_193_47# _0466_ 0
C37988 clkload4/a_110_47# clknet_1_0__leaf__0459_ 0
C37989 net64 clknet_0__0458_ 0.047f
C37990 pp[28] _1011_/a_975_413# 0
C37991 _0233_ net51 0.16744f
C37992 net67 _0288_ 0.24227f
C37993 control0.sh _1047_/a_27_47# 0
C37994 output44/a_27_47# _0220_ 0.0089f
C37995 _0181_ _0487_ 0.20771f
C37996 _0216_ _0223_ 0
C37997 _1036_/a_27_47# net24 0
C37998 _0230_ _0618_/a_79_21# 0
C37999 net86 _0775_/a_79_21# 0.01476f
C38000 _1000_/a_891_413# _0393_ 0
C38001 _0413_ _0799_/a_209_47# 0
C38002 pp[11] net246 0.00538f
C38003 _0800_/a_149_47# _0411_ 0
C38004 _0343_ net238 0.00558f
C38005 comp0.B\[12\] _1044_/a_1059_315# 0.08445f
C38006 net178 acc0.A\[8\] 0.00495f
C38007 _1066_/a_466_413# net17 0
C38008 _0269_ _0444_ 0
C38009 hold10/a_391_47# _0464_ 0.00215f
C38010 _0924_/a_27_47# _1061_/a_1059_315# 0
C38011 _0967_/a_297_297# control0.state\[2\] 0.00108f
C38012 control0.state\[2\] _0162_ 0.0037f
C38013 VPWR control0.count\[0\] 1.91463f
C38014 clknet_1_0__leaf__0462_ _0682_/a_68_297# 0.00102f
C38015 A[0] B[0] 0.11881f
C38016 comp0.B\[2\] _0475_ 0.06885f
C38017 hold57/a_285_47# _0176_ 0.03688f
C38018 _0606_/a_109_53# _0374_ 0.02076f
C38019 hold67/a_49_47# net143 0
C38020 _0414_ _0994_/a_1059_315# 0
C38021 _0990_/a_891_413# _0186_ 0
C38022 _0121_ net110 0
C38023 _1052_/a_1059_315# net73 0
C38024 _1017_/a_891_413# clknet_1_1__leaf__0461_ 0.00162f
C38025 _1000_/a_975_413# _0245_ 0
C38026 _0572_/a_27_297# _0195_ 0.14411f
C38027 _0572_/a_109_297# net210 0.00954f
C38028 net141 A[9] 0.00163f
C38029 _1006_/a_381_47# net92 0
C38030 VPWR _0974_/a_544_297# 0.01188f
C38031 _0993_/a_592_47# net246 0
C38032 acc0.A\[1\] net100 0
C38033 net33 net26 0
C38034 VPWR clknet_1_0__leaf__0457_ 3.10839f
C38035 _0286_ _0809_/a_81_21# 0
C38036 _0655_/a_215_53# _0420_ 0.03807f
C38037 _0283_ _0809_/a_299_297# 0
C38038 acc0.A\[14\] hold82/a_285_47# 0
C38039 pp[30] _0340_ 0.00106f
C38040 _0323_ _0219_ 0.03594f
C38041 net21 net129 0
C38042 _0984_/a_466_413# net70 0
C38043 _0643_/a_337_297# _0269_ 0.01086f
C38044 _0573_/a_27_47# _0180_ 0.00797f
C38045 _0347_ acc0.A\[26\] 0.4255f
C38046 _0579_/a_27_297# _0461_ 0.00873f
C38047 clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk 1.78575f
C38048 _0714_/a_51_297# _0999_/a_193_47# 0
C38049 acc0.A\[19\] _0099_ 0
C38050 _0242_ _0391_ 0.02175f
C38051 _0305_ net41 0
C38052 net122 B[5] 0
C38053 _0102_ acc0.A\[24\] 0
C38054 _0285_ _0289_ 0
C38055 _0206_ _0204_ 0
C38056 net180 _0207_ 0.16033f
C38057 VPWR _0988_/a_1059_315# 0.41589f
C38058 VPWR _0553_/a_51_297# 0.47582f
C38059 _1015_/a_466_413# clknet_1_0__leaf__0457_ 0
C38060 clkbuf_1_1__f__0461_/a_110_47# _0218_ 0.14338f
C38061 _0344_ _1031_/a_466_413# 0.00203f
C38062 _1054_/a_27_47# _0186_ 0
C38063 output37/a_27_47# VPWR 0.39009f
C38064 net168 _1054_/a_381_47# 0.01459f
C38065 _0791_/a_113_297# _0345_ 0.00123f
C38066 VPWR _0953_/a_304_297# 0.00456f
C38067 _0194_ _0085_ 0
C38068 clkbuf_1_1__f__0465_/a_110_47# net142 0
C38069 _1056_/a_891_413# _0186_ 0.03281f
C38070 net157 _1047_/a_27_47# 0.02869f
C38071 _0274_ clknet_1_0__leaf__0465_ 0
C38072 hold89/a_49_47# _0975_/a_59_75# 0
C38073 _1023_/a_891_413# acc0.A\[23\] 0.00349f
C38074 comp0.B\[10\] _1043_/a_193_47# 0
C38075 _0585_/a_109_297# _0171_ 0
C38076 _0426_ _0218_ 0.06031f
C38077 _1037_/a_975_413# _0175_ 0
C38078 _1016_/a_193_47# _0181_ 0
C38079 _0581_/a_27_297# _0242_ 0
C38080 _0476_ hold38/a_49_47# 0
C38081 _1044_/a_634_159# net20 0.01938f
C38082 hold64/a_285_47# acc0.A\[1\] 0
C38083 _0670_/a_79_21# _0670_/a_297_297# 0.01735f
C38084 _0466_ _0471_ 0.00481f
C38085 _0768_/a_27_47# _0392_ 0.00396f
C38086 _0101_ clknet_0_clk 0
C38087 _0404_ _0799_/a_209_297# 0.02807f
C38088 _0298_ _0799_/a_80_21# 0.04082f
C38089 _0216_ _0571_/a_373_47# 0.00103f
C38090 _0457_ _1015_/a_193_47# 0.03751f
C38091 net57 _0707_/a_75_199# 0.05647f
C38092 _0538_/a_240_47# _0172_ 0.02765f
C38093 net184 net20 0
C38094 _0402_ _0806_/a_113_297# 0.10773f
C38095 _1037_/a_592_47# control0.sh 0
C38096 VPWR _0635_/a_27_47# 0.00625f
C38097 _0349_ hold62/a_285_47# 0.00266f
C38098 hold22/a_285_47# net11 0
C38099 pp[28] _0334_ 0.09325f
C38100 _0757_/a_68_297# _0379_ 0.04127f
C38101 _0350_ _0756_/a_285_47# 0
C38102 _1037_/a_27_47# net29 0
C38103 _1037_/a_193_47# B[6] 0
C38104 net48 clknet_1_0__leaf__0457_ 0.00217f
C38105 _1001_/a_1059_315# VPWR 0.39724f
C38106 hold27/a_285_47# net22 0.00228f
C38107 net163 _1031_/a_381_47# 0.12224f
C38108 _0627_/a_215_53# _0291_ 0
C38109 hold36/a_49_47# clknet_0__0464_ 0.02728f
C38110 _0129_ _1031_/a_975_413# 0.00101f
C38111 _0159_ _0176_ 0
C38112 net45 _1017_/a_634_159# 0.0044f
C38113 VPWR _1062_/a_466_413# 0.25485f
C38114 _0504_/a_27_47# _0265_ 0
C38115 _0616_/a_78_199# _0240_ 0.00316f
C38116 _0616_/a_215_47# _0247_ 0.01275f
C38117 net64 net178 0.68609f
C38118 _0157_ _0506_/a_81_21# 0
C38119 net145 _0506_/a_299_297# 0.00821f
C38120 _0780_/a_35_297# _0347_ 0.00768f
C38121 _0181_ clkbuf_0__0457_/a_110_47# 0
C38122 _1039_/a_27_47# _0137_ 0.09079f
C38123 _1039_/a_1059_315# net180 0
C38124 _1039_/a_634_159# _0172_ 0
C38125 _1021_/a_193_47# VPWR 0.31734f
C38126 VPWR hold90/a_391_47# 0.16377f
C38127 _0369_ _0616_/a_78_199# 0
C38128 output57/a_27_47# _0216_ 0
C38129 _1018_/a_891_413# _0245_ 0
C38130 comp0.B\[13\] net18 0
C38131 clkbuf_1_0__f__0457_/a_110_47# _0616_/a_215_47# 0
C38132 _0762_/a_79_21# _0762_/a_510_47# 0.00844f
C38133 _0762_/a_297_297# _0762_/a_215_47# 0
C38134 hold52/a_49_47# hold52/a_391_47# 0.00188f
C38135 hold20/a_391_47# _1068_/a_891_413# 0
C38136 _0574_/a_109_47# acc0.A\[24\] 0.00267f
C38137 _0456_ _0265_ 0.00318f
C38138 _0343_ _0245_ 0.62079f
C38139 _0776_/a_109_297# _0308_ 0.01155f
C38140 VPWR _0588_/a_113_47# 0
C38141 _0260_ net170 0.00287f
C38142 _0437_ _0619_/a_150_297# 0
C38143 _0440_ clkbuf_1_0__f__0465_/a_110_47# 0.0039f
C38144 _0389_ _0719_/a_27_47# 0
C38145 output37/a_27_47# input4/a_75_212# 0.01973f
C38146 clknet_1_0__leaf__0463_ hold27/a_285_47# 0.00992f
C38147 _0197_ clkbuf_1_0__f__0464_/a_110_47# 0.00241f
C38148 _0606_/a_215_297# clkbuf_1_0__f__0460_/a_110_47# 0
C38149 _0390_ clknet_1_0__leaf__0457_ 0.00506f
C38150 _0100_ net220 0
C38151 VPWR _0561_/a_149_47# 0.00124f
C38152 _1065_/a_634_159# _1065_/a_381_47# 0
C38153 net150 _0237_ 0.04874f
C38154 _0217_ _0381_ 0.02736f
C38155 hold85/a_285_47# clknet_1_1__leaf_clk 0.01431f
C38156 _0998_/a_1059_315# _0218_ 0
C38157 _1036_/a_1059_315# _1035_/a_634_159# 0.00213f
C38158 _1036_/a_27_47# _1035_/a_381_47# 0
C38159 _1036_/a_891_413# _1035_/a_193_47# 0
C38160 net157 clknet_1_0__leaf__0461_ 0.13892f
C38161 clkbuf_1_1__f__0463_/a_110_47# comp0.B\[15\] 0
C38162 _1036_/a_27_47# input23/a_75_212# 0
C38163 _0853_/a_150_297# _0399_ 0
C38164 _1068_/a_27_47# _0484_ 0
C38165 control0.state\[0\] _0482_ 0.0015f
C38166 clknet_1_1__leaf__0458_ pp[4] 0
C38167 _0985_/a_1059_315# _0270_ 0
C38168 net237 _0219_ 0.15366f
C38169 comp0.B\[11\] _1042_/a_27_47# 0.07257f
C38170 _0266_ _0633_/a_109_297# 0
C38171 _1014_/a_27_47# _1014_/a_1059_315# 0.04875f
C38172 _1014_/a_193_47# _1014_/a_466_413# 0.07482f
C38173 net33 hold84/a_285_47# 0.03898f
C38174 net152 _0540_/a_240_47# 0
C38175 hold52/a_285_47# net52 0
C38176 control0.count\[2\] clknet_1_0__leaf_clk 0.25952f
C38177 VPWR _1047_/a_891_413# 0.19606f
C38178 clknet_1_1__leaf__0460_ _0324_ 0.31157f
C38179 _0716_/a_27_47# net228 0
C38180 output67/a_27_47# A[12] 0.07394f
C38181 _0647_/a_47_47# pp[12] 0
C38182 A[13] net5 0.00913f
C38183 _1052_/a_27_47# _0149_ 0
C38184 VPWR _1007_/a_975_413# 0.00535f
C38185 _0340_ _0339_ 0.27927f
C38186 hold34/a_391_47# A[11] 0
C38187 net133 control0.sh 0
C38188 _0312_ _0746_/a_384_47# 0
C38189 _1021_/a_193_47# net48 0
C38190 _0734_/a_129_47# VPWR 0
C38191 hold87/a_49_47# _0217_ 0
C38192 VPWR _0850_/a_68_297# 0.15153f
C38193 _0178_ _1049_/a_891_413# 0
C38194 output56/a_27_47# _1010_/a_27_47# 0
C38195 _1039_/a_27_47# comp0.B\[6\] 0
C38196 _0280_ acc0.A\[13\] 0
C38197 _1055_/a_1059_315# net16 0.01741f
C38198 _1055_/a_634_159# _0190_ 0
C38199 net55 _0317_ 0.08322f
C38200 clknet_1_1__leaf__0465_ _1060_/a_634_159# 0.00197f
C38201 net104 net149 0
C38202 hold78/a_391_47# _0219_ 0
C38203 _0830_/a_79_21# _0989_/a_193_47# 0
C38204 clkbuf_1_0__f__0459_/a_110_47# _1017_/a_27_47# 0
C38205 _0956_/a_32_297# comp0.B\[0\] 0.14415f
C38206 _1000_/a_891_413# net206 0
C38207 _0304_ _0301_ 0
C38208 _0615_/a_109_297# _0393_ 0
C38209 _0341_ output60/a_27_47# 0
C38210 net112 _1025_/a_1059_315# 0
C38211 _1026_/a_27_47# acc0.A\[25\] 0.08688f
C38212 hold78/a_49_47# hold78/a_285_47# 0.22264f
C38213 _0390_ _1001_/a_1059_315# 0
C38214 _0088_ _0988_/a_891_413# 0
C38215 net137 net12 0
C38216 VPWR _0748_/a_299_297# 0.26277f
C38217 _0585_/a_27_297# control0.sh 0
C38218 clknet_0_clk net23 0
C38219 _0151_ hold83/a_391_47# 0.03387f
C38220 _1025_/a_1059_315# acc0.A\[24\] 0.01754f
C38221 _0183_ _1059_/a_27_47# 0
C38222 clknet_1_0__leaf__0462_ _0753_/a_561_47# 0
C38223 net1 _0112_ 0.04624f
C38224 hold41/a_49_47# net3 0.01205f
C38225 _0693_/a_150_297# _0460_ 0
C38226 clknet_1_0__leaf__0459_ clknet_1_0__leaf__0457_ 0.02728f
C38227 control0.state\[0\] _0476_ 0.24702f
C38228 net120 _1032_/a_27_47# 0
C38229 output42/a_27_47# pp[15] 0.1682f
C38230 _0985_/a_1059_315# net233 0
C38231 _0985_/a_381_47# net61 0
C38232 net25 _1066_/a_634_159# 0
C38233 hold49/a_285_47# VPWR 0.35626f
C38234 _0981_/a_27_297# _0981_/a_373_47# 0.01338f
C38235 _0285_ _0418_ 0.12356f
C38236 _0686_/a_27_53# _0219_ 0
C38237 _1042_/a_27_47# _0202_ 0
C38238 _0216_ _0704_/a_68_297# 0.01048f
C38239 net106 control0.add 0
C38240 pp[27] _0216_ 0.12562f
C38241 _0222_ _1022_/a_1059_315# 0.04712f
C38242 net163 _0219_ 0
C38243 _0481_ _1070_/a_634_159# 0
C38244 VPWR hold19/a_285_47# 0.28061f
C38245 _0854_/a_510_47# _0081_ 0
C38246 _1037_/a_634_159# _1036_/a_193_47# 0
C38247 _1037_/a_27_47# _1036_/a_466_413# 0
C38248 _1037_/a_466_413# _1036_/a_27_47# 0
C38249 _0343_ net61 0.04223f
C38250 _0500_/a_27_47# hold71/a_285_47# 0
C38251 _0313_ clkbuf_1_1__f__0460_/a_110_47# 0
C38252 _0642_/a_27_413# _0436_ 0
C38253 _0642_/a_215_297# _0435_ 0
C38254 _0836_/a_68_297# net212 0
C38255 _0140_ net153 0.00578f
C38256 _0600_/a_337_297# _0366_ 0
C38257 _0817_/a_81_21# _0401_ 0.002f
C38258 net203 clkbuf_1_1__f__0463_/a_110_47# 0.02033f
C38259 _0625_/a_59_75# _0438_ 0
C38260 _0297_ _0668_/a_382_297# 0
C38261 _0234_ _0373_ 0
C38262 _0999_/a_466_413# _0352_ 0.01173f
C38263 _0983_/a_193_47# _0294_ 0
C38264 _0983_/a_27_47# _0218_ 0
C38265 hold78/a_285_47# _0129_ 0
C38266 _0344_ hold16/a_285_47# 0
C38267 _1013_/a_27_47# pp[31] 0
C38268 _0498_/a_149_47# _0498_/a_240_47# 0.06872f
C38269 _0958_/a_27_47# clknet_1_1__leaf_clk 0
C38270 net35 clknet_0_clk 0.10832f
C38271 _0640_/a_297_297# _0255_ 0.00473f
C38272 _0820_/a_79_21# _0428_ 0.13512f
C38273 pp[8] hold35/a_285_47# 0
C38274 _0730_/a_79_21# acc0.A\[29\] 0
C38275 net133 net157 0.0029f
C38276 _0467_ hold56/a_285_47# 0
C38277 _0179_ net2 0.22436f
C38278 _0275_ clknet_0__0465_ 0.2036f
C38279 _1038_/a_193_47# _0174_ 0
C38280 comp0.B\[2\] _1033_/a_193_47# 0.04134f
C38281 _0135_ VPWR 0.30989f
C38282 net36 _1040_/a_466_413# 0
C38283 net150 _1005_/a_27_47# 0.03717f
C38284 net190 _1028_/a_193_47# 0.35592f
C38285 _0195_ _1014_/a_1059_315# 0
C38286 _0216_ _1014_/a_634_159# 0
C38287 output56/a_27_47# pp[30] 0
C38288 A[11] _0181_ 0.00219f
C38289 _0289_ _0218_ 0
C38290 output67/a_27_47# _1057_/a_193_47# 0
C38291 _0992_/a_27_47# _0417_ 0
C38292 hold33/a_285_47# _0176_ 0
C38293 _0735_/a_109_297# _0328_ 0
C38294 _0845_/a_193_297# _0447_ 0.00571f
C38295 _0272_ _0350_ 0
C38296 clknet_1_0__leaf__0458_ _0447_ 0
C38297 net44 _0775_/a_79_21# 0
C38298 net43 _0400_ 0
C38299 _0977_/a_75_212# _0466_ 0
C38300 _0837_/a_585_47# clknet_0__0465_ 0
C38301 _0972_/a_250_297# _0468_ 0.00603f
C38302 net46 _0241_ 0.37564f
C38303 _0413_ _0668_/a_79_21# 0
C38304 _1003_/a_27_47# clknet_1_0__leaf__0460_ 0.05626f
C38305 control0.state\[1\] hold89/a_49_47# 0.05765f
C38306 clkbuf_0__0462_/a_110_47# hold90/a_49_47# 0.01853f
C38307 control0.state\[0\] hold89/a_285_47# 0.00421f
C38308 net1 net240 0
C38309 _1048_/a_381_47# _0148_ 0
C38310 _1048_/a_592_47# _0196_ 0
C38311 _1059_/a_27_47# acc0.A\[15\] 0.01034f
C38312 _0384_ _0369_ 0.00178f
C38313 _0504_/a_27_47# _0267_ 0
C38314 _1001_/a_1059_315# clknet_1_0__leaf__0459_ 0
C38315 _1018_/a_1059_315# net219 0.01018f
C38316 _1018_/a_634_159# net206 0.02818f
C38317 _0585_/a_27_297# net157 0.00103f
C38318 net149 _0584_/a_27_297# 0
C38319 _0551_/a_27_47# clknet_1_1__leaf__0457_ 0
C38320 _0319_ _0365_ 0
C38321 net31 input7/a_75_212# 0.00391f
C38322 _1008_/a_193_47# _1008_/a_381_47# 0.09503f
C38323 _1008_/a_634_159# _1008_/a_891_413# 0.03684f
C38324 _1008_/a_27_47# _1008_/a_561_413# 0.0027f
C38325 _0488_ _1069_/a_592_47# 0
C38326 _0976_/a_535_374# control0.count\[0\] 0.0065f
C38327 _0401_ _0084_ 0
C38328 hold56/a_285_47# comp0.B\[0\] 0.00308f
C38329 _0648_/a_27_297# VPWR 0.22284f
C38330 _0718_/a_47_47# _1011_/a_891_413# 0
C38331 output43/a_27_47# _0995_/a_466_413# 0
C38332 _1020_/a_1059_315# _1020_/a_1017_47# 0
C38333 _1020_/a_27_47# _0118_ 0.0965f
C38334 net88 _0100_ 0.16249f
C38335 output53/a_27_47# _1025_/a_1059_315# 0
C38336 net53 _1025_/a_193_47# 0.04094f
C38337 _0408_ _0406_ 0.1623f
C38338 _0744_/a_27_47# _0181_ 0
C38339 _1035_/a_1059_315# comp0.B\[5\] 0.03133f
C38340 _0559_/a_51_297# _0561_/a_240_47# 0
C38341 _1035_/a_381_47# comp0.B\[3\] 0
C38342 _0559_/a_240_47# _0561_/a_51_297# 0
C38343 _0305_ _0350_ 0
C38344 _0175_ _0173_ 0.68822f
C38345 _0349_ _0350_ 0.14917f
C38346 _0255_ hold7/a_285_47# 0
C38347 net59 _0195_ 0
C38348 _0483_ clk 0
C38349 _0770_/a_297_47# _0218_ 0
C38350 _0371_ clkbuf_1_0__f__0460_/a_110_47# 0
C38351 hold28/a_391_47# acc0.A\[3\] 0.05005f
C38352 hold85/a_391_47# VPWR 0.18776f
C38353 clknet_0__0458_ _0986_/a_466_413# 0.00221f
C38354 _0316_ clknet_1_1__leaf__0460_ 0.18428f
C38355 _0217_ clknet_0__0461_ 0.01237f
C38356 clknet_0__0457_ _1014_/a_466_413# 0.00252f
C38357 _0515_/a_81_21# net181 0.10257f
C38358 net144 clknet_1_1__leaf__0465_ 0.27443f
C38359 hold34/a_391_47# net66 0.01841f
C38360 _0371_ _0250_ 0.38292f
C38361 _1054_/a_634_159# _0518_/a_27_297# 0
C38362 _0525_/a_81_21# _0524_/a_27_297# 0.01145f
C38363 net46 _0772_/a_510_47# 0.00114f
C38364 _0386_ _0766_/a_109_297# 0.01129f
C38365 _1032_/a_193_47# comp0.B\[0\] 0
C38366 _1041_/a_891_413# _0172_ 0.00631f
C38367 _0298_ _0997_/a_1059_315# 0
C38368 _0997_/a_193_47# _0345_ 0.02662f
C38369 acc0.A\[14\] _0671_/a_113_297# 0
C38370 clknet_1_1__leaf__0460_ _0347_ 0.22897f
C38371 _1004_/a_27_47# _0758_/a_79_21# 0.00189f
C38372 _0846_/a_51_297# _0449_ 0.11686f
C38373 _0992_/a_891_413# _0345_ 0
C38374 _0533_/a_27_297# clknet_1_1__leaf__0457_ 0.02281f
C38375 output39/a_27_47# VPWR 0.2838f
C38376 hold94/a_391_47# _0345_ 0.00376f
C38377 _0216_ _0724_/a_199_47# 0
C38378 hold21/a_391_47# A[8] 0.07266f
C38379 _0991_/a_1059_315# acc0.A\[15\] 0
C38380 _0346_ hold2/a_391_47# 0
C38381 _0176_ net20 0.0274f
C38382 clkbuf_1_0__f__0459_/a_110_47# net238 0
C38383 net66 _0510_/a_27_297# 0
C38384 _0734_/a_47_47# clkbuf_0__0462_/a_110_47# 0
C38385 hold48/a_285_47# _0176_ 0
C38386 _0982_/a_193_47# net234 0
C38387 _0982_/a_891_413# _0855_/a_299_297# 0
C38388 net102 _0582_/a_109_297# 0
C38389 net185 _0215_ 0
C38390 hold42/a_391_47# _1058_/a_466_413# 0
C38391 _0578_/a_27_297# _0183_ 0.19501f
C38392 _0578_/a_109_47# _0217_ 0.00371f
C38393 _0578_/a_373_47# net150 0.00122f
C38394 clknet_1_1__leaf__0460_ _0104_ 0
C38395 pp[9] hold35/a_49_47# 0
C38396 clk control0.count\[1\] 0.00149f
C38397 VPWR _0497_/a_150_297# 0.00129f
C38398 clknet_1_0__leaf__0458_ acc0.A\[0\] 0.00891f
C38399 _0166_ net17 0
C38400 _0179_ _1059_/a_27_47# 0.01332f
C38401 VPWR _0499_/a_59_75# 0.20939f
C38402 _0238_ _0374_ 0
C38403 _0576_/a_373_47# clknet_1_0__leaf__0460_ 0
C38404 _0701_/a_209_297# _0350_ 0.00609f
C38405 _0218_ acc0.A\[3\] 0
C38406 net45 _0246_ 0
C38407 _0198_ net247 0
C38408 _0195_ _0124_ 0.06588f
C38409 hold13/a_391_47# VPWR 0.1777f
C38410 _1016_/a_193_47# clknet_1_1__leaf__0461_ 0.45314f
C38411 clknet_1_1__leaf__0458_ net13 0
C38412 _0580_/a_109_47# _0264_ 0
C38413 _0247_ _0771_/a_215_297# 0
C38414 _0679_/a_68_297# _0240_ 0
C38415 VPWR _1017_/a_634_159# 0.17862f
C38416 acc0.A\[26\] _0106_ 0
C38417 _0679_/a_68_297# _0369_ 0
C38418 _1037_/a_193_47# comp0.B\[5\] 0
C38419 _0443_ _0084_ 0
C38420 _1037_/a_27_47# comp0.B\[6\] 0
C38421 _0415_ clknet_1_1__leaf__0459_ 0
C38422 _0172_ net147 0.22654f
C38423 _0378_ _1005_/a_193_47# 0
C38424 clknet_1_1__leaf__0460_ _0745_/a_109_47# 0
C38425 net70 _0506_/a_81_21# 0
C38426 _0563_/a_51_297# _0563_/a_245_297# 0.01218f
C38427 VPWR _1060_/a_1017_47# 0
C38428 _0346_ _0826_/a_219_297# 0
C38429 output56/a_27_47# _0339_ 0.00892f
C38430 _0804_/a_79_21# VPWR 0.49222f
C38431 _1017_/a_27_47# clkbuf_0__0461_/a_110_47# 0.00199f
C38432 _0399_ _0869_/a_27_47# 0
C38433 clknet_0_clk _1063_/a_466_413# 0
C38434 _1044_/a_27_47# net19 0
C38435 _0113_ clknet_1_0__leaf__0457_ 0
C38436 _0178_ _0171_ 0.18051f
C38437 net66 _0181_ 0.27902f
C38438 _0157_ _0184_ 0
C38439 _1000_/a_381_47# _0774_/a_68_297# 0
C38440 VPWR _1050_/a_466_413# 0.2483f
C38441 clknet_1_0__leaf__0459_ hold19/a_285_47# 0.06323f
C38442 clkbuf_0__0458_/a_110_47# _0448_ 0
C38443 _0453_ _0850_/a_68_297# 0.01341f
C38444 _0311_ _0387_ 0
C38445 hold45/a_391_47# net192 0.16272f
C38446 pp[9] A[9] 0.17253f
C38447 _0252_ _0619_/a_150_297# 0
C38448 hold45/a_49_47# _0156_ 0
C38449 _1010_/a_27_47# _1010_/a_466_413# 0.27314f
C38450 _1010_/a_193_47# _1010_/a_634_159# 0.11072f
C38451 _0179_ _0991_/a_1059_315# 0
C38452 _0116_ _0242_ 0
C38453 clknet_1_0__leaf__0462_ _1004_/a_27_47# 0.01813f
C38454 _0644_/a_129_47# net42 0.00232f
C38455 _0217_ _0468_ 0
C38456 _0670_/a_215_47# _0302_ 0
C38457 _0991_/a_27_47# _0181_ 0.03663f
C38458 pp[27] _1010_/a_561_413# 0
C38459 hold36/a_49_47# hold47/a_285_47# 0
C38460 _0183_ net218 0
C38461 _0541_/a_68_297# _0541_/a_150_297# 0.00477f
C38462 net57 _0338_ 0.0347f
C38463 _0146_ _1048_/a_27_47# 0.10163f
C38464 _0198_ _1048_/a_466_413# 0
C38465 _0195_ _0335_ 0
C38466 _0713_/a_27_47# _0457_ 0.004f
C38467 _0536_/a_149_47# net157 0.00957f
C38468 VPWR _0973_/a_109_47# 0
C38469 hold96/a_391_47# _0216_ 0.06455f
C38470 _0218_ _0418_ 0
C38471 _1002_/a_193_47# _0217_ 0.0238f
C38472 _0473_ _0913_/a_27_47# 0.00125f
C38473 _0238_ acc0.A\[19\] 0.00349f
C38474 _0746_/a_299_297# _0746_/a_384_47# 0
C38475 hold88/a_391_47# _0990_/a_27_47# 0
C38476 _0376_ _0606_/a_465_297# 0
C38477 net45 net103 0.00632f
C38478 _0482_ _0478_ 0.11091f
C38479 _1020_/a_1059_315# _0461_ 0
C38480 VPWR _0160_ 0.94136f
C38481 net125 _0172_ 0.12547f
C38482 net191 hold50/a_285_47# 0
C38483 _0137_ _0953_/a_32_297# 0
C38484 _0369_ _0383_ 0.0394f
C38485 _0481_ _0479_ 0
C38486 hold91/a_285_47# net6 0
C38487 clkbuf_0__0458_/a_110_47# _0444_ 0.01019f
C38488 _0437_ _0434_ 0
C38489 _1000_/a_466_413# _0773_/a_285_297# 0
C38490 _0268_ net165 0
C38491 clknet_1_0__leaf__0462_ _0593_/a_113_47# 0
C38492 _0181_ _0350_ 0.1606f
C38493 net36 _0465_ 0.01663f
C38494 _0227_ net46 0.00982f
C38495 _1009_/a_634_159# _1009_/a_466_413# 0.23992f
C38496 _1009_/a_193_47# _1009_/a_1059_315# 0.03405f
C38497 _1009_/a_27_47# _1009_/a_891_413# 0.03224f
C38498 clknet_1_0__leaf__0460_ hold93/a_285_47# 0.01065f
C38499 VPWR _0518_/a_373_47# 0
C38500 _0243_ net149 0
C38501 hold100/a_285_47# VPWR 0.2783f
C38502 net211 acc0.A\[20\] 0
C38503 _0216_ net247 0
C38504 _1065_/a_634_159# control0.reset 0
C38505 hold5/a_391_47# net198 0
C38506 hold5/a_285_47# net18 0
C38507 pp[0] _0207_ 0
C38508 hold18/a_49_47# _0447_ 0
C38509 _0982_/a_634_159# VPWR 0.1841f
C38510 acc0.A\[2\] net36 0
C38511 _0999_/a_1017_47# net41 0
C38512 _0476_ _1066_/a_193_47# 0.03653f
C38513 _0399_ _0831_/a_35_297# 0.035f
C38514 _0279_ _0303_ 0
C38515 _0446_ _0842_/a_59_75# 0.11029f
C38516 net228 _0185_ 0.0888f
C38517 _0817_/a_81_21# _0089_ 0.08811f
C38518 _1036_/a_1059_315# net121 0.003f
C38519 comp0.B\[4\] _1035_/a_27_47# 0.00376f
C38520 net111 _1025_/a_1059_315# 0
C38521 net7 _0548_/a_512_297# 0
C38522 _0238_ _0249_ 0.26007f
C38523 _0967_/a_403_297# net1 0
C38524 _0819_/a_384_47# _0346_ 0
C38525 _0101_ _0228_ 0.02521f
C38526 _0180_ acc0.A\[15\] 0.6502f
C38527 acc0.A\[27\] _1027_/a_27_47# 0.00122f
C38528 net31 _0138_ 0
C38529 _1032_/a_27_47# net118 0.23034f
C38530 comp0.B\[1\] _0565_/a_240_47# 0.0106f
C38531 hold79/a_285_47# _0168_ 0.0361f
C38532 _0557_/a_51_297# _0211_ 0.15686f
C38533 _1014_/a_891_413# _1014_/a_1017_47# 0.00617f
C38534 _1014_/a_634_159# net100 0
C38535 _0959_/a_217_297# _0955_/a_32_297# 0
C38536 _0329_ _0729_/a_68_297# 0
C38537 _1071_/a_1059_315# _1071_/a_891_413# 0.31086f
C38538 _1071_/a_193_47# _1071_/a_975_413# 0
C38539 _1071_/a_466_413# _1071_/a_381_47# 0.03733f
C38540 acc0.A\[15\] net218 0.09433f
C38541 net48 _0973_/a_109_47# 0
C38542 _0996_/a_27_47# _0410_ 0
C38543 _0996_/a_193_47# net238 0.26883f
C38544 _1015_/a_381_47# _0208_ 0.01293f
C38545 _0130_ net201 0
C38546 _1000_/a_27_47# clkbuf_1_0__f__0461_/a_110_47# 0
C38547 clkbuf_1_1__f__0463_/a_110_47# _0176_ 0.00164f
C38548 _0985_/a_1017_47# _0458_ 0
C38549 _1013_/a_634_159# net42 0
C38550 hold10/a_49_47# hold10/a_285_47# 0.22264f
C38551 net203 _0163_ 0.00213f
C38552 _0179_ _0425_ 0
C38553 _0251_ _0830_/a_510_47# 0
C38554 _0343_ _0792_/a_303_47# 0
C38555 hold53/a_285_47# VPWR 0.33219f
C38556 _1035_/a_466_413# net26 0.00661f
C38557 hold39/a_285_47# hold39/a_391_47# 0.41909f
C38558 net139 A[6] 0
C38559 clknet_1_1__leaf__0461_ net41 0
C38560 _0670_/a_215_47# net6 0
C38561 clknet_1_1__leaf__0465_ net146 0.30533f
C38562 control0.sh _0177_ 0
C38563 _0216_ _1024_/a_193_47# 0.00628f
C38564 acc0.A\[7\] _0437_ 0.09172f
C38565 _0809_/a_299_297# _0345_ 0.01032f
C38566 _0549_/a_68_297# _0549_/a_150_297# 0.00477f
C38567 _0437_ _0989_/a_1059_315# 0
C38568 _0087_ _0989_/a_634_159# 0
C38569 hold65/a_49_47# clknet_0__0465_ 0
C38570 _0305_ _1059_/a_561_413# 0
C38571 acc0.A\[5\] net75 0
C38572 _0089_ _0084_ 0
C38573 hold98/a_391_47# pp[14] 0.00987f
C38574 net86 _0116_ 0
C38575 _1027_/a_27_47# _0364_ 0
C38576 _0343_ _0659_/a_68_297# 0.0041f
C38577 _1015_/a_891_413# net17 0
C38578 _0186_ _0523_/a_299_297# 0.04788f
C38579 VPWR _0206_ 1.27843f
C38580 net36 _1039_/a_381_47# 0.01662f
C38581 _0195_ _1048_/a_891_413# 0.00416f
C38582 net88 _1067_/a_381_47# 0
C38583 _1042_/a_891_413# _0542_/a_51_297# 0
C38584 _1012_/a_891_413# _0352_ 0.02008f
C38585 pp[26] hold9/a_391_47# 0
C38586 _0608_/a_27_47# _0240_ 0.0517f
C38587 _0112_ control0.sh 0
C38588 clknet_1_0__leaf__0458_ _0500_/a_27_47# 0
C38589 _0343_ _1016_/a_561_413# 0
C38590 _1033_/a_634_159# _0215_ 0
C38591 net180 _0472_ 0
C38592 _0172_ _0473_ 0.30748f
C38593 clknet_1_0__leaf__0459_ _1017_/a_634_159# 0
C38594 _0433_ _0271_ 0.0023f
C38595 clknet_1_1__leaf__0459_ _0812_/a_79_21# 0.01138f
C38596 _0253_ acc0.A\[6\] 0.44587f
C38597 net150 _0222_ 0
C38598 hold36/a_49_47# comp0.B\[14\] 0.33204f
C38599 _1069_/a_27_47# _1069_/a_193_47# 0.96995f
C38600 _0369_ _0825_/a_150_297# 0
C38601 input25/a_75_212# control0.sh 0
C38602 hold25/a_391_47# net7 0
C38603 _0579_/a_373_47# clknet_1_0__leaf__0457_ 0
C38604 _0981_/a_373_47# _0170_ 0
C38605 net162 _0341_ 0
C38606 pp[20] pp[23] 0.08753f
C38607 _1052_/a_561_413# _0180_ 0
C38608 hold54/a_391_47# comp0.B\[0\] 0
C38609 _0786_/a_80_21# _0296_ 0
C38610 hold89/a_285_47# _0478_ 0
C38611 _0225_ _0606_/a_109_53# 0
C38612 _0179_ _0180_ 0.72471f
C38613 _1037_/a_27_47# net161 0
C38614 _0135_ _1036_/a_27_47# 0
C38615 hold20/a_285_47# _0483_ 0.00116f
C38616 _0179_ net218 0
C38617 hold42/a_285_47# pp[10] 0
C38618 _0174_ net29 0.05776f
C38619 clkbuf_1_1__f__0464_/a_110_47# _0172_ 0.00366f
C38620 comp0.B\[7\] hold25/a_49_47# 0
C38621 _0512_/a_27_297# acc0.A\[11\] 0.06226f
C38622 net101 net23 0
C38623 _1030_/a_27_47# hold62/a_391_47# 0
C38624 _1030_/a_193_47# hold62/a_285_47# 0
C38625 _1030_/a_634_159# hold62/a_49_47# 0
C38626 _0305_ _0731_/a_299_297# 0
C38627 VPWR _0508_/a_81_21# 0.19916f
C38628 _0399_ _1060_/a_193_47# 0
C38629 _0985_/a_193_47# _0350_ 0
C38630 B[14] net152 0
C38631 _0975_/a_145_75# _0468_ 0
C38632 _0477_ clknet_1_1__leaf_clk 0.72931f
C38633 _0084_ _0986_/a_891_413# 0
C38634 _0550_/a_51_297# comp0.B\[8\] 0
C38635 _0718_/a_47_47# output56/a_27_47# 0.01669f
C38636 _0369_ net229 0
C38637 hold97/a_391_47# acc0.A\[27\] 0.00811f
C38638 hold96/a_391_47# _1024_/a_193_47# 0
C38639 hold96/a_285_47# _1024_/a_634_159# 0
C38640 _1053_/a_466_413# net9 0
C38641 _0399_ _0988_/a_381_47# 0
C38642 net36 net174 0
C38643 clkload1/Y _0257_ 0.02751f
C38644 _0216_ net100 0
C38645 _0130_ comp0.B\[2\] 0
C38646 _0260_ _0846_/a_51_297# 0
C38647 clknet_1_1__leaf__0462_ _1008_/a_466_413# 0.00192f
C38648 _0129_ clknet_1_1__leaf__0462_ 0
C38649 net157 _0177_ 0.02959f
C38650 comp0.B\[6\] _0561_/a_51_297# 0.00528f
C38651 pp[9] _1057_/a_561_413# 0
C38652 _0457_ _0399_ 0
C38653 VPWR _1046_/a_1059_315# 0.38419f
C38654 _0172_ _0186_ 0.02225f
C38655 _0231_ _0325_ 0
C38656 _1022_/a_27_47# _1022_/a_561_413# 0.0027f
C38657 _1022_/a_634_159# _1022_/a_891_413# 0.03684f
C38658 _1022_/a_193_47# _1022_/a_381_47# 0.0982f
C38659 _0645_/a_285_47# _0644_/a_47_47# 0.00217f
C38660 _0164_ _0468_ 0.0123f
C38661 _0686_/a_301_297# _0318_ 0.0018f
C38662 output47/a_27_47# acc0.A\[9\] 0
C38663 hold49/a_49_47# _0172_ 0.03348f
C38664 _0717_/a_209_297# acc0.A\[30\] 0
C38665 _0684_/a_59_75# VPWR 0.23327f
C38666 _1052_/a_634_159# _0525_/a_299_297# 0
C38667 acc0.A\[27\] net96 0
C38668 clkbuf_1_1__f__0460_/a_110_47# _0321_ 0
C38669 input7/a_75_212# net7 0.10851f
C38670 _0416_ _0281_ 0.00144f
C38671 _0275_ _0986_/a_27_47# 0.09052f
C38672 _0274_ _0986_/a_193_47# 0
C38673 _0272_ _0986_/a_634_159# 0
C38674 _0112_ net157 0
C38675 _0957_/a_220_297# _0474_ 0.01077f
C38676 _1018_/a_1017_47# _0116_ 0
C38677 net104 net206 0.35549f
C38678 net211 _1001_/a_193_47# 0.3181f
C38679 net150 net220 0
C38680 _0292_ _0812_/a_79_21# 0.03528f
C38681 clkbuf_0_clk/a_110_47# _0488_ 0
C38682 pp[7] output63/a_27_47# 0.04581f
C38683 clknet_1_1__leaf__0459_ _0347_ 0.02268f
C38684 _1055_/a_634_159# _1055_/a_592_47# 0
C38685 _0313_ _0733_/a_79_199# 0
C38686 _0505_/a_109_297# net6 0.00625f
C38687 hold43/a_49_47# hold43/a_391_47# 0.00188f
C38688 _0280_ VPWR 1.01443f
C38689 _0559_/a_240_47# _0208_ 0.07519f
C38690 _0771_/a_298_297# _0771_/a_382_47# 0
C38691 _0133_ comp0.B\[6\] 0.40116f
C38692 net89 hold12/a_391_47# 0.002f
C38693 _1003_/a_466_413# _1003_/a_381_47# 0.03733f
C38694 _1003_/a_193_47# _1003_/a_975_413# 0
C38695 _1003_/a_1059_315# _1003_/a_891_413# 0.31086f
C38696 hold14/a_391_47# _1036_/a_193_47# 0.00283f
C38697 hold14/a_285_47# _1036_/a_634_159# 0.01163f
C38698 _0466_ _1063_/a_193_47# 0
C38699 hold97/a_391_47# _0364_ 0
C38700 _0954_/a_32_297# _0540_/a_51_297# 0.00321f
C38701 VPWR _0246_ 0.5495f
C38702 VPWR _0687_/a_145_75# 0
C38703 _0248_ _0763_/a_109_47# 0.00149f
C38704 hold64/a_285_47# _0216_ 0.05351f
C38705 net171 _1040_/a_27_47# 0
C38706 _0289_ net228 0.14048f
C38707 _0168_ _0970_/a_285_47# 0
C38708 net247 _1048_/a_466_413# 0
C38709 net185 _0955_/a_304_297# 0.00164f
C38710 _0212_ _0955_/a_220_297# 0
C38711 _0558_/a_150_297# comp0.B\[5\] 0
C38712 hold58/a_49_47# net205 0.00106f
C38713 clkbuf_0__0461_/a_110_47# _0245_ 0.01098f
C38714 _0231_ _0238_ 0
C38715 net22 _1042_/a_634_159# 0
C38716 VPWR _0747_/a_510_47# 0
C38717 _1054_/a_634_159# _0191_ 0
C38718 _0525_/a_81_21# _0194_ 0.17045f
C38719 _0830_/a_297_297# clknet_1_1__leaf__0458_ 0.0014f
C38720 _0525_/a_384_47# net12 0
C38721 net29 _0208_ 0.08985f
C38722 clknet_1_1__leaf__0460_ _0106_ 0
C38723 acc0.A\[27\] _0315_ 0
C38724 net235 _0439_ 0.13594f
C38725 _0086_ _0438_ 0
C38726 _0764_/a_384_47# _0384_ 0
C38727 clkload0/a_27_47# clknet_1_0__leaf_clk 0.22611f
C38728 _0844_/a_79_21# _0844_/a_297_47# 0.03259f
C38729 _1004_/a_891_413# _0347_ 0
C38730 _1004_/a_634_159# _0352_ 0
C38731 _1004_/a_193_47# _0102_ 0.53656f
C38732 hold59/a_285_47# _0459_ 0
C38733 net74 acc0.A\[6\] 0.00295f
C38734 _0151_ net9 0
C38735 net53 _0313_ 0.31005f
C38736 _0199_ clknet_1_1__leaf__0457_ 0.29862f
C38737 VPWR net235 0.15815f
C38738 _0244_ _0181_ 0
C38739 _0502_/a_27_47# clknet_1_0__leaf__0464_ 0.02195f
C38740 _0534_/a_81_21# _0531_/a_109_297# 0
C38741 clknet_0__0458_ _0369_ 0.00364f
C38742 _0442_ acc0.A\[5\] 0.08083f
C38743 net70 _0184_ 0.00241f
C38744 net66 _0187_ 0
C38745 net23 _1065_/a_27_47# 0.02657f
C38746 VPWR _0270_ 0.4389f
C38747 _1054_/a_466_413# _1053_/a_891_413# 0
C38748 _0765_/a_79_21# hold73/a_49_47# 0.00163f
C38749 _1012_/a_193_47# _0350_ 0
C38750 VPWR _0987_/a_466_413# 0.27368f
C38751 _1024_/a_27_47# _1024_/a_634_159# 0.14145f
C38752 _1058_/a_891_413# net189 0.00134f
C38753 _0276_ _0788_/a_150_297# 0
C38754 _0557_/a_245_297# net160 0
C38755 _0858_/a_27_47# VPWR 0.29884f
C38756 hold64/a_391_47# clknet_0__0457_ 0.00268f
C38757 input32/a_75_212# _1042_/a_27_47# 0
C38758 _0292_ _0347_ 0
C38759 clknet_1_0__leaf__0458_ _0275_ 0
C38760 output61/a_27_47# acc0.A\[6\] 0
C38761 _0664_/a_297_47# _0296_ 0.00964f
C38762 _1059_/a_561_413# _0181_ 0
C38763 _1000_/a_466_413# _0244_ 0
C38764 _1000_/a_193_47# _0388_ 0
C38765 _1000_/a_634_159# _0386_ 0
C38766 VPWR _1029_/a_466_413# 0.2739f
C38767 _0462_ _0218_ 0
C38768 _0315_ _0364_ 0
C38769 hold59/a_391_47# clknet_1_0__leaf__0461_ 0.00305f
C38770 _1055_/a_1059_315# net142 0
C38771 _0540_/a_51_297# _0540_/a_245_297# 0.01218f
C38772 _0982_/a_634_159# _0453_ 0
C38773 _0982_/a_891_413# _0452_ 0
C38774 hold61/a_285_47# hold61/a_391_47# 0.41909f
C38775 _1048_/a_634_159# _1048_/a_1059_315# 0
C38776 _1048_/a_27_47# _1048_/a_381_47# 0.06222f
C38777 _1048_/a_193_47# _1048_/a_891_413# 0.19489f
C38778 _0786_/a_80_21# _0811_/a_81_21# 0.01709f
C38779 _1034_/a_27_47# clknet_1_1__leaf__0463_ 0.06548f
C38780 _0195_ _0790_/a_35_297# 0
C38781 VPWR net103 1.01518f
C38782 _0399_ _0796_/a_79_21# 0.13746f
C38783 net235 output62/a_27_47# 0
C38784 _0833_/a_215_47# pp[4] 0
C38785 clkbuf_1_0__f__0461_/a_110_47# acc0.A\[19\] 0.01503f
C38786 _0607_/a_109_297# _0780_/a_35_297# 0
C38787 _0232_ _0742_/a_384_47# 0
C38788 net116 _0219_ 0.04208f
C38789 net220 control0.add 0
C38790 _0555_/a_240_47# VPWR 0.01074f
C38791 _0312_ _1007_/a_466_413# 0
C38792 _0981_/a_27_297# clknet_1_0__leaf_clk 0.02779f
C38793 net120 _0562_/a_68_297# 0
C38794 clknet_1_0__leaf__0457_ _0345_ 0.16186f
C38795 hold11/a_285_47# hold11/a_391_47# 0.41909f
C38796 _0179_ hold70/a_285_47# 0
C38797 _0680_/a_217_297# clkbuf_0__0460_/a_110_47# 0
C38798 VPWR _1033_/a_1017_47# 0
C38799 _0387_ _0677_/a_285_47# 0
C38800 clknet_0_clk _0161_ 0.65151f
C38801 net1 _0721_/a_27_47# 0.0168f
C38802 _0343_ net209 0
C38803 hold59/a_285_47# _0265_ 0
C38804 _0402_ _0399_ 0
C38805 _0390_ _0246_ 0
C38806 clknet_0__0459_ net228 0.01493f
C38807 _0252_ _0434_ 0.03161f
C38808 _0518_/a_109_297# acc0.A\[6\] 0.05658f
C38809 net187 hold73/a_285_47# 0.00161f
C38810 net45 _0774_/a_68_297# 0.10943f
C38811 net233 VPWR 0.19258f
C38812 _0172_ _0497_/a_68_297# 0.03122f
C38813 net152 _0544_/a_51_297# 0.05982f
C38814 _0151_ _1054_/a_891_413# 0
C38815 hold76/a_285_47# hold76/a_391_47# 0.41909f
C38816 clknet_0__0463_ _0560_/a_68_297# 0.00134f
C38817 _1010_/a_193_47# net96 0.00549f
C38818 _1010_/a_1059_315# _1010_/a_1017_47# 0
C38819 _0348_ net57 0.03012f
C38820 _0153_ acc0.A\[8\] 0
C38821 hold6/a_49_47# _0546_/a_240_47# 0
C38822 _0130_ _1015_/a_193_47# 0
C38823 hold55/a_391_47# _1015_/a_1059_315# 0.00124f
C38824 hold55/a_285_47# _1015_/a_891_413# 0.00163f
C38825 hold92/a_285_47# _0219_ 0
C38826 net165 net222 0
C38827 clknet_1_1__leaf__0461_ _0350_ 0
C38828 _1040_/a_634_159# _1040_/a_592_47# 0
C38829 hold74/a_49_47# acc0.A\[16\] 0.34605f
C38830 _0768_/a_109_297# _0310_ 0.01151f
C38831 _0410_ _0794_/a_27_47# 0
C38832 _0266_ _0451_ 0
C38833 _0111_ clknet_1_1__leaf__0461_ 0.00378f
C38834 _0432_ _0441_ 0.00644f
C38835 _1072_/a_27_47# _1072_/a_634_159# 0.13601f
C38836 hold88/a_285_47# clknet_1_1__leaf__0465_ 0
C38837 _0527_/a_27_297# net154 0.06634f
C38838 _0216_ _1027_/a_891_413# 0.05528f
C38839 _0853_/a_150_297# _0346_ 0.00144f
C38840 comp0.B\[1\] _0171_ 0
C38841 net88 net150 0
C38842 _1002_/a_1017_47# _0183_ 0
C38843 _0328_ _0323_ 0.0481f
C38844 _0273_ _0829_/a_27_47# 0
C38845 VPWR _1019_/a_1059_315# 0.39924f
C38846 control0.state\[1\] _0469_ 0.00101f
C38847 _0765_/a_79_21# _0181_ 0
C38848 _0749_/a_299_297# net92 0
C38849 input19/a_75_212# net10 0.00381f
C38850 net1 _0760_/a_285_47# 0
C38851 _0743_/a_240_47# hold90/a_285_47# 0
C38852 _0635_/a_27_47# _0345_ 0.01089f
C38853 acc0.A\[14\] _0996_/a_381_47# 0
C38854 _0218_ _0297_ 0.05769f
C38855 _0343_ hold72/a_49_47# 0
C38856 comp0.B\[5\] input27/a_75_212# 0
C38857 _1067_/a_634_159# _1067_/a_592_47# 0
C38858 _0174_ _0137_ 0.07096f
C38859 net34 _0468_ 0.05093f
C38860 hold1/a_391_47# net154 0
C38861 clknet_1_0__leaf__0465_ _0433_ 0.039f
C38862 _0244_ _1018_/a_27_47# 0.00102f
C38863 _0458_ net9 0
C38864 _0251_ _0989_/a_193_47# 0.03166f
C38865 _0800_/a_240_47# _0410_ 0
C38866 hold31/a_49_47# hold31/a_285_47# 0.22264f
C38867 net178 _0369_ 0.00526f
C38868 clknet_1_1__leaf__0460_ _1011_/a_27_47# 0.01039f
C38869 hold35/a_285_47# A[10] 0.00865f
C38870 hold12/a_285_47# net35 0.08238f
C38871 _1071_/a_634_159# _0169_ 0.00101f
C38872 net199 _0102_ 0
C38873 control0.count\[3\] net49 0
C38874 hold90/a_391_47# _0345_ 0.0282f
C38875 _1004_/a_1059_315# _0757_/a_68_297# 0.00151f
C38876 acc0.A\[7\] _0252_ 0.79653f
C38877 _0086_ clknet_1_1__leaf__0465_ 0
C38878 net57 _0332_ 0
C38879 control0.state\[1\] _1002_/a_634_159# 0
C38880 _0717_/a_80_21# _0717_/a_303_47# 0.01146f
C38881 _0717_/a_209_297# _0717_/a_209_47# 0
C38882 _0252_ _0989_/a_1059_315# 0.05378f
C38883 net65 _0989_/a_561_413# 0
C38884 _0343_ hold87/a_49_47# 0
C38885 _0989_/a_466_413# _0989_/a_561_413# 0.00772f
C38886 _0989_/a_634_159# _0989_/a_975_413# 0
C38887 _0997_/a_27_47# _0997_/a_634_159# 0.13601f
C38888 _1020_/a_193_47# clknet_1_0__leaf__0461_ 0
C38889 net228 _0418_ 0
C38890 _0129_ hold92/a_49_47# 0
C38891 _0412_ _0218_ 0
C38892 _0181_ _0986_/a_634_159# 0.00119f
C38893 _0544_/a_149_47# _1042_/a_27_47# 0
C38894 _0544_/a_51_297# _1042_/a_466_413# 0.00193f
C38895 _0248_ _0616_/a_215_47# 0.00446f
C38896 net68 VPWR 0.3817f
C38897 _0292_ clkbuf_0__0465_/a_110_47# 0
C38898 hold30/a_49_47# net46 0.02196f
C38899 acc0.A\[16\] _0583_/a_27_297# 0.1318f
C38900 _0992_/a_193_47# _0992_/a_592_47# 0.00135f
C38901 _0992_/a_466_413# _0992_/a_561_413# 0.00772f
C38902 _0992_/a_634_159# _0992_/a_975_413# 0
C38903 VPWR _1051_/a_27_47# 0.69912f
C38904 _0749_/a_81_21# _0369_ 0
C38905 clkbuf_1_1__f__0459_/a_110_47# net41 0
C38906 _0498_/a_51_297# acc0.A\[15\] 0
C38907 net26 _0561_/a_51_297# 0
C38908 net7 _0138_ 0.25977f
C38909 _0678_/a_68_297# _0240_ 0
C38910 _1002_/a_1059_315# _0603_/a_68_297# 0
C38911 VPWR _1045_/a_634_159# 0.18102f
C38912 _0402_ _0808_/a_266_297# 0.00253f
C38913 net158 net247 0
C38914 _0125_ _1027_/a_975_413# 0.00111f
C38915 _0766_/a_109_297# _0240_ 0
C38916 _0337_ pp[27] 0.03678f
C38917 _0280_ _0283_ 0.14285f
C38918 clkbuf_1_0__f__0458_/a_110_47# _0841_/a_215_47# 0
C38919 _0355_ _1029_/a_891_413# 0
C38920 _0109_ _1029_/a_193_47# 0
C38921 hold13/a_49_47# comp0.B\[5\] 0.3337f
C38922 clkbuf_0__0463_/a_110_47# _0493_/a_27_47# 0
C38923 clknet_1_1__leaf__0464_ net148 0
C38924 _0793_/a_149_47# _0792_/a_80_21# 0
C38925 clknet_0__0458_ _0846_/a_240_47# 0
C38926 _0963_/a_117_297# _0466_ 0
C38927 hold1/a_285_47# hold7/a_49_47# 0
C38928 _0465_ _1061_/a_27_47# 0.00204f
C38929 _0935_/a_27_47# _1061_/a_891_413# 0
C38930 _0983_/a_634_159# _0116_ 0
C38931 _1061_/a_27_47# _1061_/a_381_47# 0.06222f
C38932 _1061_/a_193_47# _1061_/a_891_413# 0.19685f
C38933 _1061_/a_634_159# _1061_/a_1059_315# 0
C38934 _0680_/a_217_297# _1009_/a_27_47# 0
C38935 net51 _0754_/a_51_297# 0.00604f
C38936 net46 _0352_ 0.07341f
C38937 net69 acc0.A\[14\] 0
C38938 net66 _0990_/a_193_47# 0.03042f
C38939 acc0.A\[8\] _0990_/a_27_47# 0.02599f
C38940 _0133_ net26 0.0312f
C38941 _0554_/a_150_297# net28 0
C38942 _0314_ clknet_1_1__leaf__0460_ 0
C38943 net64 _0153_ 0
C38944 _0216_ _1026_/a_975_413# 0.00121f
C38945 _0195_ _1026_/a_1017_47# 0
C38946 _0124_ _1026_/a_381_47# 0.11825f
C38947 _1007_/a_1059_315# _0219_ 0
C38948 _0174_ comp0.B\[6\] 0.06003f
C38949 _0428_ _0465_ 0
C38950 _0689_/a_150_297# _0364_ 0
C38951 VPWR net143 0.69303f
C38952 _1065_/a_466_413# _1063_/a_27_47# 0
C38953 _0180_ hold83/a_49_47# 0.03225f
C38954 _1035_/a_27_47# _1035_/a_193_47# 0.96668f
C38955 pp[18] _0714_/a_51_297# 0
C38956 _0483_ _0964_/a_109_297# 0
C38957 VPWR output41/a_27_47# 0.29681f
C38958 _0850_/a_68_297# _0345_ 0.05124f
C38959 _0648_/a_277_297# _0277_ 0.00104f
C38960 _0558_/a_68_297# net26 0.01224f
C38961 _0137_ _0208_ 0.00551f
C38962 clkload1/Y clknet_1_1__leaf__0458_ 0.00239f
C38963 net199 _0574_/a_109_47# 0
C38964 _0092_ _0801_/a_113_47# 0
C38965 hold2/a_285_47# _1047_/a_1059_315# 0.00229f
C38966 clkbuf_1_1__f__0462_/a_110_47# _1011_/a_193_47# 0
C38967 _0217_ _1014_/a_381_47# 0.01457f
C38968 _0183_ _1014_/a_1059_315# 0.00259f
C38969 _0787_/a_80_21# _0091_ 0.12356f
C38970 _0787_/a_209_47# _0419_ 0.00297f
C38971 net88 control0.add 0.08502f
C38972 _0489_ _1069_/a_193_47# 0.03652f
C38973 _1065_/a_1059_315# clknet_1_0__leaf__0457_ 0.0026f
C38974 _0372_ clkbuf_0__0460_/a_110_47# 0
C38975 net204 _0175_ 0.00159f
C38976 _0661_/a_27_297# _0423_ 0.01134f
C38977 _0459_ _0219_ 0.03117f
C38978 _0768_/a_109_297# _0768_/a_27_47# 0
C38979 _0328_ net237 0
C38980 VPWR _0637_/a_311_297# 0.00348f
C38981 hold58/a_49_47# net160 0
C38982 net119 _0215_ 0.20416f
C38983 _0984_/a_1017_47# acc0.A\[15\] 0
C38984 clknet_1_0__leaf__0459_ net103 0.23366f
C38985 net76 _0990_/a_634_159# 0
C38986 _0956_/a_32_297# control0.sh 0
C38987 _0343_ _0991_/a_381_47# 0.00987f
C38988 net24 net171 0
C38989 VPWR _1028_/a_975_413# 0.00473f
C38990 _1069_/a_466_413# _1069_/a_592_47# 0.00553f
C38991 _1069_/a_634_159# _1069_/a_1017_47# 0
C38992 _1056_/a_193_47# net66 0
C38993 VPWR _0723_/a_207_413# 0.15716f
C38994 _0402_ _0295_ 0
C38995 net102 _0158_ 0
C38996 _0718_/a_285_47# pp[30] 0
C38997 _0243_ net206 0
C38998 hold69/a_391_47# _0324_ 0
C38999 _1059_/a_1059_315# acc0.A\[13\] 0.14049f
C39000 _1059_/a_193_47# net5 0
C39001 _0954_/a_304_297# comp0.B\[12\] 0
C39002 pp[16] hold78/a_391_47# 0
C39003 _0753_/a_79_21# _0223_ 0
C39004 _0343_ _0600_/a_103_199# 0.01037f
C39005 _1062_/a_27_47# hold84/a_285_47# 0
C39006 VPWR input3/a_75_212# 0.24854f
C39007 _0225_ _0238_ 0.00875f
C39008 _1041_/a_1059_315# _1040_/a_634_159# 0
C39009 _1041_/a_891_413# _1040_/a_193_47# 0
C39010 _1031_/a_381_47# _0220_ 0.02068f
C39011 comp0.B\[3\] _0160_ 0
C39012 _0200_ _0172_ 0.00227f
C39013 net31 net22 0.04412f
C39014 _0997_/a_193_47# _0411_ 0
C39015 _0399_ _1017_/a_1059_315# 0
C39016 hold66/a_391_47# _0383_ 0
C39017 net213 _0762_/a_510_47# 0
C39018 hold55/a_285_47# net87 0
C39019 hold64/a_49_47# hold64/a_391_47# 0.00188f
C39020 _0482_ VPWR 0.34741f
C39021 _0990_/a_193_47# _0350_ 0
C39022 hold23/a_49_47# VPWR 0.32549f
C39023 clknet_1_0__leaf__0460_ _1063_/a_27_47# 0
C39024 _1030_/a_381_47# net209 0.12224f
C39025 B[12] hold51/a_285_47# 0.00238f
C39026 _0386_ _0242_ 0
C39027 _1018_/a_891_413# clknet_0__0461_ 0
C39028 _0397_ clknet_0__0461_ 0
C39029 _1051_/a_891_413# net9 0.00466f
C39030 hold22/a_49_47# net63 0
C39031 _0172_ comp0.B\[8\] 0.03553f
C39032 _1002_/a_381_47# _0181_ 0.00308f
C39033 hold89/a_49_47# _0479_ 0
C39034 hold96/a_285_47# net110 0.00192f
C39035 hold12/a_391_47# clkbuf_0_clk/a_110_47# 0.01439f
C39036 _0217_ _1022_/a_634_159# 0
C39037 _0183_ _1022_/a_27_47# 0.0097f
C39038 acc0.A\[22\] _1022_/a_193_47# 0.00604f
C39039 _0343_ clknet_0__0461_ 0.02157f
C39040 _0561_/a_51_297# hold84/a_285_47# 0
C39041 clknet_0__0457_ clkbuf_1_1__f__0457_/a_110_47# 0.32353f
C39042 _0538_/a_245_297# net183 0
C39043 _0538_/a_149_47# _0201_ 0.00154f
C39044 _0538_/a_51_297# net21 0.09158f
C39045 hold6/a_285_47# _0176_ 0
C39046 _0462_ _0099_ 0
C39047 hold30/a_285_47# VPWR 0.28219f
C39048 comp0.B\[6\] _0208_ 0.16324f
C39049 _0524_/a_27_297# _0524_/a_109_297# 0.17136f
C39050 hold67/a_285_47# acc0.A\[9\] 0.00546f
C39051 clknet_1_0__leaf__0463_ net31 0.02755f
C39052 _1022_/a_1059_315# net151 0
C39053 net53 _0572_/a_109_297# 0
C39054 _1065_/a_466_413# _1062_/a_1059_315# 0
C39055 _1065_/a_381_47# _1062_/a_193_47# 0
C39056 hold22/a_285_47# net15 0.00631f
C39057 _0357_ _0329_ 0.0725f
C39058 net64 _0990_/a_27_47# 0
C39059 clknet_1_0__leaf__0459_ _1019_/a_1059_315# 0.01352f
C39060 clkbuf_1_0__f__0462_/a_110_47# _0219_ 0.01645f
C39061 hold12/a_49_47# net159 0
C39062 _1003_/a_193_47# _0974_/a_79_199# 0
C39063 _0987_/a_193_47# acc0.A\[6\] 0
C39064 net199 _1025_/a_1059_315# 0
C39065 _0328_ _0686_/a_27_53# 0.0016f
C39066 _0994_/a_634_159# _0994_/a_592_47# 0
C39067 acc0.A\[26\] _0360_ 0
C39068 _0259_ _0819_/a_384_47# 0
C39069 _1020_/a_561_413# clknet_1_0__leaf__0457_ 0
C39070 _0358_ _0327_ 0
C39071 _0285_ _0417_ 0.22815f
C39072 _0579_/a_27_297# net223 0
C39073 _0779_/a_215_47# _0396_ 0.00549f
C39074 _0779_/a_79_21# _0097_ 0.05919f
C39075 _0289_ _0090_ 0
C39076 _0462_ _0359_ 0.74164f
C39077 _0305_ _0195_ 0.03505f
C39078 _0260_ _0643_/a_253_297# 0
C39079 VPWR _0739_/a_510_47# 0.00109f
C39080 _0803_/a_68_297# _0279_ 0
C39081 _1023_/a_1059_315# net51 0.00114f
C39082 _0337_ _0216_ 0
C39083 _0349_ _0195_ 0.0242f
C39084 _0835_/a_292_297# _0256_ 0.00443f
C39085 _0835_/a_78_199# _0271_ 0
C39086 _0464_ _1046_/a_27_47# 0.0016f
C39087 comp0.B\[15\] _0584_/a_27_297# 0
C39088 hold22/a_285_47# _1053_/a_1059_315# 0.0054f
C39089 _0855_/a_299_297# _0350_ 0.05906f
C39090 VPWR _0102_ 0.46882f
C39091 net169 net63 0
C39092 hold14/a_49_47# net161 0
C39093 _1003_/a_381_47# _0101_ 0.1311f
C39094 net36 _1047_/a_975_413# 0
C39095 _0993_/a_27_47# _0993_/a_634_159# 0.14145f
C39096 input3/a_75_212# input4/a_75_212# 0
C39097 _1058_/a_193_47# net192 0
C39098 _1065_/a_27_47# _0213_ 0
C39099 _1039_/a_634_159# _1039_/a_1059_315# 0
C39100 _1039_/a_27_47# _1039_/a_381_47# 0.05761f
C39101 _1039_/a_193_47# _1039_/a_891_413# 0.19226f
C39102 _0476_ VPWR 1.63107f
C39103 _0357_ _0221_ 0.06108f
C39104 hold33/a_391_47# net173 0
C39105 _0258_ _0640_/a_215_297# 0
C39106 net7 net134 0
C39107 _1020_/a_891_413# _0457_ 0
C39108 _0279_ _0672_/a_215_47# 0
C39109 net193 _0172_ 0.00871f
C39110 net22 net128 0
C39111 net140 _0191_ 0
C39112 _0985_/a_1059_315# net170 0
C39113 _1056_/a_27_47# net64 0
C39114 _0372_ _1009_/a_27_47# 0
C39115 A[12] _0512_/a_27_297# 0.07631f
C39116 hold27/a_285_47# net157 0.01449f
C39117 _0172_ _1046_/a_466_413# 0.01794f
C39118 _1010_/a_1059_315# _0332_ 0
C39119 _0257_ _0989_/a_1017_47# 0
C39120 _0447_ _0448_ 0.04068f
C39121 hold14/a_49_47# net26 0.00287f
C39122 input26/a_75_212# B[4] 0.00567f
C39123 _1026_/a_634_159# _1026_/a_466_413# 0.23992f
C39124 _1026_/a_193_47# _1026_/a_1059_315# 0.03405f
C39125 _1026_/a_27_47# _1026_/a_891_413# 0.03224f
C39126 net33 _1062_/a_381_47# 0
C39127 VPWR A[4] 0.19433f
C39128 _0733_/a_79_199# _0321_ 0.00759f
C39129 _0733_/a_222_93# _0360_ 0.09853f
C39130 _0343_ _0082_ 0.02731f
C39131 _0985_/a_466_413# clknet_1_0__leaf__0458_ 0.00188f
C39132 hold10/a_49_47# _1047_/a_27_47# 0.02457f
C39133 _0750_/a_27_47# _0228_ 0
C39134 _1021_/a_634_159# clknet_1_0__leaf__0460_ 0.00959f
C39135 net162 acc0.A\[30\] 0.00266f
C39136 VPWR _0774_/a_68_297# 0.14832f
C39137 net61 acc0.A\[6\] 0.02434f
C39138 hold59/a_391_47# _0218_ 0.01854f
C39139 net169 _1053_/a_891_413# 0.00171f
C39140 net140 _1053_/a_381_47# 0
C39141 _0982_/a_1059_315# _0399_ 0
C39142 _0258_ _0465_ 0.01302f
C39143 _0715_/a_27_47# _0662_/a_81_21# 0
C39144 _1032_/a_891_413# clknet_1_1__leaf_clk 0
C39145 VPWR A[1] 0.24657f
C39146 comp0.B\[4\] _0959_/a_80_21# 0.00759f
C39147 VPWR _0085_ 0.39259f
C39148 _0217_ _1067_/a_1059_315# 0
C39149 _1024_/a_891_413# _1024_/a_975_413# 0.00851f
C39150 _1024_/a_27_47# net110 0.23044f
C39151 _1024_/a_381_47# _1024_/a_561_413# 0.00123f
C39152 net45 hold72/a_391_47# 0.01474f
C39153 net227 _0723_/a_297_47# 0
C39154 acc0.A\[20\] _0461_ 0.00277f
C39155 _0995_/a_891_413# A[13] 0
C39156 _0718_/a_285_47# _0339_ 0.00953f
C39157 _1014_/a_27_47# _0181_ 0.00207f
C39158 _1021_/a_891_413# _1020_/a_466_413# 0
C39159 _0121_ hold29/a_49_47# 0.00236f
C39160 clknet_1_1__leaf__0464_ _0542_/a_240_47# 0
C39161 _0220_ _0219_ 0.04015f
C39162 _0438_ net66 0
C39163 net244 _0321_ 0
C39164 net246 _0281_ 0.00571f
C39165 hold97/a_285_47# hold97/a_391_47# 0.41909f
C39166 net217 clknet_1_1__leaf__0465_ 0
C39167 _0098_ _0244_ 0.00165f
C39168 VPWR net191 0.45691f
C39169 _0574_/a_109_47# VPWR 0
C39170 hold89/a_285_47# VPWR 0.2765f
C39171 _0151_ hold22/a_391_47# 0
C39172 _0180_ _1049_/a_891_413# 0.00815f
C39173 _0786_/a_80_21# _0992_/a_634_159# 0
C39174 _0786_/a_217_297# _0992_/a_193_47# 0
C39175 A[11] clknet_1_1__leaf__0465_ 0.03578f
C39176 _0731_/a_81_21# clknet_0__0460_ 0
C39177 _0540_/a_512_297# net20 0
C39178 clk _1064_/a_975_413# 0
C39179 _0268_ acc0.A\[3\] 0.00136f
C39180 control0.add _0771_/a_298_297# 0
C39181 net53 _0321_ 0.00997f
C39182 _0402_ _0811_/a_299_297# 0.06342f
C39183 pp[6] VPWR 0.58888f
C39184 acc0.A\[14\] _0300_ 0
C39185 B[13] _1043_/a_193_47# 0
C39186 hold11/a_49_47# _0142_ 0
C39187 _0464_ _0178_ 0
C39188 _1068_/a_466_413# _0468_ 0.02224f
C39189 _1041_/a_27_47# _1041_/a_193_47# 0.9657f
C39190 _0343_ _1013_/a_466_413# 0
C39191 net1 _0182_ 0
C39192 _0234_ _0751_/a_111_297# 0
C39193 _0223_ clkbuf_1_0__f__0460_/a_110_47# 0.00977f
C39194 _0312_ _0105_ 0.00381f
C39195 _0170_ clknet_1_0__leaf_clk 0.0365f
C39196 _0416_ _0803_/a_68_297# 0.10709f
C39197 _0415_ _0803_/a_150_297# 0
C39198 _0399_ _0451_ 0.24503f
C39199 _0787_/a_80_21# _0346_ 0
C39200 _0748_/a_299_297# net52 0
C39201 _0340_ _0708_/a_150_297# 0.00134f
C39202 _1015_/a_634_159# comp0.B\[15\] 0
C39203 _0744_/a_27_47# clknet_1_1__leaf__0465_ 0
C39204 _0248_ _0771_/a_215_297# 0
C39205 _0223_ _0250_ 0
C39206 _1057_/a_27_47# _0514_/a_27_297# 0
C39207 hold76/a_49_47# _1001_/a_27_47# 0
C39208 clkbuf_1_0__f__0457_/a_110_47# _0603_/a_68_297# 0
C39209 clkbuf_1_0__f__0457_/a_110_47# hold73/a_391_47# 0
C39210 net185 net33 0
C39211 _0139_ _0204_ 0
C39212 net32 net18 0.1939f
C39213 net167 _0974_/a_222_93# 0
C39214 _0607_/a_109_47# acc0.A\[17\] 0
C39215 clknet_0__0464_ _1061_/a_27_47# 0
C39216 _0118_ net23 0
C39217 clknet_0__0460_ _1006_/a_193_47# 0
C39218 _0616_/a_78_199# acc0.A\[19\] 0
C39219 hold69/a_391_47# _0104_ 0
C39220 _1056_/a_381_47# _0189_ 0
C39221 hold6/a_391_47# _0139_ 0.05234f
C39222 _1040_/a_975_413# net174 0
C39223 _0607_/a_27_297# clkbuf_1_1__f__0461_/a_110_47# 0
C39224 _1053_/a_561_413# acc0.A\[6\] 0
C39225 _1057_/a_193_47# _0512_/a_27_297# 0
C39226 hold44/a_49_47# _1029_/a_27_47# 0.01435f
C39227 output64/a_27_47# pp[4] 0.04597f
C39228 _0438_ _0350_ 0.06772f
C39229 _0249_ _1006_/a_891_413# 0
C39230 _0250_ _1006_/a_1059_315# 0
C39231 _1072_/a_891_413# _1072_/a_975_413# 0.00851f
C39232 _1072_/a_381_47# _1072_/a_561_413# 0.00123f
C39233 _0437_ _0186_ 0.0504f
C39234 _0343_ _0984_/a_193_47# 0.02689f
C39235 _0124_ net156 0
C39236 _0841_/a_510_47# _0445_ 0.00404f
C39237 _0369_ _0675_/a_68_297# 0
C39238 _0137_ comp0.B\[9\] 0
C39239 hold39/a_49_47# clknet_0__0463_ 0
C39240 net65 _0831_/a_35_297# 0.01354f
C39241 hold38/a_391_47# hold39/a_49_47# 0.0012f
C39242 hold38/a_285_47# hold39/a_285_47# 0.01958f
C39243 hold38/a_49_47# hold39/a_391_47# 0.0012f
C39244 output57/a_27_47# _0333_ 0
C39245 _0267_ _0219_ 0.02218f
C39246 _1013_/a_634_159# net60 0
C39247 hold68/a_285_47# _0347_ 0
C39248 _0471_ _1062_/a_193_47# 0
C39249 hold36/a_285_47# clknet_1_0__leaf__0465_ 0.00808f
C39250 VPWR _1025_/a_1059_315# 0.4575f
C39251 _0537_/a_68_297# net184 0
C39252 _1067_/a_891_413# control0.add 0.00293f
C39253 acc0.A\[27\] _0691_/a_150_297# 0
C39254 net61 _0624_/a_59_75# 0
C39255 comp0.B\[4\] _0173_ 0.00283f
C39256 net161 _0208_ 0
C39257 VPWR clkbuf_0__0463_/a_110_47# 1.31379f
C39258 _1041_/a_891_413# _0207_ 0
C39259 _0239_ _0097_ 0
C39260 _1012_/a_634_159# _0722_/a_215_47# 0
C39261 net136 _0172_ 0
C39262 _0195_ _0181_ 0.37221f
C39263 _0476_ _0559_/a_245_297# 0
C39264 _0891_/a_27_47# _0457_ 0.01068f
C39265 _0217_ _1024_/a_891_413# 0
C39266 _1004_/a_975_413# _0380_ 0
C39267 control0.state\[1\] net88 0
C39268 hold75/a_285_47# net233 0
C39269 _0997_/a_891_413# _0997_/a_975_413# 0.00851f
C39270 _0997_/a_381_47# _0997_/a_561_413# 0.00123f
C39271 _0805_/a_27_47# acc0.A\[10\] 0
C39272 _1053_/a_193_47# _0150_ 0
C39273 _1037_/a_466_413# net24 0
C39274 _0810_/a_113_47# _0420_ 0
C39275 _0664_/a_382_297# _0346_ 0
C39276 clknet_1_0__leaf__0457_ hold93/a_49_47# 0.00213f
C39277 _0140_ _1042_/a_193_47# 0.39029f
C39278 net198 _1042_/a_891_413# 0.00238f
C39279 net18 _1042_/a_1059_315# 0
C39280 net46 _0237_ 0
C39281 VPWR _1044_/a_193_47# 0.29969f
C39282 acc0.A\[16\] _0114_ 0.0428f
C39283 acc0.A\[14\] _0404_ 0.00689f
C39284 hold100/a_285_47# _0345_ 0.00323f
C39285 VPWR _0815_/a_113_297# 0.18988f
C39286 _0349_ _1010_/a_891_413# 0.03842f
C39287 net26 _0208_ 0.28473f
C39288 VPWR net131 0.49952f
C39289 _0402_ _0091_ 0.04155f
C39290 hold88/a_49_47# _0399_ 0
C39291 _0783_/a_297_297# _0352_ 0.00581f
C39292 output65/a_27_47# _0828_/a_113_297# 0
C39293 _0254_ _0428_ 0
C39294 clknet_0__0458_ _0084_ 0.00479f
C39295 _0218_ _0417_ 0
C39296 _0243_ _0773_/a_35_297# 0.00628f
C39297 _0756_/a_47_47# _0756_/a_129_47# 0.00369f
C39298 _1000_/a_193_47# _0216_ 0
C39299 _0343_ net145 0
C39300 _0407_ _0405_ 0.09867f
C39301 _0793_/a_240_47# _0408_ 0.04114f
C39302 _1001_/a_193_47# _0461_ 0.00964f
C39303 clkbuf_1_1__f__0465_/a_110_47# _0812_/a_79_21# 0.00183f
C39304 _1027_/a_466_413# _1027_/a_561_413# 0.00772f
C39305 _1027_/a_634_159# _1027_/a_975_413# 0
C39306 _0643_/a_103_199# _0643_/a_253_297# 0.01483f
C39307 _0366_ _0315_ 0.29696f
C39308 hold87/a_285_47# net234 0.0097f
C39309 _0257_ _0261_ 0
C39310 clknet_1_0__leaf__0463_ _0548_/a_240_47# 0
C39311 _0384_ _0374_ 0
C39312 VPWR _0849_/a_297_297# 0.00964f
C39313 net66 clknet_1_1__leaf__0465_ 0.05526f
C39314 net10 net18 0.13032f
C39315 VPWR _1032_/a_381_47# 0.07714f
C39316 net69 _0116_ 0
C39317 _0362_ _0776_/a_27_47# 0
C39318 _0217_ _1072_/a_891_413# 0
C39319 _1061_/a_1059_315# net147 0
C39320 clknet_1_0__leaf__0465_ _0522_/a_109_47# 0
C39321 _0305_ _1009_/a_381_47# 0
C39322 comp0.B\[5\] B[2] 0.00138f
C39323 net51 _0219_ 0.0635f
C39324 _0798_/a_113_297# _0277_ 0
C39325 _0555_/a_512_297# comp0.B\[5\] 0.0022f
C39326 clknet_1_0__leaf__0459_ _0774_/a_68_297# 0
C39327 _0143_ net154 0
C39328 net125 _0214_ 0
C39329 hold21/a_285_47# VPWR 0.2798f
C39330 hold10/a_49_47# net133 0.00194f
C39331 _0346_ _0460_ 0.05913f
C39332 _1065_/a_27_47# _0161_ 0
C39333 _0991_/a_27_47# clknet_1_1__leaf__0465_ 0
C39334 _1035_/a_466_413# _1035_/a_592_47# 0.00553f
C39335 _1035_/a_634_159# _1035_/a_1017_47# 0
C39336 _0668_/a_79_21# _0668_/a_382_297# 0.00145f
C39337 pp[18] net225 0
C39338 _0362_ _0219_ 0.34387f
C39339 clknet_1_0__leaf__0465_ _0835_/a_78_199# 0.00114f
C39340 _1035_/a_466_413# B[15] 0
C39341 output37/a_27_47# _0156_ 0
C39342 _1053_/a_466_413# A[7] 0
C39343 _1053_/a_381_47# input14/a_75_212# 0
C39344 hold76/a_285_47# clknet_1_0__leaf__0461_ 0.00256f
C39345 clknet_1_0__leaf__0462_ net215 0.01689f
C39346 net17 _1064_/a_891_413# 0
C39347 _0946_/a_30_53# _1064_/a_27_47# 0
C39348 _0399_ _0271_ 0
C39349 _1000_/a_891_413# _0247_ 0.05149f
C39350 _0217_ acc0.A\[0\] 0.12321f
C39351 hold7/a_285_47# hold7/a_391_47# 0.41909f
C39352 _0809_/a_81_21# _0809_/a_384_47# 0.00138f
C39353 _0172_ _1045_/a_193_47# 0.03223f
C39354 hold69/a_49_47# _0326_ 0
C39355 VPWR _0533_/a_109_297# 0.19652f
C39356 _0289_ _0401_ 0.56188f
C39357 _0293_ _0423_ 0.26007f
C39358 _0287_ _0290_ 0.08081f
C39359 _0292_ _0425_ 0
C39360 _0983_/a_27_47# net222 0
C39361 VPWR hold71/a_49_47# 0.30223f
C39362 _1048_/a_891_413# acc0.A\[15\] 0
C39363 _1030_/a_27_47# _0334_ 0
C39364 clknet_1_1__leaf__0459_ _1013_/a_193_47# 0
C39365 _1010_/a_891_413# _0701_/a_209_297# 0
C39366 _0460_ hold94/a_49_47# 0
C39367 _0457_ _0346_ 0
C39368 _0718_/a_47_47# _0718_/a_285_47# 0.01755f
C39369 VPWR _0546_/a_512_297# 0.00733f
C39370 _0343_ net67 0
C39371 acc0.A\[29\] _1029_/a_975_413# 0
C39372 _0127_ _1029_/a_891_413# 0
C39373 _1011_/a_1059_315# _0726_/a_51_297# 0.00125f
C39374 _1011_/a_27_47# _0726_/a_240_47# 0
C39375 _1011_/a_193_47# _0726_/a_149_47# 0
C39376 pp[27] _0333_ 0.06139f
C39377 _1069_/a_381_47# control0.count\[0\] 0
C39378 _1033_/a_27_47# _1065_/a_466_413# 0
C39379 clknet_1_1__leaf__0460_ _0360_ 0.00327f
C39380 net152 _1043_/a_27_47# 0
C39381 _0081_ _0181_ 0.05607f
C39382 hold11/a_285_47# clknet_1_1__leaf__0457_ 0
C39383 _1052_/a_466_413# _0524_/a_109_297# 0
C39384 clknet_0__0465_ _0088_ 0
C39385 B[11] clknet_1_1__leaf__0464_ 0.0016f
C39386 _0328_ _0320_ 0.03966f
C39387 hold78/a_49_47# _0218_ 0
C39388 _0700_/a_113_47# _0332_ 0.00957f
C39389 net22 net7 0
C39390 clknet_1_1__leaf__0465_ _0350_ 0.03584f
C39391 _1041_/a_466_413# net174 0.00278f
C39392 clkload3/Y acc0.A\[16\] 0.02683f
C39393 net45 _0341_ 0.03249f
C39394 acc0.A\[27\] hold50/a_391_47# 0.04929f
C39395 net125 _1061_/a_1059_315# 0.00152f
C39396 _0398_ _1016_/a_193_47# 0
C39397 _0399_ _1016_/a_27_47# 0
C39398 _0985_/a_193_47# _0195_ 0
C39399 _0384_ acc0.A\[19\] 0
C39400 _0488_ _0487_ 0.00444f
C39401 _0466_ _0485_ 0.03429f
C39402 _0577_/a_109_47# _0183_ 0.00283f
C39403 output38/a_27_47# pp[11] 0.16612f
C39404 _0577_/a_373_47# acc0.A\[22\] 0.00122f
C39405 _0577_/a_27_297# _0120_ 0.10878f
C39406 _0195_ _1018_/a_27_47# 0.44265f
C39407 hold54/a_391_47# control0.sh 0
C39408 _0180_ _0171_ 0.02273f
C39409 _0553_/a_51_297# net171 0.09082f
C39410 net58 _0988_/a_27_47# 0.03928f
C39411 _0640_/a_297_297# clknet_1_1__leaf__0458_ 0
C39412 _1001_/a_381_47# _0346_ 0
C39413 _0467_ _1067_/a_193_47# 0
C39414 _0568_/a_27_297# net209 0.00576f
C39415 _0481_ _1064_/a_1059_315# 0
C39416 hold20/a_391_47# clkload0/a_27_47# 0
C39417 _0181_ _0505_/a_373_47# 0.00122f
C39418 _0645_/a_47_47# _0302_ 0.01433f
C39419 _0663_/a_207_413# VPWR 0.17264f
C39420 net150 net151 0
C39421 _0426_ _0089_ 0
C39422 _0508_/a_81_21# _0345_ 0
C39423 _0563_/a_245_297# _0173_ 0.00149f
C39424 _0579_/a_27_297# clkbuf_0__0457_/a_110_47# 0
C39425 hold58/a_49_47# _1034_/a_193_47# 0
C39426 hold58/a_285_47# _1034_/a_27_47# 0
C39427 _0325_ _0462_ 0
C39428 clknet_1_0__leaf__0463_ net7 0.28635f
C39429 net106 _1015_/a_1059_315# 0
C39430 clknet_1_0__leaf__0462_ _0695_/a_80_21# 0
C39431 _0524_/a_109_297# _0194_ 0.01813f
C39432 _0524_/a_373_47# net12 0
C39433 _0151_ A[7] 0.00484f
C39434 _0693_/a_68_297# _0350_ 0
C39435 net9 _0528_/a_81_21# 0.01201f
C39436 pp[11] _0993_/a_1059_315# 0
C39437 _1065_/a_1059_315# _0160_ 0
C39438 _0129_ _0218_ 0
C39439 net87 net105 0
C39440 _0608_/a_109_297# _0307_ 0
C39441 _0465_ net72 0.00601f
C39442 comp0.B\[12\] _0542_/a_512_297# 0
C39443 _0475_ _0563_/a_240_47# 0.04282f
C39444 net211 _1019_/a_193_47# 0
C39445 _0217_ _0580_/a_109_297# 0.0113f
C39446 _0298_ _0798_/a_113_297# 0.10996f
C39447 net180 input30/a_75_212# 0
C39448 net232 comp0.B\[4\] 0
C39449 clkbuf_1_1__f__0460_/a_110_47# _0332_ 0.0133f
C39450 _0982_/a_891_413# net36 0.04326f
C39451 VPWR hold72/a_391_47# 0.18789f
C39452 _0476_ _1036_/a_27_47# 0
C39453 _0902_/a_27_47# _0352_ 0
C39454 _0431_ acc0.A\[6\] 0
C39455 net45 _1013_/a_891_413# 0.01738f
C39456 hold91/a_49_47# acc0.A\[13\] 0
C39457 _0179_ _1048_/a_891_413# 0
C39458 _0220_ hold61/a_49_47# 0.00537f
C39459 _0664_/a_79_21# _0421_ 0
C39460 _1043_/a_634_159# _1042_/a_193_47# 0.01011f
C39461 _1043_/a_27_47# _1042_/a_466_413# 0
C39462 _1043_/a_193_47# _1042_/a_634_159# 0.01011f
C39463 _1043_/a_466_413# _1042_/a_27_47# 0
C39464 clkbuf_1_1__f__0460_/a_110_47# _0685_/a_68_297# 0.01121f
C39465 _0777_/a_285_47# _0347_ 0.00312f
C39466 hold7/a_285_47# clknet_1_1__leaf__0458_ 0.08245f
C39467 acc0.A\[1\] _0526_/a_27_47# 0
C39468 clkbuf_0__0461_/a_110_47# hold72/a_49_47# 0.02131f
C39469 _0769_/a_384_47# VPWR 0
C39470 net93 acc0.A\[23\] 0
C39471 net17 hold84/a_49_47# 0
C39472 clkbuf_1_1__f__0462_/a_110_47# _0321_ 0.00104f
C39473 _0993_/a_891_413# _0993_/a_975_413# 0.00851f
C39474 _0993_/a_381_47# _0993_/a_561_413# 0.00123f
C39475 clkload1/Y _0218_ 0
C39476 _0280_ _0345_ 0.0837f
C39477 hold87/a_391_47# VPWR 0.1826f
C39478 _0341_ _0587_/a_27_47# 0.0014f
C39479 clknet_0__0463_ _0159_ 0.00111f
C39480 hold85/a_49_47# _0471_ 0
C39481 _0458_ _0255_ 0
C39482 _1039_/a_1059_315# net125 0
C39483 output45/a_27_47# _1013_/a_27_47# 0
C39484 _0742_/a_81_21# _0366_ 0.00419f
C39485 _0258_ _0254_ 0.01744f
C39486 _0238_ _0462_ 0.11265f
C39487 VPWR _0529_/a_109_297# 0.19343f
C39488 _0730_/a_79_21# _0730_/a_297_297# 0.01735f
C39489 _1039_/a_381_47# _0953_/a_32_297# 0
C39490 _0973_/a_373_47# clknet_1_0__leaf__0460_ 0
C39491 _0677_/a_47_47# _0240_ 0.03773f
C39492 _0673_/a_253_47# _0347_ 0.00826f
C39493 _0343_ _0707_/a_201_297# 0.00385f
C39494 hold20/a_285_47# _0981_/a_109_297# 0
C39495 _0677_/a_47_47# _0369_ 0
C39496 _0363_ _0371_ 0
C39497 _0724_/a_199_47# _0333_ 0.00101f
C39498 _0452_ _0350_ 0.00422f
C39499 _0714_/a_51_297# _1031_/a_193_47# 0
C39500 net63 _0830_/a_79_21# 0.02045f
C39501 _0485_ _1064_/a_193_47# 0.00291f
C39502 _0487_ _1064_/a_27_47# 0
C39503 net135 _0196_ 0
C39504 _0549_/a_150_297# _0173_ 0
C39505 _1026_/a_466_413# net112 0
C39506 _1059_/a_1059_315# VPWR 0.41392f
C39507 _1054_/a_1059_315# acc0.A\[5\] 0
C39508 _0985_/a_891_413# _0449_ 0
C39509 _0083_ clknet_1_0__leaf__0458_ 0
C39510 _0465_ _1047_/a_634_159# 0.0046f
C39511 _0234_ _0103_ 0.036f
C39512 _0999_/a_27_47# _0779_/a_215_47# 0
C39513 _1072_/a_27_47# _0486_ 0
C39514 _0472_ _1061_/a_634_159# 0
C39515 _0432_ _0435_ 0
C39516 _0111_ _0567_/a_27_297# 0
C39517 _0817_/a_81_21# _0817_/a_368_297# 0.01485f
C39518 _0181_ _1009_/a_381_47# 0.00393f
C39519 _0402_ _0346_ 0.3051f
C39520 _0383_ _0374_ 0.00112f
C39521 _0312_ _0359_ 0.0944f
C39522 _1024_/a_1017_47# _0122_ 0
C39523 _0542_/a_51_297# net20 0.04123f
C39524 _0081_ _1018_/a_27_47# 0
C39525 _0473_ _0207_ 0
C39526 _0270_ _0345_ 0
C39527 _0537_/a_68_297# _0176_ 0.10435f
C39528 _1021_/a_891_413# _0118_ 0
C39529 _0230_ _0754_/a_149_47# 0.01046f
C39530 _0598_/a_79_21# _0219_ 0.0234f
C39531 _0216_ _0333_ 0.06928f
C39532 clknet_1_1__leaf__0459_ hold70/a_285_47# 0.01576f
C39533 _0645_/a_47_47# net6 0
C39534 _0536_/a_51_297# _1061_/a_27_47# 0
C39535 hold99/a_285_47# pp[11] 0.00222f
C39536 hold36/a_391_47# net184 0.00647f
C39537 _0573_/a_27_47# _0181_ 0.00127f
C39538 _0174_ _1040_/a_466_413# 0.00894f
C39539 net34 _0978_/a_109_297# 0
C39540 _1037_/a_634_159# _1037_/a_1059_315# 0
C39541 _1037_/a_27_47# _1037_/a_381_47# 0.06222f
C39542 _1037_/a_193_47# _1037_/a_891_413# 0.19212f
C39543 hold53/a_285_47# net52 0
C39544 _0469_ clknet_1_1__leaf_clk 0
C39545 _0182_ acc0.A\[3\] 0
C39546 net20 _0142_ 0.12484f
C39547 _0767_/a_145_75# _0462_ 0
C39548 comp0.B\[10\] _1040_/a_891_413# 0.02136f
C39549 _0953_/a_32_297# net174 0.00219f
C39550 _0369_ _0507_/a_109_47# 0
C39551 _0252_ _0186_ 0.03236f
C39552 output59/a_27_47# _1030_/a_27_47# 0
C39553 _0785_/a_384_47# _0401_ 0
C39554 net126 _0137_ 0.0025f
C39555 _0182_ control0.sh 0.09406f
C39556 net67 net38 0
C39557 VPWR _1005_/a_193_47# 0.35241f
C39558 _0790_/a_35_297# acc0.A\[15\] 0.07604f
C39559 _0790_/a_117_297# net42 0.0103f
C39560 _0166_ _0468_ 0.37881f
C39561 _0369_ hold82/a_285_47# 0.03178f
C39562 net120 net186 0.02538f
C39563 _1041_/a_466_413# _1041_/a_592_47# 0.00553f
C39564 _0247_ _0615_/a_109_297# 0.01217f
C39565 VPWR _0991_/a_975_413# 0.00601f
C39566 _0690_/a_68_297# _1008_/a_1059_315# 0
C39567 B[2] B[3] 0
C39568 net22 comp0.B\[11\] 0
C39569 net54 _0737_/a_35_297# 0
C39570 _1054_/a_466_413# _0180_ 0.02636f
C39571 _0504_/a_27_47# net218 0
C39572 hold30/a_285_47# _1023_/a_27_47# 0
C39573 _0172_ net73 0
C39574 VPWR _0600_/a_337_297# 0.0029f
C39575 _1057_/a_27_47# _0189_ 0
C39576 _1057_/a_634_159# net2 0
C39577 hold86/a_285_47# _0843_/a_68_297# 0
C39578 _1038_/a_193_47# net8 0
C39579 _0176_ _1043_/a_381_47# 0
C39580 _0718_/a_129_47# net162 0
C39581 _1030_/a_27_47# _0724_/a_113_297# 0
C39582 _1039_/a_1059_315# _0473_ 0.00199f
C39583 hold9/a_49_47# _1008_/a_193_47# 0.00115f
C39584 acc0.A\[12\] acc0.A\[10\] 0.32983f
C39585 acc0.A\[29\] net114 0
C39586 net175 net10 0
C39587 _0216_ clkbuf_1_0__f__0460_/a_110_47# 0.04059f
C39588 _1051_/a_1059_315# _0193_ 0
C39589 net233 _0345_ 0.04786f
C39590 _0195_ clknet_1_1__leaf__0461_ 0.16793f
C39591 net35 clknet_1_0__leaf_clk 0.00486f
C39592 hold42/a_49_47# net3 0
C39593 _0369_ _0242_ 0.10747f
C39594 _0315_ acc0.A\[24\] 0.19456f
C39595 _0461_ _0585_/a_109_47# 0
C39596 _0216_ _0250_ 0.02522f
C39597 VPWR _1011_/a_1059_315# 0.40634f
C39598 _0292_ hold70/a_285_47# 0
C39599 hold59/a_285_47# _0347_ 0.00108f
C39600 _1055_/a_193_47# net62 0
C39601 hold88/a_49_47# _0190_ 0
C39602 net53 _1024_/a_1059_315# 0
C39603 _1029_/a_193_47# _1008_/a_27_47# 0
C39604 _1029_/a_27_47# _1008_/a_193_47# 0
C39605 _0476_ comp0.B\[3\] 0.04077f
C39606 _0995_/a_27_47# _0400_ 0
C39607 clknet_1_0__leaf__0465_ _0399_ 0
C39608 _0277_ net41 0.32962f
C39609 _0963_/a_35_297# _1069_/a_891_413# 0.01244f
C39610 _0195_ _1030_/a_193_47# 0.04084f
C39611 _0255_ clkbuf_1_1__f__0458_/a_110_47# 0.00825f
C39612 _0230_ _0228_ 0
C39613 net48 _1005_/a_193_47# 0.03864f
C39614 _0644_/a_47_47# _0996_/a_1059_315# 0
C39615 clkbuf_0__0461_/a_110_47# clknet_0__0461_ 1.86296f
C39616 _0135_ net171 0.00482f
C39617 A[10] _0515_/a_384_47# 0
C39618 _0289_ _0089_ 0
C39619 _1019_/a_1059_315# _0345_ 0.01149f
C39620 _0361_ _1009_/a_466_413# 0
C39621 _0985_/a_1059_315# _0846_/a_51_297# 0.01354f
C39622 _0985_/a_27_47# _0846_/a_240_47# 0
C39623 output67/a_27_47# _1058_/a_634_159# 0.0014f
C39624 _0804_/a_79_21# _0994_/a_27_47# 0
C39625 net67 hold81/a_285_47# 0.00548f
C39626 _0182_ net157 0.23141f
C39627 clknet_1_0__leaf__0459_ hold72/a_391_47# 0.03301f
C39628 VPWR _0264_ 0.68721f
C39629 _1012_/a_891_413# _0110_ 0
C39630 _0143_ clknet_0__0464_ 0.02884f
C39631 net22 _0202_ 0
C39632 _0413_ pp[14] 0
C39633 hold33/a_285_47# clknet_0__0463_ 0
C39634 _0275_ _0444_ 0
C39635 _0274_ _0445_ 0
C39636 net213 _0217_ 0
C39637 control0.state\[0\] _0972_/a_93_21# 0.01463f
C39638 _0218_ _0799_/a_209_47# 0.00109f
C39639 _0487_ _1065_/a_193_47# 0
C39640 _0135_ net24 0
C39641 _0324_ _0219_ 0.13959f
C39642 _0689_/a_68_297# _0689_/a_150_297# 0.00477f
C39643 hold26/a_49_47# clknet_1_0__leaf__0465_ 0
C39644 _0146_ _1049_/a_1059_315# 0
C39645 acc0.A\[29\] _0365_ 0
C39646 _0650_/a_68_297# acc0.A\[10\] 0.18009f
C39647 net95 _1009_/a_193_47# 0.00453f
C39648 _0261_ _0263_ 0.93852f
C39649 _0246_ net52 0
C39650 net68 _0345_ 0
C39651 _0960_/a_27_47# _0480_ 0.01342f
C39652 _0661_/a_277_297# _0288_ 0
C39653 pp[7] _0435_ 0
C39654 _0287_ _0656_/a_59_75# 0
C39655 _1003_/a_193_47# acc0.A\[21\] 0
C39656 _0175_ _0562_/a_68_297# 0.10913f
C39657 _0495_/a_150_297# _0171_ 0
C39658 _0098_ _0195_ 0
C39659 _0461_ _0772_/a_297_297# 0
C39660 _0983_/a_381_47# _0264_ 0
C39661 _1027_/a_561_413# net156 0
C39662 _0643_/a_253_47# _0274_ 0.01507f
C39663 _0643_/a_337_297# _0275_ 0.00257f
C39664 net44 _0342_ 0.01276f
C39665 _0606_/a_297_297# _0219_ 0
C39666 comp0.B\[8\] _1040_/a_193_47# 0.08522f
C39667 _0206_ _1040_/a_27_47# 0.42459f
C39668 VPWR net170 0.35512f
C39669 hold97/a_391_47# _0698_/a_113_297# 0
C39670 _1059_/a_1059_315# clknet_1_0__leaf__0459_ 0
C39671 hold76/a_285_47# _0218_ 0.00436f
C39672 _0697_/a_217_297# _0352_ 0
C39673 _0957_/a_32_297# _0957_/a_304_297# 0.00167f
C39674 _0747_/a_510_47# net52 0.00153f
C39675 _0119_ _0891_/a_27_47# 0
C39676 _0749_/a_384_47# _0372_ 0
C39677 _0341_ VPWR 1.39685f
C39678 clknet_1_0__leaf__0462_ _1023_/a_1017_47# 0
C39679 clknet_1_0__leaf__0460_ _0758_/a_79_21# 0.0375f
C39680 _0471_ net17 0.05781f
C39681 VPWR _0845_/a_109_297# 0.00454f
C39682 _1041_/a_27_47# comp0.B\[10\] 0
C39683 _0855_/a_81_21# _1014_/a_193_47# 0
C39684 _0855_/a_299_297# _1014_/a_27_47# 0
C39685 hold23/a_285_47# net71 0.00201f
C39686 _0478_ _1071_/a_891_413# 0
C39687 _1007_/a_634_159# _1007_/a_466_413# 0.23992f
C39688 _1007_/a_193_47# _1007_/a_1059_315# 0.03202f
C39689 _1007_/a_27_47# _1007_/a_891_413# 0.03224f
C39690 _1052_/a_193_47# _1052_/a_381_47# 0.09503f
C39691 _1052_/a_634_159# _1052_/a_891_413# 0.03684f
C39692 _1052_/a_27_47# _1052_/a_561_413# 0.00163f
C39693 net44 _0334_ 0
C39694 _1035_/a_592_47# _0133_ 0.00164f
C39695 _0343_ pp[30] 0.0361f
C39696 _0967_/a_109_93# net33 0
C39697 hold87/a_391_47# _0453_ 0.00139f
C39698 hold10/a_49_47# _0177_ 0
C39699 _1012_/a_1059_315# acc0.A\[30\] 0
C39700 net121 net23 0
C39701 _0195_ _0531_/a_27_297# 0
C39702 net186 _1034_/a_466_413# 0
C39703 _0133_ B[15] 0
C39704 _0973_/a_27_297# hold93/a_391_47# 0
C39705 _1058_/a_466_413# _1058_/a_381_47# 0.03733f
C39706 _1058_/a_193_47# _1058_/a_975_413# 0
C39707 _1058_/a_1059_315# _1058_/a_891_413# 0.31086f
C39708 _0973_/a_109_297# hold93/a_285_47# 0
C39709 _0172_ _1044_/a_27_47# 0.07649f
C39710 _0461_ _0208_ 0.22368f
C39711 _0179_ _1052_/a_27_47# 0.38151f
C39712 hold13/a_49_47# control0.reset 0
C39713 _0570_/a_27_297# _1027_/a_193_47# 0
C39714 net86 _0240_ 0.00468f
C39715 net34 _0480_ 0
C39716 clknet_1_0__leaf__0462_ hold52/a_49_47# 0.00938f
C39717 _1051_/a_1017_47# _0172_ 0.00134f
C39718 clk _0489_ 0
C39719 net86 _0369_ 0
C39720 clknet_0__0458_ _0442_ 0
C39721 _0298_ net41 0
C39722 _0083_ hold18/a_49_47# 0
C39723 _0399_ _0400_ 0.00807f
C39724 _0626_/a_68_297# net62 0.03947f
C39725 _1050_/a_27_47# net154 0.02682f
C39726 _0680_/a_80_21# _0311_ 0.11437f
C39727 _0680_/a_472_297# _0305_ 0.00107f
C39728 hold12/a_391_47# _0487_ 0.01194f
C39729 VPWR _0722_/a_79_21# 0.45761f
C39730 _0559_/a_51_297# _0176_ 0
C39731 acc0.A\[12\] _0510_/a_109_297# 0.0105f
C39732 net47 clknet_1_1__leaf__0458_ 0.00807f
C39733 _0353_ hold62/a_285_47# 0.00146f
C39734 VPWR _0139_ 0.51959f
C39735 _1011_/a_634_159# _0109_ 0.04584f
C39736 _1011_/a_381_47# _0355_ 0
C39737 _1011_/a_891_413# net227 0.00102f
C39738 _1011_/a_561_413# _0354_ 0
C39739 net46 _0222_ 0.03271f
C39740 VPWR _1013_/a_891_413# 0.1845f
C39741 clknet_0__0465_ _0516_/a_109_297# 0
C39742 net36 clkbuf_0__0457_/a_110_47# 0
C39743 _0343_ _0771_/a_215_297# 0
C39744 net119 _1065_/a_193_47# 0
C39745 _1002_/a_466_413# VPWR 0.24815f
C39746 _0949_/a_145_75# clknet_0_clk 0
C39747 _0182_ _1015_/a_975_413# 0
C39748 _0229_ clknet_1_0__leaf__0460_ 0
C39749 _0305_ _0183_ 0.02143f
C39750 _1052_/a_381_47# net12 0.01141f
C39751 hold75/a_391_47# _0849_/a_79_21# 0.00134f
C39752 _0983_/a_27_47# _0854_/a_215_47# 0
C39753 _0742_/a_81_21# acc0.A\[24\] 0.01257f
C39754 _0538_/a_512_297# comp0.B\[14\] 0.00178f
C39755 _0174_ _0465_ 0
C39756 _0328_ _1007_/a_1059_315# 0
C39757 _1058_/a_27_47# _0186_ 0.00459f
C39758 _0176_ input29/a_75_212# 0
C39759 _0327_ _0727_/a_109_47# 0
C39760 acc0.A\[9\] _0990_/a_891_413# 0.00407f
C39761 _0254_ net72 0
C39762 hold13/a_391_47# net24 0
C39763 _0128_ net209 0.23816f
C39764 hold70/a_49_47# _0418_ 0
C39765 hold70/a_391_47# _0281_ 0
C39766 VPWR _0525_/a_81_21# 0.22718f
C39767 _0575_/a_373_47# _0216_ 0.00121f
C39768 pp[18] _0340_ 0.00916f
C39769 _1021_/a_1059_315# acc0.A\[20\] 0
C39770 _0974_/a_222_93# _0974_/a_448_47# 0.00596f
C39771 _0258_ _0625_/a_59_75# 0
C39772 net205 _1034_/a_891_413# 0
C39773 clknet_1_0__leaf__0462_ clknet_1_0__leaf__0460_ 0.13895f
C39774 net47 _0263_ 0
C39775 net76 _0399_ 0.02155f
C39776 clknet_0__0458_ net165 0
C39777 _0984_/a_466_413# VPWR 0.25097f
C39778 clkbuf_0__0458_/a_110_47# _0842_/a_59_75# 0.00575f
C39779 _0985_/a_891_413# _0260_ 0
C39780 net167 _0481_ 0
C39781 _0746_/a_299_297# _0359_ 0.06532f
C39782 _0994_/a_891_413# _0218_ 0.003f
C39783 net59 _1012_/a_975_413# 0
C39784 comp0.B\[12\] _0141_ 0.11031f
C39785 net111 _1026_/a_466_413# 0
C39786 _0995_/a_975_413# pp[14] 0
C39787 _0501_/a_27_47# VPWR 0.23901f
C39788 _0570_/a_27_297# _1026_/a_1059_315# 0
C39789 net168 net14 0.00675f
C39790 _0369_ _0990_/a_27_47# 0
C39791 _0217_ _0583_/a_27_297# 0.09814f
C39792 _0343_ _0302_ 0
C39793 clkbuf_1_0__f__0462_/a_110_47# _1007_/a_193_47# 0.00675f
C39794 _1002_/a_466_413# net48 0
C39795 VPWR _1042_/a_561_413# 0.00221f
C39796 _0251_ _0642_/a_215_297# 0.01581f
C39797 _0776_/a_27_47# _0347_ 0
C39798 net58 _0267_ 0.02485f
C39799 _0343_ _0795_/a_299_297# 0
C39800 _1056_/a_891_413# acc0.A\[9\] 0
C39801 _0544_/a_245_297# _0202_ 0
C39802 _0982_/a_1059_315# _0346_ 0
C39803 _0518_/a_109_47# _0252_ 0
C39804 _0195_ _0855_/a_299_297# 0.00179f
C39805 _0316_ _0219_ 0.00216f
C39806 control0.sh _0495_/a_68_297# 0.12706f
C39807 output55/a_27_47# VPWR 0.30803f
C39808 _0691_/a_68_297# _0315_ 0.17796f
C39809 output54/a_27_47# net155 0
C39810 pp[26] _0572_/a_373_47# 0
C39811 _1043_/a_193_47# net128 0
C39812 clknet_1_1__leaf__0464_ _0140_ 0
C39813 net141 net74 0
C39814 _0998_/a_891_413# net83 0
C39815 _0217_ _0603_/a_68_297# 0
C39816 _0305_ acc0.A\[15\] 0.03616f
C39817 _1030_/a_1059_315# acc0.A\[30\] 0.13354f
C39818 _0273_ _0989_/a_634_159# 0
C39819 _0988_/a_634_159# _0988_/a_381_47# 0
C39820 hold3/a_391_47# _0219_ 0
C39821 _0347_ _0219_ 0.30566f
C39822 acc0.A\[12\] _0188_ 0
C39823 clkbuf_0_clk/a_110_47# _1062_/a_27_47# 0
C39824 _0730_/a_215_47# _0108_ 0
C39825 hold64/a_391_47# acc0.A\[19\] 0.03198f
C39826 net1 _0383_ 0
C39827 _0465_ _0208_ 0
C39828 VPWR _0532_/a_81_21# 0.21325f
C39829 _0343_ _0339_ 1.03886f
C39830 net10 _1043_/a_1017_47# 0
C39831 hold20/a_391_47# _0170_ 0
C39832 _0695_/a_300_47# _0326_ 0
C39833 _0312_ _0325_ 0
C39834 net225 _1031_/a_193_47# 0
C39835 _0496_/a_27_47# _0494_/a_27_47# 0
C39836 _1056_/a_27_47# _0369_ 0
C39837 _0104_ _0219_ 0.00132f
C39838 hold38/a_49_47# net231 0
C39839 _1026_/a_1017_47# acc0.A\[26\] 0
C39840 _0328_ clkbuf_1_0__f__0462_/a_110_47# 0
C39841 _1001_/a_1059_315# clknet_1_0__leaf__0457_ 0.01021f
C39842 net85 _0779_/a_79_21# 0.0015f
C39843 _0999_/a_466_413# _0097_ 0.00167f
C39844 _0460_ _1062_/a_193_47# 0
C39845 clknet_0__0457_ _0855_/a_81_21# 0
C39846 _0472_ net147 0.03287f
C39847 _0346_ _0451_ 0.02249f
C39848 clknet_1_1__leaf__0460_ _1009_/a_1017_47# 0
C39849 _0331_ hold95/a_391_47# 0
C39850 net17 control0.reset 0
C39851 _1035_/a_1059_315# net27 0
C39852 _1021_/a_193_47# clknet_1_0__leaf__0457_ 0.01213f
C39853 _0316_ _1008_/a_634_159# 0
C39854 _0455_ net104 0
C39855 _0453_ _0264_ 0.34349f
C39856 input6/a_75_212# pp[13] 0
C39857 net47 clknet_1_0__leaf__0461_ 0.00289f
C39858 _0191_ _0087_ 0
C39859 _0458_ _0843_/a_68_297# 0
C39860 pp[26] acc0.A\[27\] 0.12329f
C39861 hold36/a_391_47# net130 0
C39862 net44 output59/a_27_47# 0.03959f
C39863 _0279_ _0994_/a_466_413# 0
C39864 _0795_/a_81_21# net5 0.04858f
C39865 clknet_1_1__leaf__0460_ _0741_/a_109_297# 0.00413f
C39866 _0792_/a_209_297# _0219_ 0.01013f
C39867 net43 net42 0.9449f
C39868 clkbuf_1_1__f__0463_/a_110_47# clknet_0__0463_ 0.43882f
C39869 _0347_ _1008_/a_634_159# 0.00231f
C39870 _0174_ net174 0.03071f
C39871 _0399_ _0849_/a_510_47# 0.00166f
C39872 _1037_/a_466_413# _0135_ 0.03882f
C39873 _0745_/a_109_47# _0219_ 0
C39874 _0531_/a_27_297# _1048_/a_193_47# 0
C39875 _0531_/a_109_297# _1048_/a_27_47# 0
C39876 pp[0] input30/a_75_212# 0
C39877 VPWR net37 0.8826f
C39878 _0195_ _0998_/a_561_413# 0.00115f
C39879 hold38/a_49_47# hold38/a_285_47# 0.22264f
C39880 _0238_ _0312_ 0.00637f
C39881 clknet_1_0__leaf__0462_ _0576_/a_109_297# 0.00729f
C39882 pp[30] _1030_/a_381_47# 0.00628f
C39883 clkbuf_1_0__f__0465_/a_110_47# _0826_/a_27_53# 0.00864f
C39884 net191 _0345_ 0.00454f
C39885 _0305_ _0179_ 0.23913f
C39886 _0557_/a_51_297# control0.sh 0.0139f
C39887 hold89/a_49_47# _1064_/a_1059_315# 0
C39888 _0999_/a_27_47# net42 0
C39889 _0343_ net6 0
C39890 net8 net29 0
C39891 _0207_ comp0.B\[8\] 0
C39892 net171 _0206_ 0.00183f
C39893 hold24/a_285_47# _0209_ 0.00123f
C39894 VPWR hold91/a_49_47# 0.27016f
C39895 _0985_/a_466_413# _0448_ 0
C39896 _0959_/a_472_297# net23 0
C39897 net169 _0180_ 0.03941f
C39898 _0218_ _0668_/a_79_21# 0.00714f
C39899 net88 clknet_1_1__leaf_clk 0
C39900 pp[8] _0186_ 0.00338f
C39901 _1001_/a_634_159# _1001_/a_381_47# 0
C39902 _0604_/a_113_47# _0248_ 0
C39903 _0183_ _0181_ 0.29488f
C39904 net221 _1060_/a_193_47# 0
C39905 _0101_ net51 0.00278f
C39906 _1035_/a_27_47# input25/a_75_212# 0
C39907 _1062_/a_634_159# _1062_/a_1059_315# 0
C39908 _1062_/a_27_47# _1062_/a_381_47# 0.06222f
C39909 _1062_/a_193_47# _1062_/a_891_413# 0.1932f
C39910 VPWR _0385_ 0.17147f
C39911 net125 _0472_ 0.00395f
C39912 _0340_ _0567_/a_109_47# 0
C39913 _1011_/a_193_47# _0725_/a_209_297# 0
C39914 _1021_/a_27_47# _1021_/a_634_159# 0.14145f
C39915 _0587_/a_27_47# acc0.A\[30\] 0
C39916 _0831_/a_35_297# _0253_ 0.09566f
C39917 _0608_/a_27_47# clkbuf_1_1__f__0461_/a_110_47# 0
C39918 _1003_/a_634_159# net49 0
C39919 net61 _0626_/a_150_297# 0.00108f
C39920 control0.add _0610_/a_59_75# 0
C39921 _0575_/a_109_297# _1024_/a_466_413# 0
C39922 hold41/a_49_47# hold41/a_391_47# 0.00188f
C39923 _0419_ _0807_/a_150_297# 0
C39924 net64 _0827_/a_27_47# 0.00219f
C39925 clkbuf_1_1__f__0465_/a_110_47# _0425_ 0
C39926 _0275_ _0424_ 0
C39927 _0467_ _0951_/a_109_93# 0
C39928 _0198_ net9 0.07303f
C39929 _0146_ net175 0.25439f
C39930 _1049_/a_891_413# _1048_/a_891_413# 0
C39931 net189 net3 0
C39932 _0248_ _0603_/a_68_297# 0
C39933 _0996_/a_27_47# _0670_/a_79_21# 0.00686f
C39934 VPWR _1006_/a_1017_47# 0
C39935 _0248_ hold73/a_391_47# 0
C39936 _0285_ _0787_/a_303_47# 0
C39937 _1000_/a_891_413# _0217_ 0
C39938 _0346_ _0373_ 0.19781f
C39939 _0536_/a_51_297# _0953_/a_32_297# 0
C39940 _0963_/a_285_297# _0167_ 0
C39941 _0963_/a_285_47# clknet_1_0__leaf_clk 0
C39942 hold88/a_49_47# _0346_ 0
C39943 hold47/a_285_47# _0143_ 0.00297f
C39944 _0331_ acc0.A\[28\] 0.01735f
C39945 input4/a_75_212# net37 0
C39946 hold4/a_285_47# net51 0
C39947 _0856_/a_79_21# VPWR 0.43751f
C39948 control0.state\[0\] _0975_/a_59_75# 0.04508f
C39949 clknet_1_1__leaf__0464_ _1043_/a_634_159# 0.04454f
C39950 VPWR _0986_/a_1017_47# 0
C39951 _0195_ _1015_/a_27_47# 0
C39952 _0749_/a_81_21# acc0.A\[19\] 0
C39953 hold52/a_391_47# _0352_ 0
C39954 net180 _0176_ 0.05461f
C39955 net45 _0779_/a_79_21# 0.00412f
C39956 _0742_/a_384_47# _0368_ 0.0012f
C39957 VPWR _0670_/a_297_297# 0.0081f
C39958 _1020_/a_193_47# _0721_/a_27_47# 0.00875f
C39959 acc0.A\[13\] _0184_ 0
C39960 _0951_/a_109_93# comp0.B\[0\] 0.02512f
C39961 _0092_ _0994_/a_193_47# 0.22714f
C39962 hold55/a_49_47# _0461_ 0
C39963 _0130_ _0891_/a_27_47# 0
C39964 net44 _0240_ 0.52445f
C39965 hold34/a_391_47# _0179_ 0
C39966 _0186_ _0988_/a_891_413# 0
C39967 _0373_ hold94/a_49_47# 0
C39968 _1004_/a_561_413# _0216_ 0
C39969 _0850_/a_68_297# _0635_/a_27_47# 0
C39970 net44 _0369_ 0
C39971 _0714_/a_51_297# _0344_ 0.09849f
C39972 hold78/a_285_47# _0714_/a_240_47# 0
C39973 _0149_ _0150_ 0
C39974 _0676_/a_113_47# net43 0
C39975 control0.state\[0\] net231 0.23055f
C39976 _0361_ _0315_ 0.09098f
C39977 _0181_ acc0.A\[15\] 0.12477f
C39978 net48 _0385_ 0.19953f
C39979 _1072_/a_466_413# _1068_/a_891_413# 0
C39980 _1072_/a_381_47# _1068_/a_634_159# 0
C39981 _1072_/a_1059_315# _1068_/a_1059_315# 0
C39982 VPWR _0762_/a_215_47# 0.00167f
C39983 _0251_ _0833_/a_510_47# 0
C39984 _0219_ hold95/a_49_47# 0.01299f
C39985 hold13/a_285_47# _1037_/a_1059_315# 0.00197f
C39986 net99 net60 0
C39987 _0174_ clknet_0__0464_ 0.00225f
C39988 output44/a_27_47# _0335_ 0
C39989 _0346_ _0271_ 0.10921f
C39990 net185 _1062_/a_27_47# 0
C39991 _0102_ net52 0.00772f
C39992 hold30/a_391_47# clknet_1_0__leaf__0460_ 0.00114f
C39993 _0399_ clkbuf_0__0459_/a_110_47# 0.00101f
C39994 _0179_ _0510_/a_27_297# 0.00621f
C39995 net154 _0987_/a_27_47# 0.00182f
C39996 _1036_/a_193_47# net122 0.00707f
C39997 _1036_/a_466_413# clknet_1_1__leaf__0463_ 0.01239f
C39998 _0457_ _0782_/a_27_47# 0.02861f
C39999 _1052_/a_27_47# hold83/a_49_47# 0.01463f
C40000 _1050_/a_27_47# clknet_0__0464_ 0
C40001 net187 _0713_/a_27_47# 0.00647f
C40002 _0738_/a_68_297# net244 0.12849f
C40003 _0461_ _1019_/a_193_47# 0.03916f
C40004 _0538_/a_240_47# _1046_/a_891_413# 0
C40005 _0815_/a_113_297# _0345_ 0.04785f
C40006 net160 _1034_/a_891_413# 0
C40007 _0749_/a_81_21# _0249_ 0
C40008 _0956_/a_32_297# _0563_/a_51_297# 0.00112f
C40009 _1035_/a_592_47# _0208_ 0
C40010 hold67/a_49_47# hold67/a_285_47# 0.22264f
C40011 _1041_/a_193_47# net153 0.28645f
C40012 _0087_ clkbuf_1_0__f__0465_/a_110_47# 0
C40013 _1041_/a_634_159# net127 0
C40014 _1047_/a_466_413# _1047_/a_561_413# 0.00772f
C40015 _1047_/a_634_159# _1047_/a_975_413# 0
C40016 clknet_1_1__leaf__0459_ net81 0.13062f
C40017 _0185_ net229 0.05764f
C40018 net83 _0793_/a_240_47# 0.00128f
C40019 _0305_ _0780_/a_35_297# 0.01988f
C40020 hold39/a_285_47# clknet_1_1__leaf_clk 0
C40021 _0473_ _0472_ 0.33717f
C40022 _0714_/a_149_47# net163 0
C40023 control0.state\[1\] hold38/a_49_47# 0
C40024 _0131_ _0563_/a_512_297# 0
C40025 _1041_/a_1059_315# _0136_ 0
C40026 _0639_/a_109_297# _0465_ 0
C40027 net185 _0561_/a_51_297# 0.09296f
C40028 hold85/a_285_47# _1063_/a_27_47# 0
C40029 _0343_ _0718_/a_47_47# 0.00994f
C40030 _0216_ _0526_/a_27_47# 0.07838f
C40031 net58 _0833_/a_510_47# 0.00116f
C40032 _0183_ _1018_/a_27_47# 0.01055f
C40033 _0217_ _1018_/a_634_159# 0.01328f
C40034 _0456_ _1014_/a_1059_315# 0.00281f
C40035 _0797_/a_297_47# net5 0
C40036 _1007_/a_466_413# net93 0
C40037 _1007_/a_634_159# _0105_ 0
C40038 net243 _1004_/a_634_159# 0.01849f
C40039 VPWR _0454_ 0.17577f
C40040 _0837_/a_368_297# _0441_ 0.01665f
C40041 _0837_/a_266_47# _0440_ 0.04268f
C40042 _0165_ hold93/a_391_47# 0.01483f
C40043 _1020_/a_975_413# _0352_ 0.00108f
C40044 _0293_ _0369_ 0
C40045 acc0.A\[25\] net50 0
C40046 _0126_ _1027_/a_193_47# 0
C40047 net190 _1027_/a_1059_315# 0
C40048 net48 _0762_/a_215_47# 0.00244f
C40049 _1021_/a_381_47# clknet_1_0__leaf__0461_ 0
C40050 input19/a_75_212# _0203_ 0
C40051 VPWR _0498_/a_240_47# 0.0026f
C40052 clknet_1_1__leaf__0460_ _0678_/a_150_297# 0
C40053 hold74/a_285_47# hold74/a_391_47# 0.41909f
C40054 _0212_ net121 0
C40055 net185 _0133_ 0.03023f
C40056 _0234_ hold66/a_49_47# 0
C40057 acc0.A\[4\] _0527_/a_27_297# 0
C40058 _0179_ _0181_ 0.20199f
C40059 hold32/a_285_47# pp[1] 0
C40060 _0971_/a_81_21# _0163_ 0.11458f
C40061 _0971_/a_384_47# _0181_ 0.01003f
C40062 A[14] net6 0.00552f
C40063 _0574_/a_109_47# net52 0
C40064 net97 _0109_ 0.00435f
C40065 net57 _0355_ 0.03535f
C40066 _0195_ _0354_ 0.08145f
C40067 _0225_ _0383_ 0
C40068 _0172_ _0196_ 0
C40069 VPWR _0505_/a_27_297# 0.23811f
C40070 _0294_ _0582_/a_373_47# 0
C40071 _0100_ VPWR 0.33298f
C40072 clknet_1_0__leaf__0461_ _0173_ 0
C40073 _0558_/a_68_297# net185 0.17637f
C40074 _1061_/a_381_47# comp0.B\[9\] 0
C40075 _1057_/a_27_47# net67 0.03297f
C40076 _0459_ _0796_/a_215_47# 0
C40077 pp[15] net41 0.01455f
C40078 _0328_ net51 0
C40079 clkbuf_1_1__f__0460_/a_110_47# clknet_0__0460_ 0.31131f
C40080 acc0.A\[4\] hold1/a_391_47# 0.02501f
C40081 _0464_ _0180_ 0
C40082 _0243_ _0247_ 0.05457f
C40083 _0329_ _0356_ 0.06532f
C40084 _0283_ net37 0.10267f
C40085 _0983_/a_466_413# _0081_ 0.00716f
C40086 _0983_/a_381_47# _0454_ 0
C40087 _0983_/a_891_413# _0455_ 0
C40088 net69 _0854_/a_79_21# 0
C40089 _0143_ comp0.B\[14\] 0.1746f
C40090 _0323_ _0370_ 0.00295f
C40091 net36 _0350_ 0.04047f
C40092 _1063_/a_1059_315# _1063_/a_891_413# 0.31086f
C40093 _1063_/a_193_47# _1063_/a_975_413# 0
C40094 _1063_/a_466_413# _1063_/a_381_47# 0.03733f
C40095 _0833_/a_79_21# _0988_/a_27_47# 0.00172f
C40096 _0555_/a_240_47# net171 0
C40097 _0965_/a_47_47# _1072_/a_27_47# 0.05847f
C40098 _1019_/a_381_47# _0346_ 0.00546f
C40099 _0362_ _0328_ 0
C40100 hold75/a_49_47# clknet_1_0__leaf__0458_ 0.00121f
C40101 _1037_/a_381_47# _0208_ 0
C40102 net159 _1063_/a_891_413# 0
C40103 _0959_/a_80_21# _0959_/a_217_297# 0.12661f
C40104 acc0.A\[20\] net223 0
C40105 _1063_/a_1017_47# clknet_1_0__leaf__0457_ 0
C40106 _0251_ net63 0.09437f
C40107 _0462_ _1006_/a_891_413# 0.0043f
C40108 net36 _0463_ 0.01573f
C40109 _0165_ control0.reset 0
C40110 _0748_/a_81_21# _0748_/a_384_47# 0.00138f
C40111 _0137_ net8 0.51144f
C40112 _1039_/a_975_413# _0177_ 0
C40113 hold11/a_285_47# net135 0
C40114 hold11/a_49_47# _0147_ 0
C40115 net158 _1049_/a_561_413# 0
C40116 _0343_ _0790_/a_285_297# 0.00883f
C40117 _1028_/a_27_47# net113 0
C40118 _1028_/a_634_159# clknet_1_1__leaf__0462_ 0.0242f
C40119 net64 net16 0.00816f
C40120 _0356_ _0221_ 0.02926f
C40121 _0663_/a_207_413# _0345_ 0.01188f
C40122 _0211_ _0209_ 0
C40123 VPWR _0506_/a_81_21# 0.23055f
C40124 net46 _0771_/a_298_297# 0
C40125 _0642_/a_215_297# _0831_/a_285_297# 0
C40126 control0.count\[3\] _1071_/a_634_159# 0
C40127 _0483_ _1071_/a_27_47# 0
C40128 _0733_/a_79_199# _0368_ 0
C40129 _0176_ _0545_/a_150_297# 0
C40130 _0490_ _0482_ 0
C40131 _0515_/a_81_21# net66 0.01072f
C40132 clknet_1_0__leaf__0463_ net123 0.10497f
C40133 _1011_/a_592_47# acc0.A\[29\] 0
C40134 hold18/a_285_47# _0266_ 0.00212f
C40135 _0337_ _0333_ 0.01455f
C40136 _0217_ _0114_ 0
C40137 VPWR _1010_/a_634_159# 0.20276f
C40138 _1000_/a_27_47# _1000_/a_634_159# 0.13646f
C40139 _0100_ net48 0.23776f
C40140 _0576_/a_373_47# _0352_ 0
C40141 VPWR acc0.A\[30\] 1.27392f
C40142 _1060_/a_1059_315# _1060_/a_891_413# 0.31086f
C40143 _1060_/a_193_47# _1060_/a_975_413# 0
C40144 _1060_/a_466_413# _1060_/a_381_47# 0.03733f
C40145 net198 net20 0.049f
C40146 _0733_/a_448_47# _0319_ 0.00273f
C40147 acc0.A\[28\] _1008_/a_27_47# 0
C40148 clkbuf_0__0457_/a_110_47# hold60/a_391_47# 0.01103f
C40149 _0294_ clknet_1_0__leaf__0461_ 0
C40150 hold48/a_49_47# net18 0
C40151 hold49/a_49_47# hold49/a_391_47# 0.00188f
C40152 _0192_ _0520_/a_27_297# 0.11183f
C40153 net45 _0239_ 0.00453f
C40154 _0462_ _0616_/a_78_199# 0.00257f
C40155 _1053_/a_466_413# net11 0.0017f
C40156 _0143_ _1050_/a_381_47# 0
C40157 _1039_/a_1059_315# _0555_/a_149_47# 0
C40158 hold69/a_285_47# clkbuf_0__0460_/a_110_47# 0
C40159 net203 _1065_/a_466_413# 0
C40160 VPWR _0846_/a_51_297# 0.50624f
C40161 hold26/a_285_47# _0176_ 0.00606f
C40162 clknet_1_1__leaf__0463_ comp0.B\[6\] 0.04853f
C40163 clkbuf_1_1__f__0462_/a_110_47# _0332_ 0.00486f
C40164 _0988_/a_381_47# net74 0
C40165 _0269_ _0826_/a_219_297# 0
C40166 _0553_/a_149_47# _0174_ 0.02197f
C40167 _1067_/a_891_413# clknet_1_1__leaf_clk 0
C40168 _0399_ _0986_/a_193_47# 0.03171f
C40169 _0661_/a_27_297# _0817_/a_81_21# 0
C40170 _0973_/a_109_297# _1063_/a_27_47# 0
C40171 _0973_/a_27_297# _1063_/a_193_47# 0
C40172 control0.state\[0\] control0.state\[1\] 0.39002f
C40173 VPWR _1009_/a_466_413# 0.24729f
C40174 _0698_/a_113_297# _0698_/a_199_47# 0
C40175 _0579_/a_109_297# net187 0.01052f
C40176 _0467_ _0486_ 0.00129f
C40177 hold19/a_49_47# hold19/a_391_47# 0.00188f
C40178 _0156_ net143 0
C40179 _0280_ _0809_/a_299_297# 0
C40180 _1041_/a_381_47# _0206_ 0
C40181 net53 _0368_ 0
C40182 _0235_ _0603_/a_68_297# 0.12525f
C40183 _0152_ acc0.A\[6\] 0
C40184 _0982_/a_1017_47# _0465_ 0
C40185 _0195_ _0452_ 0.00187f
C40186 _0233_ _0756_/a_285_47# 0
C40187 _0218_ net47 0.7184f
C40188 _0234_ acc0.A\[22\] 0
C40189 _0583_/a_27_297# _0583_/a_373_47# 0.01338f
C40190 _1071_/a_27_47# control0.count\[1\] 0
C40191 VPWR _1014_/a_975_413# 0.00461f
C40192 _1071_/a_891_413# VPWR 0.20416f
C40193 _0973_/a_27_297# _0460_ 0.01068f
C40194 _0459_ _0775_/a_79_21# 0
C40195 net195 net19 0.39016f
C40196 _0195_ _0567_/a_27_297# 0.15514f
C40197 _0289_ net229 0
C40198 _0985_/a_193_47# _0179_ 0.04226f
C40199 net8 comp0.B\[6\] 0
C40200 _0856_/a_510_47# _0452_ 0
C40201 hold39/a_391_47# VPWR 0.18826f
C40202 acc0.A\[15\] _0507_/a_373_47# 0
C40203 _0780_/a_35_297# _0181_ 0.0141f
C40204 _0500_/a_27_47# _1049_/a_466_413# 0
C40205 _1059_/a_27_47# _0219_ 0
C40206 _1021_/a_1017_47# _0460_ 0
C40207 clknet_0__0458_ _0832_/a_113_47# 0
C40208 comp0.B\[13\] clknet_0__0464_ 0
C40209 acc0.A\[15\] hold82/a_391_47# 0.00265f
C40210 _0573_/a_27_47# _1015_/a_27_47# 0
C40211 comp0.B\[9\] net174 0.02301f
C40212 hold20/a_391_47# net35 0.01562f
C40213 _1067_/a_381_47# clkbuf_1_1__f_clk/a_110_47# 0
C40214 _0739_/a_79_21# _0318_ 0
C40215 clknet_0__0464_ _1046_/a_193_47# 0.19239f
C40216 clkbuf_0__0464_/a_110_47# _1046_/a_381_47# 0.00121f
C40217 _1071_/a_193_47# clkbuf_1_0__f_clk/a_110_47# 0.00826f
C40218 _0183_ clknet_1_1__leaf__0461_ 0.00473f
C40219 net226 clknet_1_0__leaf_clk 0.14269f
C40220 _1008_/a_1059_315# _0365_ 0
C40221 net54 _1027_/a_193_47# 0.03467f
C40222 _1008_/a_634_159# _0106_ 0.04794f
C40223 _0959_/a_217_297# _0173_ 0
C40224 VPWR _0954_/a_32_297# 0.41198f
C40225 _0558_/a_150_297# net27 0.00159f
C40226 _0305_ clkload3/a_110_47# 0
C40227 _0347_ net94 0
C40228 _0678_/a_68_297# clkbuf_1_1__f__0461_/a_110_47# 0
C40229 _0458_ _0257_ 0
C40230 _0718_/a_285_47# _1030_/a_466_413# 0
C40231 net9 _1048_/a_466_413# 0.01533f
C40232 _0151_ net11 0
C40233 comp0.B\[11\] _1043_/a_193_47# 0
C40234 comp0.B\[12\] _1043_/a_27_47# 0
C40235 output57/a_27_47# acc0.A\[29\] 0.00285f
C40236 VPWR B[5] 0.27284f
C40237 _1020_/a_27_47# _0578_/a_27_297# 0
C40238 pp[8] net62 0
C40239 net243 net46 0.00102f
C40240 _0276_ _0300_ 0.06915f
C40241 clkbuf_1_0__f__0459_/a_110_47# net6 0
C40242 _0538_/a_149_47# _1045_/a_1059_315# 0
C40243 _0538_/a_240_47# _1045_/a_466_413# 0
C40244 _0201_ _1045_/a_27_47# 0
C40245 net149 _1047_/a_1059_315# 0
C40246 clknet_1_0__leaf__0465_ _0527_/a_109_297# 0
C40247 hold13/a_285_47# _0472_ 0.0144f
C40248 hold13/a_49_47# _0475_ 0
C40249 VPWR _1022_/a_1059_315# 0.38685f
C40250 clknet_1_0__leaf__0465_ _0346_ 0.08409f
C40251 pp[30] _0568_/a_27_297# 0.00495f
C40252 net23 _0178_ 0.00134f
C40253 clknet_1_1__leaf__0460_ _0305_ 0.12596f
C40254 _0349_ clknet_1_1__leaf__0460_ 0
C40255 _0553_/a_149_47# _0208_ 0
C40256 VPWR _0779_/a_79_21# 0.45527f
C40257 clknet_1_1__leaf__0459_ _0993_/a_466_413# 0
C40258 _0852_/a_35_297# _0452_ 0.07102f
C40259 _0610_/a_59_75# _0610_/a_145_75# 0.00658f
C40260 _0993_/a_891_413# net38 0.00629f
C40261 input22/a_75_212# hold6/a_391_47# 0
C40262 _0999_/a_634_159# _0999_/a_466_413# 0.23992f
C40263 _0999_/a_193_47# _0999_/a_1059_315# 0.03405f
C40264 _0999_/a_27_47# _0999_/a_891_413# 0.03224f
C40265 _0820_/a_215_47# _0401_ 0
C40266 net17 _1063_/a_193_47# 0.03506f
C40267 _0992_/a_193_47# _0422_ 0
C40268 _0992_/a_634_159# net217 0
C40269 _0083_ _0448_ 0
C40270 _1017_/a_1059_315# net221 0.00158f
C40271 _1001_/a_193_47# net223 0.01299f
C40272 _1001_/a_27_47# _0391_ 0.00189f
C40273 clknet_1_0__leaf__0465_ net65 0
C40274 VPWR _0310_ 1.35058f
C40275 _0340_ _1031_/a_193_47# 0
C40276 _0555_/a_51_297# _0957_/a_32_297# 0.0018f
C40277 _0478_ _0975_/a_59_75# 0
C40278 _1004_/a_27_47# _0217_ 0
C40279 _0991_/a_975_413# _0345_ 0
C40280 net120 _1034_/a_466_413# 0
C40281 _0115_ _1060_/a_561_413# 0
C40282 hold86/a_285_47# _0263_ 0
C40283 control0.count\[3\] _0978_/a_27_297# 0
C40284 _1062_/a_466_413# _0160_ 0.00106f
C40285 net17 _0460_ 0.08714f
C40286 clknet_0__0458_ _0622_/a_109_47# 0
C40287 output56/a_27_47# net208 0
C40288 acc0.A\[12\] _0647_/a_285_47# 0.03533f
C40289 clknet_1_0__leaf__0465_ _0935_/a_27_47# 0
C40290 _0600_/a_337_297# _0345_ 0
C40291 clknet_1_0__leaf__0465_ _1061_/a_193_47# 0.00102f
C40292 _0691_/a_68_297# _0691_/a_150_297# 0.00477f
C40293 _1021_/a_381_47# _1021_/a_561_413# 0.00123f
C40294 _1021_/a_891_413# _1021_/a_975_413# 0.00851f
C40295 net89 net49 0
C40296 hold24/a_391_47# _1038_/a_1059_315# 0
C40297 hold24/a_285_47# _1038_/a_891_413# 0.00152f
C40298 _0454_ _0453_ 0.01682f
C40299 _0575_/a_109_297# _0122_ 0.00169f
C40300 _0081_ _0452_ 0
C40301 _0591_/a_109_297# clknet_1_0__leaf__0460_ 0
C40302 _0308_ _0350_ 0
C40303 acc0.A\[3\] _1048_/a_1059_315# 0
C40304 clknet_0__0459_ net229 0
C40305 _0180_ _0830_/a_79_21# 0
C40306 acc0.A\[16\] _0096_ 0
C40307 hold41/a_285_47# net4 0
C40308 clknet_1_1__leaf__0461_ acc0.A\[15\] 0
C40309 _0729_/a_68_297# _0352_ 0.01968f
C40310 _0179_ hold82/a_391_47# 0.03411f
C40311 _0174_ _0536_/a_51_297# 0.11188f
C40312 clknet_1_1__leaf__0459_ _0790_/a_35_297# 0
C40313 VPWR _0540_/a_245_297# 0.00614f
C40314 clknet_0__0464_ _0987_/a_27_47# 0
C40315 _0996_/a_193_47# _0302_ 0
C40316 acc0.A\[31\] net60 0.34495f
C40317 _0459_ _0158_ 0
C40318 clkbuf_1_1__f__0462_/a_110_47# _0738_/a_68_297# 0
C40319 comp0.B\[5\] _0560_/a_68_297# 0.01724f
C40320 _0098_ _0183_ 0
C40321 hold43/a_391_47# net115 0
C40322 hold43/a_285_47# net191 0.00276f
C40323 _1056_/a_634_159# acc0.A\[12\] 0
C40324 _0369_ _0829_/a_109_297# 0
C40325 _0457_ net17 0.23312f
C40326 net62 _0988_/a_891_413# 0.02057f
C40327 _1043_/a_193_47# _0202_ 0
C40328 VPWR net173 0.2706f
C40329 net40 net42 0.0024f
C40330 _1011_/a_27_47# _0219_ 0.01792f
C40331 hold11/a_391_47# VPWR 0.17188f
C40332 clknet_1_0__leaf__0459_ _0506_/a_81_21# 0
C40333 clknet_1_1__leaf__0464_ net129 0.31906f
C40334 net132 _1061_/a_891_413# 0
C40335 net157 net7 0
C40336 comp0.B\[10\] _0547_/a_150_297# 0
C40337 _0953_/a_304_297# _0206_ 0
C40338 _0817_/a_368_297# _0426_ 0
C40339 _0384_ _0462_ 0.02941f
C40340 _0673_/a_103_199# acc0.A\[9\] 0
C40341 net1 clkbuf_1_1__f__0457_/a_110_47# 0.00344f
C40342 _0728_/a_59_75# _1011_/a_27_47# 0.00255f
C40343 VPWR _0978_/a_373_47# 0
C40344 _0168_ _0978_/a_109_297# 0.0021f
C40345 hold26/a_391_47# _0139_ 0
C40346 clknet_1_0__leaf__0464_ _1046_/a_27_47# 0
C40347 hold19/a_391_47# _1017_/a_193_47# 0
C40348 hold19/a_49_47# _1017_/a_466_413# 0
C40349 clknet_1_0__leaf__0458_ net71 0.18075f
C40350 clknet_1_0__leaf__0465_ _0538_/a_149_47# 0
C40351 control0.count\[2\] _1071_/a_193_47# 0.16628f
C40352 _0984_/a_891_413# _0399_ 0
C40353 net225 _0344_ 0.00185f
C40354 _1055_/a_634_159# _0189_ 0
C40355 _0210_ _0209_ 0
C40356 clknet_0__0464_ comp0.B\[9\] 0
C40357 hold37/a_49_47# _0143_ 0.29946f
C40358 hold47/a_49_47# _1050_/a_193_47# 0.00148f
C40359 _0561_/a_240_47# _0132_ 0
C40360 VPWR _1067_/a_381_47# 0.07807f
C40361 _0264_ _0345_ 0.35499f
C40362 _0222_ _1023_/a_193_47# 0.00443f
C40363 acc0.A\[12\] _0806_/a_113_297# 0.01779f
C40364 _1050_/a_1059_315# _0186_ 0
C40365 _0725_/a_209_297# _0707_/a_75_199# 0
C40366 hold31/a_285_47# VPWR 0.28386f
C40367 net17 _1062_/a_891_413# 0
C40368 hold28/a_285_47# hold28/a_391_47# 0.41909f
C40369 hold99/a_391_47# net38 0.07739f
C40370 _1033_/a_1059_315# clknet_1_0__leaf__0461_ 0.01273f
C40371 pp[9] input2/a_75_212# 0
C40372 acc0.A\[21\] _0460_ 0.05644f
C40373 pp[27] acc0.A\[29\] 0.02025f
C40374 _0276_ _0404_ 0.03113f
C40375 _0324_ _1007_/a_193_47# 0
C40376 _0382_ clknet_1_0__leaf__0460_ 0
C40377 net58 _0347_ 0.02615f
C40378 _0459_ _0391_ 0
C40379 _0179_ _0187_ 0.01239f
C40380 _0618_/a_79_21# _0249_ 0.11245f
C40381 net186 _0175_ 0.18366f
C40382 net161 clknet_1_1__leaf__0463_ 0.32037f
C40383 _0346_ _0400_ 0.00117f
C40384 _0226_ acc0.A\[20\] 0.18788f
C40385 _0343_ _0275_ 0.07911f
C40386 _0416_ _0787_/a_209_297# 0
C40387 hold14/a_285_47# net27 0
C40388 VPWR _1027_/a_27_47# 0.65831f
C40389 input27/a_75_212# net27 0.10859f
C40390 _0314_ _0219_ 0.00216f
C40391 _1041_/a_592_47# comp0.B\[9\] 0
C40392 _0257_ clkbuf_1_1__f__0458_/a_110_47# 0
C40393 hold100/a_285_47# _0850_/a_68_297# 0
C40394 _0350_ _1008_/a_381_47# 0
C40395 _1047_/a_561_413# _0145_ 0
C40396 _1000_/a_27_47# _0242_ 0
C40397 _1003_/a_1059_315# _0760_/a_285_47# 0
C40398 _0997_/a_27_47# _0405_ 0.0011f
C40399 hold46/a_49_47# _0174_ 0
C40400 output55/a_27_47# net56 0.00592f
C40401 _0707_/a_201_297# _0128_ 0
C40402 _0339_ _0568_/a_27_297# 0.00263f
C40403 output51/a_27_47# net51 0.21401f
C40404 _0459_ _0581_/a_27_297# 0.0148f
C40405 clknet_0__0458_ acc0.A\[3\] 0
C40406 net168 net63 0.00736f
C40407 clknet_0__0465_ _0434_ 0.00324f
C40408 net157 _1048_/a_1059_315# 0
C40409 _0343_ hold74/a_49_47# 0.01023f
C40410 acc0.A\[14\] _0459_ 0.21779f
C40411 net185 _0208_ 0.0179f
C40412 net170 _0345_ 0
C40413 _0343_ _0311_ 0
C40414 VPWR _0768_/a_27_47# 0.00744f
C40415 _0557_/a_51_297# _1036_/a_891_413# 0.00713f
C40416 clknet_1_1__leaf__0463_ net26 0.09249f
C40417 _0546_/a_51_297# _1040_/a_634_159# 0
C40418 _0341_ _0345_ 0.02288f
C40419 _0710_/a_109_47# _0219_ 0.00239f
C40420 _0217_ net104 0.03246f
C40421 _0567_/a_373_47# acc0.A\[30\] 0
C40422 _0476_ net24 0.05589f
C40423 net232 _0959_/a_217_297# 0
C40424 hold85/a_49_47# _0470_ 0
C40425 net93 _0105_ 0.00173f
C40426 net55 _0730_/a_79_21# 0.05091f
C40427 _0513_/a_384_47# net4 0
C40428 _0513_/a_81_21# _0187_ 0
C40429 acc0.A\[8\] _0989_/a_193_47# 0.03472f
C40430 acc0.A\[8\] hold1/a_285_47# 0
C40431 _0753_/a_297_297# _0374_ 0
C40432 _0200_ _0472_ 0
C40433 _0311_ net95 0
C40434 clknet_1_0__leaf__0457_ _0246_ 0
C40435 net44 hold15/a_285_47# 0.01553f
C40436 _0328_ _0324_ 0.7989f
C40437 clkload3/a_110_47# _0181_ 0
C40438 _0996_/a_193_47# net6 0
C40439 A[1] net171 0
C40440 _0291_ _0992_/a_27_47# 0
C40441 _0712_/a_297_297# _0340_ 0.05525f
C40442 pp[0] _0176_ 0
C40443 _0487_ _0880_/a_27_47# 0
C40444 _0544_/a_51_297# _0544_/a_240_47# 0.03076f
C40445 net61 _0831_/a_35_297# 0
C40446 _0531_/a_27_297# acc0.A\[15\] 0
C40447 _0535_/a_68_297# comp0.B\[14\] 0.17558f
C40448 _0956_/a_304_297# control0.reset 0
C40449 _0376_ net213 0
C40450 _0747_/a_297_297# _0460_ 0.00172f
C40451 _0472_ comp0.B\[8\] 0.00187f
C40452 VPWR _0524_/a_109_297# 0.18998f
C40453 _1034_/a_634_159# _1034_/a_1059_315# 0
C40454 _1034_/a_27_47# _1034_/a_381_47# 0.05658f
C40455 _1034_/a_193_47# _1034_/a_891_413# 0.19524f
C40456 _0536_/a_245_297# _0536_/a_240_47# 0
C40457 _0581_/a_109_297# clknet_1_0__leaf__0461_ 0.00158f
C40458 net76 _0346_ 0
C40459 _0796_/a_79_21# net238 0.11962f
C40460 net162 _1030_/a_891_413# 0
C40461 clknet_1_1__leaf__0460_ _0181_ 0.06531f
C40462 _1021_/a_466_413# acc0.A\[21\] 0
C40463 _0679_/a_68_297# _0462_ 0
C40464 net168 _1053_/a_891_413# 0.01274f
C40465 _0559_/a_149_47# hold58/a_391_47# 0
C40466 VPWR _0972_/a_93_21# 0.13536f
C40467 VPWR _0184_ 0.37265f
C40468 _0626_/a_150_297# _0269_ 0
C40469 _0464_ _0498_/a_51_297# 0
C40470 _0239_ VPWR 0.47882f
C40471 _0428_ net66 0.03476f
C40472 _0427_ acc0.A\[8\] 0.00457f
C40473 _0982_/a_561_413# clknet_1_0__leaf__0461_ 0
C40474 acc0.A\[20\] clkbuf_0__0457_/a_110_47# 0
C40475 _0183_ _0855_/a_299_297# 0
C40476 _1013_/a_193_47# _0219_ 0.02057f
C40477 _0516_/a_373_47# acc0.A\[9\] 0
C40478 clknet_1_0__leaf__0459_ _0310_ 0
C40479 control0.state\[0\] _1066_/a_634_159# 0
C40480 _0570_/a_27_297# _0570_/a_373_47# 0.01338f
C40481 _0343_ _0583_/a_27_297# 0.02124f
C40482 net45 _0309_ 0
C40483 _0086_ _0988_/a_193_47# 0.18109f
C40484 _1063_/a_381_47# _0161_ 0.13197f
C40485 _0225_ _0756_/a_129_47# 0.0011f
C40486 _0231_ _0692_/a_113_47# 0
C40487 _0607_/a_109_297# _0219_ 0
C40488 net34 _1068_/a_27_47# 0
C40489 control0.state\[0\] _1068_/a_634_159# 0
C40490 control0.state\[1\] _1068_/a_193_47# 0
C40491 _0129_ _0710_/a_109_297# 0
C40492 VPWR _1026_/a_466_413# 0.27212f
C40493 _0483_ _1072_/a_634_159# 0
C40494 _0848_/a_109_297# _0848_/a_27_47# 0
C40495 control0.count\[3\] _1072_/a_1059_315# 0.14735f
C40496 output35/a_27_47# pp[21] 0
C40497 net78 _0992_/a_1059_315# 0
C40498 _0750_/a_27_47# net51 0.00338f
C40499 _0724_/a_199_47# acc0.A\[29\] 0
C40500 acc0.A\[14\] _0265_ 0.00405f
C40501 VPWR _1024_/a_561_413# 0.00306f
C40502 hold32/a_49_47# hold32/a_391_47# 0.00188f
C40503 _0399_ hold91/a_391_47# 0.02842f
C40504 _0218_ _0848_/a_109_297# 0
C40505 _0517_/a_299_297# _0517_/a_384_47# 0
C40506 _0174_ comp0.B\[14\] 0.17263f
C40507 _0999_/a_193_47# _0397_ 0
C40508 _0361_ _0691_/a_150_297# 0
C40509 hold97/a_391_47# VPWR 0.17419f
C40510 net46 net151 0
C40511 net248 acc0.A\[6\] 0
C40512 acc0.A\[17\] net43 0.52433f
C40513 _0294_ _0218_ 0.31989f
C40514 VPWR _1048_/a_592_47# 0
C40515 net18 _0203_ 0.18756f
C40516 _0204_ net19 0
C40517 control0.state\[1\] _0478_ 0
C40518 clknet_1_0__leaf__0460_ _1005_/a_634_159# 0.01117f
C40519 A[10] _0186_ 0
C40520 net114 clknet_1_1__leaf__0462_ 0.14465f
C40521 _0967_/a_109_93# _1062_/a_27_47# 0
C40522 _1017_/a_27_47# _1017_/a_1059_315# 0.04864f
C40523 _1017_/a_193_47# _1017_/a_466_413# 0.07911f
C40524 _0487_ _1062_/a_27_47# 0.03385f
C40525 net58 clkbuf_0__0465_/a_110_47# 0.04617f
C40526 _0259_ _0271_ 0
C40527 hold47/a_49_47# net194 0
C40528 _0473_ _1046_/a_891_413# 0.01976f
C40529 _0216_ acc0.A\[29\] 0.3629f
C40530 _0179_ _0531_/a_27_297# 0.01192f
C40531 _1004_/a_891_413# _0122_ 0
C40532 VPWR net96 0.4839f
C40533 _1000_/a_381_47# _1000_/a_561_413# 0.00123f
C40534 _1000_/a_27_47# net86 0.23437f
C40535 _1000_/a_891_413# _1000_/a_975_413# 0.00851f
C40536 _0507_/a_27_297# _0507_/a_109_47# 0.00393f
C40537 _0600_/a_253_47# clknet_1_0__leaf__0460_ 0.00338f
C40538 _1033_/a_1017_47# clknet_1_0__leaf__0457_ 0
C40539 _1060_/a_381_47# _0158_ 0.13437f
C40540 _0477_ _1063_/a_27_47# 0
C40541 _1051_/a_891_413# net11 0.01899f
C40542 _0195_ _0398_ 0.01539f
C40543 _0129_ _1013_/a_27_47# 0
C40544 _0176_ hold51/a_391_47# 0.00134f
C40545 _0168_ _0480_ 0
C40546 _0671_/a_199_47# acc0.A\[15\] 0.0109f
C40547 _0428_ _0350_ 0
C40548 _1072_/a_561_413# VPWR 0.00243f
C40549 net126 net174 0
C40550 _0143_ acc0.A\[4\] 0.0587f
C40551 net36 clkbuf_1_0__f__0463_/a_110_47# 0
C40552 clkbuf_0__0463_/a_110_47# _1061_/a_466_413# 0
C40553 _0462_ _0383_ 0
C40554 clknet_1_1__leaf__0458_ _0987_/a_975_413# 0
C40555 _0786_/a_472_297# net228 0.00137f
C40556 _0174_ _0543_/a_68_297# 0.04199f
C40557 comp0.B\[10\] net153 0
C40558 _0536_/a_51_297# _1046_/a_193_47# 0.00227f
C40559 output55/a_27_47# _0345_ 0.00238f
C40560 _0520_/a_27_297# clknet_1_0__leaf__0465_ 0.03208f
C40561 _0293_ _0817_/a_81_21# 0.17085f
C40562 _0292_ _0817_/a_266_47# 0
C40563 _0289_ _0817_/a_368_297# 0
C40564 _0165_ _1063_/a_193_47# 0
C40565 net240 _1063_/a_1059_315# 0
C40566 clkbuf_1_1__f__0461_/a_110_47# _0675_/a_68_297# 0.01503f
C40567 _0216_ _0699_/a_68_297# 0
C40568 _0582_/a_109_297# _0347_ 0
C40569 _0317_ _0330_ 0.08496f
C40570 acc0.A\[11\] acc0.A\[10\] 0.0439f
C40571 _0290_ _0992_/a_27_47# 0
C40572 _0347_ _1007_/a_193_47# 0.00592f
C40573 net9 net148 0.37175f
C40574 clknet_1_0__leaf__0460_ _1006_/a_27_47# 0.01734f
C40575 _0857_/a_27_47# net119 0
C40576 _0963_/a_35_297# _0481_ 0.17423f
C40577 _0231_ _0618_/a_79_21# 0.04283f
C40578 _0751_/a_29_53# clknet_1_0__leaf__0460_ 0.00308f
C40579 _0548_/a_51_297# _0545_/a_68_297# 0
C40580 net53 clknet_0__0460_ 0
C40581 clknet_1_0__leaf__0465_ clkbuf_0__0464_/a_110_47# 0.02934f
C40582 hold55/a_285_47# _0457_ 0.02023f
C40583 _0583_/a_373_47# _0114_ 0
C40584 _0165_ _0460_ 0.03958f
C40585 _1072_/a_27_47# clknet_0_clk 0.05102f
C40586 _1050_/a_634_159# _1050_/a_1059_315# 0
C40587 _1050_/a_27_47# _1050_/a_381_47# 0.06222f
C40588 _1050_/a_193_47# _1050_/a_891_413# 0.19497f
C40589 _0643_/a_253_297# VPWR 0.00207f
C40590 VPWR _0315_ 0.74893f
C40591 _1019_/a_1059_315# clknet_1_0__leaf__0457_ 0.04561f
C40592 _0557_/a_149_47# comp0.B\[5\] 0.00208f
C40593 output47/a_27_47# VPWR 0.46506f
C40594 hold50/a_285_47# hold50/a_391_47# 0.41909f
C40595 _1032_/a_1059_315# control0.reset 0
C40596 clkbuf_0__0463_/a_110_47# net24 0
C40597 _0294_ _0775_/a_215_47# 0.00284f
C40598 clknet_1_1__leaf__0462_ _0365_ 0.06519f
C40599 _0221_ _1011_/a_891_413# 0.00739f
C40600 _0958_/a_27_47# _0958_/a_197_47# 0.00167f
C40601 hold21/a_391_47# acc0.A\[7\] 0.02564f
C40602 _0179_ _1049_/a_592_47# 0.00124f
C40603 _1051_/a_891_413# hold7/a_391_47# 0.00107f
C40604 _0427_ _0423_ 0
C40605 _0177_ _0173_ 0
C40606 _0316_ _0328_ 0.00957f
C40607 _0565_/a_51_297# _0565_/a_245_297# 0.01218f
C40608 clknet_1_0__leaf__0462_ hold90/a_285_47# 0.00134f
C40609 _0715_/a_27_47# _0350_ 0
C40610 _0458_ _0263_ 0.00175f
C40611 _0718_/a_129_47# VPWR 0
C40612 _0998_/a_634_159# net43 0.00125f
C40613 clknet_1_0__leaf__0459_ _0768_/a_27_47# 0
C40614 _0457_ _0165_ 0
C40615 _0748_/a_299_297# _0246_ 0
C40616 _1054_/a_27_47# _1052_/a_466_413# 0
C40617 net94 _0106_ 0.00849f
C40618 _0559_/a_240_47# _0134_ 0
C40619 net224 _1009_/a_1059_315# 0.00651f
C40620 _0328_ _0347_ 0
C40621 _0982_/a_193_47# net149 0
C40622 _1039_/a_27_47# _0463_ 0.02954f
C40623 _1039_/a_466_413# clkbuf_0__0463_/a_110_47# 0
C40624 net150 VPWR 1.01408f
C40625 _1056_/a_193_47# _0179_ 0.39535f
C40626 net46 _0378_ 0.00561f
C40627 acc0.A\[14\] _1060_/a_381_47# 0
C40628 hold65/a_285_47# hold65/a_391_47# 0.41909f
C40629 _1020_/a_891_413# net187 0.00665f
C40630 pp[28] _0725_/a_303_47# 0
C40631 net25 _0561_/a_240_47# 0.05778f
C40632 hold46/a_49_47# comp0.B\[13\] 0.30527f
C40633 net248 _0624_/a_59_75# 0
C40634 net1 _0486_ 0
C40635 _0486_ _1068_/a_381_47# 0.01755f
C40636 _0143_ _1045_/a_891_413# 0
C40637 hold58/a_49_47# _1036_/a_1059_315# 0
C40638 _0531_/a_373_47# clknet_1_1__leaf__0457_ 0
C40639 _0606_/a_465_297# _0460_ 0
C40640 net37 _0345_ 0.0038f
C40641 hold46/a_285_47# _1046_/a_27_47# 0
C40642 hold46/a_49_47# _1046_/a_193_47# 0
C40643 pp[30] _0128_ 0.00652f
C40644 _0946_/a_184_297# clk 0
C40645 output47/a_27_47# output62/a_27_47# 0.00151f
C40646 clknet_1_0__leaf__0463_ _0209_ 0
C40647 _0343_ _1000_/a_891_413# 0.00108f
C40648 pp[12] _0218_ 0.0058f
C40649 _0137_ _0492_/a_27_47# 0
C40650 _1033_/a_891_413# _0173_ 0
C40651 acc0.A\[10\] hold81/a_391_47# 0
C40652 _0183_ _1015_/a_27_47# 0
C40653 acc0.A\[19\] _0242_ 0.05764f
C40654 clkbuf_1_1__f__0459_/a_110_47# acc0.A\[15\] 0.05881f
C40655 _0999_/a_466_413# net85 0.00131f
C40656 net239 _0352_ 0.02642f
C40657 _1001_/a_466_413# _1019_/a_891_413# 0.00388f
C40658 _0487_ net107 0
C40659 hold76/a_285_47# clkbuf_1_0__f__0461_/a_110_47# 0.02333f
C40660 _0772_/a_79_21# _0391_ 0.12553f
C40661 clknet_1_0__leaf__0459_ _0184_ 0
C40662 VPWR _0993_/a_561_413# 0.0036f
C40663 _1054_/a_891_413# net148 0
C40664 net172 net7 0
C40665 _1016_/a_27_47# net221 0.42477f
C40666 _0239_ clknet_1_0__leaf__0459_ 0
C40667 clknet_1_0__leaf__0462_ _1007_/a_561_413# 0.00164f
C40668 comp0.B\[7\] net29 0.00159f
C40669 _0697_/a_300_47# _0321_ 0
C40670 _0256_ _0186_ 0
C40671 hold91/a_49_47# _0345_ 0.02337f
C40672 _0983_/a_891_413# _0217_ 0
C40673 _0775_/a_79_21# _0775_/a_510_47# 0.00844f
C40674 _0775_/a_297_297# _0775_/a_215_47# 0
C40675 _0186_ _0987_/a_1059_315# 0
C40676 _0195_ _0353_ 0.00352f
C40677 _0536_/a_51_297# comp0.B\[9\] 0.01198f
C40678 acc0.A\[1\] hold60/a_49_47# 0
C40679 hold74/a_391_47# net45 0.00261f
C40680 _0133_ net119 0
C40681 _0556_/a_68_297# _1036_/a_466_413# 0.00123f
C40682 hold20/a_49_47# hold20/a_285_47# 0.22264f
C40683 B[9] net198 0
C40684 acc0.A\[14\] _0267_ 0.14374f
C40685 hold38/a_49_47# _0564_/a_68_297# 0.01017f
C40686 _0818_/a_109_47# _0291_ 0.00113f
C40687 comp0.B\[1\] net23 0.04374f
C40688 hold32/a_49_47# _0153_ 0.29658f
C40689 _1033_/a_193_47# net17 0.00103f
C40690 _0961_/a_113_297# _0486_ 0
C40691 _1016_/a_634_159# _0459_ 0.00221f
C40692 hold88/a_49_47# _0253_ 0
C40693 _0648_/a_205_297# _0278_ 0.00272f
C40694 _0648_/a_27_297# _0280_ 0.10255f
C40695 _0343_ hold65/a_49_47# 0.00125f
C40696 pp[8] _0512_/a_109_47# 0
C40697 clknet_1_1__leaf__0460_ _1012_/a_193_47# 0.00109f
C40698 net150 net48 0.08959f
C40699 hold17/a_391_47# net164 0.13552f
C40700 _0598_/a_79_21# _0750_/a_27_47# 0.01104f
C40701 _1051_/a_891_413# clknet_1_1__leaf__0458_ 0
C40702 hold38/a_49_47# clknet_1_1__leaf_clk 0
C40703 _0249_ _0242_ 0
C40704 clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ 1.72358f
C40705 net231 clkbuf_1_1__f_clk/a_110_47# 0.03397f
C40706 _1006_/a_381_47# _0219_ 0
C40707 _0814_/a_109_47# acc0.A\[9\] 0
C40708 _0482_ control0.count\[0\] 0
C40709 _0258_ _0350_ 0
C40710 net64 net142 0
C40711 _0614_/a_29_53# _0245_ 0.09443f
C40712 _0856_/a_79_21# _0345_ 0.11851f
C40713 _0510_/a_109_297# acc0.A\[11\] 0
C40714 hold100/a_49_47# hold100/a_391_47# 0.00188f
C40715 _0985_/a_466_413# _0985_/a_381_47# 0.03733f
C40716 _0985_/a_193_47# _0985_/a_975_413# 0
C40717 _0985_/a_1059_315# _0985_/a_891_413# 0.31086f
C40718 _0304_ _0288_ 0
C40719 acc0.A\[22\] hold29/a_391_47# 0.00107f
C40720 _0183_ hold29/a_285_47# 0
C40721 comp0.B\[13\] comp0.B\[14\] 0.84171f
C40722 hold19/a_285_47# net103 0.00623f
C40723 _1018_/a_193_47# _1018_/a_381_47# 0.09503f
C40724 _1018_/a_634_159# _1018_/a_891_413# 0.03684f
C40725 _1018_/a_27_47# _1018_/a_561_413# 0.00163f
C40726 net36 _1014_/a_27_47# 0
C40727 _0794_/a_326_47# net6 0
C40728 _0985_/a_193_47# _1049_/a_891_413# 0
C40729 _0243_ _0217_ 0
C40730 comp0.B\[14\] _1046_/a_193_47# 0
C40731 net50 _1022_/a_381_47# 0
C40732 _0642_/a_298_297# _0273_ 0.04879f
C40733 VPWR control0.add 2.14753f
C40734 _0982_/a_193_47# _0982_/a_466_413# 0.07482f
C40735 _0982_/a_27_47# _0982_/a_1059_315# 0.04875f
C40736 VPWR _0742_/a_81_21# 0.22875f
C40737 _0725_/a_80_21# _0339_ 0
C40738 _0725_/a_209_47# _0335_ 0
C40739 _1049_/a_27_47# _1049_/a_466_413# 0.27314f
C40740 _1049_/a_193_47# _1049_/a_634_159# 0.11072f
C40741 _0250_ clkbuf_1_0__f__0460_/a_110_47# 0.02188f
C40742 _0983_/a_466_413# acc0.A\[15\] 0.0021f
C40743 clknet_1_1__leaf__0460_ _0732_/a_209_47# 0.00207f
C40744 _0119_ net17 0
C40745 net105 _0869_/a_27_47# 0
C40746 output37/a_27_47# input3/a_75_212# 0
C40747 _1060_/a_1059_315# net228 0
C40748 VPWR _0689_/a_150_297# 0.00115f
C40749 _0753_/a_381_47# _0233_ 0.00969f
C40750 _0753_/a_297_297# _0231_ 0.05011f
C40751 _0172_ _0540_/a_51_297# 0.14467f
C40752 _0552_/a_68_297# _0552_/a_150_297# 0.00477f
C40753 clkload3/a_110_47# clknet_1_1__leaf__0461_ 0
C40754 _0690_/a_68_297# _0690_/a_150_297# 0.00477f
C40755 _1054_/a_193_47# A[8] 0
C40756 _1019_/a_466_413# _0586_/a_27_47# 0
C40757 hold46/a_49_47# comp0.B\[9\] 0
C40758 hold11/a_285_47# _0172_ 0.00549f
C40759 _1038_/a_891_413# _0210_ 0
C40760 clknet_1_0__leaf__0462_ clknet_0__0462_ 0.00292f
C40761 hold56/a_391_47# net23 0
C40762 _1066_/a_27_47# _1066_/a_466_413# 0.27314f
C40763 _1066_/a_193_47# _1066_/a_634_159# 0.12497f
C40764 hold37/a_49_47# _1050_/a_27_47# 0
C40765 _0331_ _1010_/a_27_47# 0
C40766 net56 _1010_/a_634_159# 0
C40767 net56 acc0.A\[30\] 0
C40768 _0183_ clknet_1_1__leaf__0465_ 0
C40769 net45 _0999_/a_466_413# 0.00653f
C40770 VPWR _0309_ 0.34717f
C40771 VPWR _1052_/a_1059_315# 0.403f
C40772 _0833_/a_79_21# _0833_/a_510_47# 0.00844f
C40773 _0833_/a_297_297# _0833_/a_215_47# 0
C40774 _1031_/a_634_159# acc0.A\[30\] 0
C40775 _0339_ _0128_ 0.02795f
C40776 clknet_1_1__leaf__0460_ clknet_1_1__leaf__0461_ 0.00242f
C40777 _1023_/a_27_47# _1022_/a_1059_315# 0
C40778 output67/a_27_47# A[11] 0.03346f
C40779 _0967_/a_297_297# clk 0
C40780 _1068_/a_27_47# _1068_/a_466_413# 0.26005f
C40781 _1068_/a_193_47# _1068_/a_634_159# 0.11897f
C40782 net8 _1040_/a_466_413# 0
C40783 _0459_ _0116_ 0.01191f
C40784 clk _0162_ 0.05824f
C40785 _0294_ _0359_ 0
C40786 _0677_/a_129_47# acc0.A\[17\] 0
C40787 net32 _1040_/a_466_413# 0
C40788 VPWR input22/a_75_212# 0.26942f
C40789 _1019_/a_592_47# clknet_1_0__leaf__0461_ 0
C40790 net178 pp[4] 0
C40791 clkbuf_1_1__f__0464_/a_110_47# _1045_/a_466_413# 0
C40792 net157 clkbuf_1_1__f__0457_/a_110_47# 0.02071f
C40793 net187 _0891_/a_27_47# 0
C40794 _0982_/a_1059_315# _0446_ 0
C40795 hold58/a_391_47# comp0.B\[5\] 0.00962f
C40796 _0731_/a_81_21# _0346_ 0.00885f
C40797 _0255_ _0825_/a_68_297# 0
C40798 pp[9] _0512_/a_109_297# 0.0452f
C40799 _0797_/a_27_413# _0297_ 0.20915f
C40800 _0804_/a_510_47# _0279_ 0.00245f
C40801 _0720_/a_150_297# _0350_ 0
C40802 _1032_/a_634_159# net23 0
C40803 net36 hold18/a_391_47# 0
C40804 net48 control0.add 0
C40805 _0223_ acc0.A\[23\] 0.08774f
C40806 VPWR _0975_/a_59_75# 0.20908f
C40807 _0818_/a_109_47# _0290_ 0
C40808 _0344_ _0340_ 0.09492f
C40809 hold78/a_391_47# _0342_ 0
C40810 hold53/a_49_47# hold53/a_391_47# 0.00188f
C40811 _0544_/a_512_297# _0140_ 0
C40812 _0219_ _0360_ 0.06605f
C40813 _0471_ _0468_ 0.63712f
C40814 _0519_/a_81_21# acc0.A\[7\] 0.03901f
C40815 _0519_/a_299_297# net65 0
C40816 _0357_ _0352_ 0.01362f
C40817 _0108_ _0347_ 0.23435f
C40818 _0625_/a_145_75# net63 0
C40819 _0313_ _0318_ 0.00534f
C40820 net101 clknet_0__0457_ 0.00236f
C40821 acc0.A\[10\] _0281_ 0.12392f
C40822 _0268_ _0261_ 0.12059f
C40823 _1051_/a_193_47# _0186_ 0.03354f
C40824 _1034_/a_27_47# comp0.B\[2\] 0.43399f
C40825 _0557_/a_512_297# net26 0.00124f
C40826 hold6/a_285_47# net198 0
C40827 _0188_ acc0.A\[11\] 0.12559f
C40828 output65/a_27_47# net65 0.22757f
C40829 _0410_ _0094_ 0
C40830 _0119_ acc0.A\[21\] 0
C40831 net14 net139 0.03713f
C40832 net25 B[4] 0.00146f
C40833 B[2] net27 0.13945f
C40834 _0440_ _0433_ 0.11234f
C40835 VPWR net231 0.26381f
C40836 _1056_/a_27_47# hold32/a_49_47# 0
C40837 _0480_ _0976_/a_439_47# 0
C40838 _0169_ _0976_/a_505_21# 0
C40839 _0979_/a_27_297# _0466_ 0.19564f
C40840 _0979_/a_109_297# _0488_ 0.0056f
C40841 _0461_ net202 0.00236f
C40842 _0181_ _0171_ 0
C40843 _0390_ control0.add 0.03335f
C40844 net36 _0195_ 0.16359f
C40845 _0789_/a_544_297# net6 0.00499f
C40846 hold89/a_285_47# control0.count\[0\] 0
C40847 net197 net190 0.51881f
C40848 _0225_ _0618_/a_79_21# 0.04879f
C40849 _0228_ _0369_ 0.02607f
C40850 control0.state\[0\] clknet_1_1__leaf_clk 0.0259f
C40851 _0570_/a_373_47# _0126_ 0
C40852 _0343_ _0114_ 0.04418f
C40853 _0343_ _0615_/a_109_297# 0
C40854 _0534_/a_81_21# _1047_/a_466_413# 0.00453f
C40855 clknet_1_1__leaf__0465_ acc0.A\[15\] 0.0391f
C40856 _0346_ _1006_/a_193_47# 0.46579f
C40857 hold57/a_49_47# comp0.B\[6\] 0.30159f
C40858 hold57/a_285_47# comp0.B\[5\] 0
C40859 comp0.B\[14\] comp0.B\[9\] 0.00135f
C40860 acc0.A\[20\] _0350_ 0
C40861 _0446_ _0451_ 0.00263f
C40862 _0292_ _0181_ 0.08732f
C40863 _0344_ _1013_/a_381_47# 0.00124f
C40864 _0255_ _0841_/a_79_21# 0
C40865 _1001_/a_891_413# _0352_ 0.00143f
C40866 _0793_/a_240_47# _0406_ 0
C40867 pp[30] _1031_/a_1059_315# 0.00463f
C40868 _0422_ _0420_ 0
C40869 _0346_ _0986_/a_193_47# 0
C40870 _1032_/a_27_47# clknet_1_0__leaf__0461_ 0.04189f
C40871 _0999_/a_193_47# _0793_/a_51_297# 0
C40872 pp[15] _1013_/a_975_413# 0
C40873 clknet_0_clk _0972_/a_584_47# 0
C40874 clkbuf_1_0__f__0464_/a_110_47# _1046_/a_27_47# 0
C40875 _1071_/a_561_413# _0466_ 0
C40876 net21 B[13] 0.00552f
C40877 _0716_/a_27_47# _0671_/a_113_297# 0
C40878 _0183_ _0452_ 0
C40879 net117 clknet_1_1__leaf__0462_ 0.12817f
C40880 _0389_ _0372_ 0
C40881 _0243_ _0248_ 0
C40882 _0993_/a_381_47# _0286_ 0
C40883 hold38/a_285_47# VPWR 0.29711f
C40884 net81 _0995_/a_381_47# 0
C40885 hold77/a_391_47# _1009_/a_1059_315# 0.01554f
C40886 clknet_1_0__leaf__0460_ net91 0.27997f
C40887 _1050_/a_381_47# _0987_/a_27_47# 0
C40888 _0172_ _0524_/a_27_297# 0
C40889 _1050_/a_27_47# _0987_/a_381_47# 0
C40890 _1017_/a_891_413# _1017_/a_1017_47# 0.00617f
C40891 _1017_/a_634_159# net103 0.02387f
C40892 _0751_/a_29_53# hold94/a_285_47# 0.00155f
C40893 _0708_/a_68_297# net60 0.11126f
C40894 _1058_/a_1059_315# net3 0
C40895 _1017_/a_27_47# _1016_/a_27_47# 0
C40896 net16 _0369_ 0
C40897 _1052_/a_592_47# net9 0.00255f
C40898 _0429_ _0621_/a_285_297# 0
C40899 acc0.A\[8\] _0988_/a_27_47# 0
C40900 VPWR clknet_1_1__leaf__0457_ 2.22184f
C40901 pp[2] _0253_ 0.00197f
C40902 comp0.B\[7\] _0137_ 0.09562f
C40903 net187 _0346_ 0
C40904 net103 _1060_/a_1017_47# 0
C40905 _0679_/a_68_297# _0312_ 0
C40906 control0.state\[1\] clkbuf_1_1__f_clk/a_110_47# 0.02858f
C40907 _0507_/a_109_47# _0185_ 0
C40908 _0543_/a_68_297# comp0.B\[9\] 0
C40909 _1000_/a_561_413# net45 0
C40910 control0.state\[0\] _0479_ 0
C40911 net125 comp0.B\[15\] 0
C40912 _0804_/a_510_47# _0416_ 0.00134f
C40913 hold82/a_285_47# _0185_ 0
C40914 acc0.A\[30\] _0345_ 0.06217f
C40915 _0476_ _0561_/a_149_47# 0
C40916 output56/a_27_47# _0221_ 0
C40917 net36 _0852_/a_35_297# 0
C40918 _0521_/a_81_21# net230 0.05769f
C40919 _0521_/a_299_297# _0192_ 0.08337f
C40920 _0200_ _1046_/a_891_413# 0.00796f
C40921 _1033_/a_1059_315# _1033_/a_891_413# 0.31086f
C40922 _1033_/a_193_47# _1033_/a_975_413# 0
C40923 _1033_/a_466_413# _1033_/a_381_47# 0.03733f
C40924 hold36/a_391_47# _0142_ 0
C40925 _0758_/a_510_47# net51 0
C40926 _1012_/a_1059_315# _1012_/a_891_413# 0.31086f
C40927 _1012_/a_193_47# _1012_/a_975_413# 0
C40928 _1012_/a_466_413# _1012_/a_381_47# 0.03733f
C40929 _1039_/a_634_159# _0176_ 0.02157f
C40930 clknet_1_0__leaf__0459_ control0.add 0
C40931 _0528_/a_81_21# net11 0.00212f
C40932 _0148_ _0527_/a_109_297# 0.01113f
C40933 hold55/a_391_47# _1033_/a_27_47# 0
C40934 hold23/a_285_47# _0186_ 0
C40935 _0327_ net57 0
C40936 _0846_/a_51_297# _0345_ 0.11384f
C40937 net36 hold25/a_285_47# 0.00925f
C40938 hold79/a_391_47# _0484_ 0
C40939 net226 _0970_/a_27_297# 0
C40940 hold79/a_285_47# _0485_ 0
C40941 _0216_ _1031_/a_975_413# 0
C40942 _0107_ _1009_/a_891_413# 0
C40943 net46 _0610_/a_59_75# 0.1726f
C40944 _0179_ clknet_1_1__leaf__0465_ 1.23421f
C40945 comp0.B\[8\] _1046_/a_891_413# 0.00107f
C40946 _1002_/a_193_47# hold93/a_391_47# 0
C40947 _0749_/a_81_21# _0462_ 0.00464f
C40948 hold86/a_285_47# hold86/a_391_47# 0.41909f
C40949 _0662_/a_81_21# _0991_/a_891_413# 0
C40950 _0268_ net47 0
C40951 _1050_/a_27_47# acc0.A\[4\] 0.05751f
C40952 hold67/a_285_47# VPWR 0.28954f
C40953 _0452_ acc0.A\[15\] 0
C40954 _0343_ clkload3/Y 0.00241f
C40955 _0343_ _1030_/a_466_413# 0
C40956 _1055_/a_193_47# acc0.A\[9\] 0
C40957 _0990_/a_975_413# _0181_ 0.0011f
C40958 hold47/a_49_47# net132 0
C40959 net36 _0081_ 0
C40960 _0326_ _0460_ 0.03729f
C40961 _1041_/a_1059_315# _0546_/a_240_47# 0
C40962 _1041_/a_891_413# _0546_/a_149_47# 0
C40963 _0766_/a_109_297# _0462_ 0
C40964 _0485_ net17 0
C40965 _0958_/a_197_47# _0477_ 0
C40966 _0350_ _0988_/a_193_47# 0.00134f
C40967 A[3] net10 0.01933f
C40968 hold26/a_391_47# net173 0.13057f
C40969 acc0.A\[5\] hold7/a_285_47# 0
C40970 _0259_ net76 0
C40971 _0565_/a_149_47# net201 0.01613f
C40972 _0458_ hold28/a_391_47# 0
C40973 _0730_/a_510_47# _0350_ 0.00105f
C40974 comp0.B\[7\] comp0.B\[6\] 0.003f
C40975 hold74/a_391_47# VPWR 0.17276f
C40976 hold96/a_49_47# output52/a_27_47# 0
C40977 _0586_/a_27_47# _0352_ 0.04333f
C40978 clknet_1_0__leaf__0460_ _0247_ 0
C40979 _0544_/a_149_47# _1043_/a_193_47# 0
C40980 _0369_ _0830_/a_510_47# 0.00103f
C40981 _0813_/a_109_297# _0288_ 0
C40982 _0646_/a_47_47# _0797_/a_207_413# 0
C40983 net84 net43 0.12431f
C40984 hold16/a_49_47# acc0.A\[30\] 0.0013f
C40985 _0129_ _0704_/a_150_297# 0
C40986 comp0.B\[13\] hold37/a_49_47# 0
C40987 _0230_ net51 0.15686f
C40988 net169 _1052_/a_27_47# 0
C40989 net140 _1052_/a_193_47# 0
C40990 net120 _0175_ 0
C40991 _0513_/a_81_21# clknet_1_1__leaf__0465_ 0.03422f
C40992 _0457_ net105 0.00203f
C40993 _0409_ _0300_ 0.49403f
C40994 hold24/a_49_47# net36 0.04213f
C40995 _0176_ _1040_/a_1017_47# 0.00191f
C40996 _0311_ clkbuf_0__0461_/a_110_47# 0
C40997 net21 _1044_/a_561_413# 0
C40998 _0504_/a_27_47# _0181_ 0
C40999 _0463_ _0953_/a_32_297# 0.00185f
C41000 _0956_/a_32_297# _0173_ 0
C41001 _0718_/a_47_47# _0128_ 0
C41002 clknet_1_0__leaf__0458_ _0629_/a_145_75# 0
C41003 _0241_ net206 0
C41004 net64 _0988_/a_27_47# 0.02619f
C41005 net45 _1018_/a_1059_315# 0.01202f
C41006 _0995_/a_381_47# _0797_/a_207_413# 0
C41007 net59 _0219_ 0.0399f
C41008 _0108_ hold95/a_49_47# 0
C41009 _1031_/a_1059_315# _0339_ 0.00373f
C41010 _1031_/a_891_413# _0338_ 0
C41011 net205 _1036_/a_975_413# 0
C41012 _0256_ net62 0.2119f
C41013 _0625_/a_59_75# clkbuf_1_0__f__0465_/a_110_47# 0.01355f
C41014 net193 _1046_/a_891_413# 0
C41015 _0144_ _0177_ 0
C41016 net8 _0465_ 0.00247f
C41017 _0456_ _0181_ 0.02304f
C41018 net72 _0350_ 0
C41019 comp0.B\[1\] _0213_ 0
C41020 _0251_ _0432_ 0.00111f
C41021 _1054_/a_381_47# net75 0
C41022 _0432_ _0640_/a_109_53# 0.01556f
C41023 _0443_ _0640_/a_297_297# 0.00214f
C41024 _1001_/a_193_47# _0350_ 0
C41025 _1012_/a_381_47# net98 0
C41026 _0518_/a_27_297# acc0.A\[4\] 0
C41027 pp[30] _0712_/a_561_47# 0
C41028 _1046_/a_634_159# _1046_/a_381_47# 0
C41029 _0475_ _0956_/a_304_297# 0
C41030 A[12] acc0.A\[10\] 0
C41031 _0991_/a_634_159# _0263_ 0
C41032 net233 hold100/a_285_47# 0
C41033 net40 net5 0.08339f
C41034 net123 control0.sh 0.01645f
C41035 acc0.A\[21\] _0373_ 0.00285f
C41036 _0481_ _0484_ 0.00606f
C41037 _0557_/a_51_297# _0549_/a_68_297# 0
C41038 pp[26] _0570_/a_109_297# 0
C41039 net54 _0570_/a_373_47# 0
C41040 _1032_/a_381_47# clknet_1_0__leaf__0457_ 0.00101f
C41041 net140 net12 0.22539f
C41042 _0174_ _1045_/a_891_413# 0.00107f
C41043 net166 _0582_/a_373_47# 0
C41044 _1016_/a_381_47# _0115_ 0.01975f
C41045 _0119_ _0165_ 0
C41046 control0.state\[1\] VPWR 3.31106f
C41047 _0221_ _0707_/a_315_47# 0.00416f
C41048 _0403_ _0654_/a_207_413# 0
C41049 VPWR _0698_/a_199_47# 0
C41050 hold68/a_285_47# _0122_ 0.00271f
C41051 hold68/a_391_47# net110 0.01793f
C41052 _0753_/a_297_297# _0225_ 0.00698f
C41053 _0180_ hold7/a_49_47# 0
C41054 _1051_/a_193_47# _1050_/a_634_159# 0
C41055 _1051_/a_634_159# _1050_/a_193_47# 0
C41056 _1051_/a_27_47# _1050_/a_466_413# 0.00126f
C41057 _1051_/a_466_413# _1050_/a_27_47# 0.00126f
C41058 _1039_/a_27_47# clkbuf_1_0__f__0463_/a_110_47# 0.00567f
C41059 _0623_/a_109_297# net63 0.00122f
C41060 VPWR _0583_/a_109_47# 0
C41061 _0957_/a_32_297# _0496_/a_27_47# 0.00184f
C41062 _0284_ _0422_ 0
C41063 _0404_ _0993_/a_27_47# 0
C41064 _0458_ _0218_ 0.0025f
C41065 _0985_/a_634_159# net175 0
C41066 clknet_1_0__leaf__0462_ hold53/a_49_47# 0
C41067 VPWR net19 0.40963f
C41068 _1050_/a_891_413# _1045_/a_27_47# 0
C41069 _0634_/a_113_47# _0264_ 0
C41070 hold58/a_285_47# net26 0.00237f
C41071 hold9/a_49_47# _1028_/a_27_47# 0.03548f
C41072 _0208_ clkbuf_0__0457_/a_110_47# 0
C41073 _0984_/a_891_413# _0346_ 0
C41074 _0559_/a_51_297# clknet_0__0463_ 0.01739f
C41075 _0996_/a_561_413# acc0.A\[15\] 0
C41076 clknet_1_0__leaf__0463_ _1038_/a_891_413# 0
C41077 _0785_/a_299_297# _0181_ 0.0056f
C41078 net196 _0542_/a_149_47# 0
C41079 hold33/a_391_47# _0172_ 0.04207f
C41080 _0531_/a_27_297# _1049_/a_891_413# 0
C41081 pp[28] _0728_/a_145_75# 0
C41082 hold34/a_49_47# input16/a_75_212# 0.06919f
C41083 pp[2] output61/a_27_47# 0.08165f
C41084 output58/a_27_47# pp[3] 0
C41085 _0998_/a_466_413# clknet_1_1__leaf__0461_ 0.00241f
C41086 _0662_/a_384_47# _0401_ 0
C41087 _0661_/a_27_297# _0426_ 0
C41088 _0554_/a_68_297# comp0.B\[6\] 0
C41089 _0775_/a_79_21# _0347_ 0.14299f
C41090 _0457_ _1032_/a_1059_315# 0.04527f
C41091 _0130_ net17 0.01925f
C41092 net58 _0432_ 0.00486f
C41093 net44 _0999_/a_561_413# 0
C41094 hold76/a_285_47# _0616_/a_78_199# 0
C41095 pp[30] hold16/a_391_47# 0.00769f
C41096 _0290_ clknet_1_1__leaf__0458_ 0
C41097 _1016_/a_466_413# _0218_ 0
C41098 VPWR _0610_/a_145_75# 0
C41099 VPWR _0999_/a_466_413# 0.26934f
C41100 clkload3/Y _0998_/a_193_47# 0
C41101 _1052_/a_634_159# acc0.A\[6\] 0.04235f
C41102 acc0.A\[12\] _0399_ 0.02649f
C41103 _0581_/a_27_297# _0581_/a_373_47# 0.01338f
C41104 _0229_ _0227_ 0.1933f
C41105 net55 _0690_/a_68_297# 0
C41106 _0179_ _0522_/a_109_297# 0
C41107 clknet_1_1__leaf__0459_ _0187_ 0
C41108 net10 net154 0
C41109 _0311_ hold69/a_49_47# 0.00297f
C41110 VPWR _0691_/a_150_297# 0.00213f
C41111 acc0.A\[22\] net50 0.3056f
C41112 _1039_/a_381_47# net8 0.0126f
C41113 net188 VPWR 0.13999f
C41114 _0985_/a_381_47# _0083_ 0.1291f
C41115 _0287_ hold82/a_49_47# 0
C41116 _0325_ net93 0
C41117 hold85/a_391_47# _0476_ 0.04124f
C41118 _0343_ _0990_/a_466_413# 0.00819f
C41119 _0985_/a_27_47# acc0.A\[3\] 0.1493f
C41120 _0967_/a_215_297# _0970_/a_27_297# 0
C41121 _0404_ _0409_ 0.52393f
C41122 output58/a_27_47# _0273_ 0
C41123 clknet_1_1__leaf__0459_ clknet_1_1__leaf__0461_ 0.64991f
C41124 _1053_/a_193_47# _0191_ 0
C41125 hold101/a_49_47# _0346_ 0.059f
C41126 _0982_/a_193_47# _0080_ 0.17469f
C41127 _0982_/a_891_413# _0982_/a_1017_47# 0.00617f
C41128 _0982_/a_634_159# net68 0
C41129 control0.reset _0560_/a_68_297# 0
C41130 _0343_ net104 0
C41131 _1049_/a_27_47# _0147_ 0.09543f
C41132 _1049_/a_193_47# net135 0.01355f
C41133 _1049_/a_1059_315# _1049_/a_1017_47# 0
C41134 _0653_/a_113_47# net38 0
C41135 _0795_/a_81_21# _0669_/a_29_53# 0
C41136 clknet_1_0__leaf__0462_ _0227_ 0
C41137 clknet_0__0465_ _0186_ 0
C41138 _0483_ _0486_ 0
C41139 input6/a_75_212# A[14] 0.19704f
C41140 _0985_/a_193_47# _0504_/a_27_47# 0
C41141 _0606_/a_215_297# _0606_/a_109_53# 0.08065f
C41142 _1070_/a_27_47# _1070_/a_466_413# 0.27314f
C41143 _1070_/a_193_47# _1070_/a_634_159# 0.12729f
C41144 _0399_ _0445_ 0.10945f
C41145 _1052_/a_1059_315# _0523_/a_81_21# 0.00146f
C41146 _1053_/a_193_47# _1053_/a_381_47# 0.10164f
C41147 _1053_/a_634_159# _1053_/a_891_413# 0.03684f
C41148 _1053_/a_27_47# _1053_/a_561_413# 0.0027f
C41149 output44/a_27_47# _1030_/a_193_47# 0
C41150 _0381_ _0460_ 0.00287f
C41151 _1057_/a_193_47# acc0.A\[10\] 0.03363f
C41152 _0578_/a_27_297# net23 0
C41153 clknet_1_0__leaf__0465_ _1050_/a_193_47# 0.00345f
C41154 _0714_/a_240_47# _0218_ 0.05008f
C41155 hold54/a_285_47# clknet_1_0__leaf__0461_ 0.02913f
C41156 _0156_ net37 0.02249f
C41157 net45 _0998_/a_27_47# 0.00998f
C41158 _0996_/a_466_413# _0181_ 0
C41159 _0236_ net51 0
C41160 _1066_/a_193_47# clknet_1_1__leaf_clk 0.0042f
C41161 _1066_/a_1059_315# _1066_/a_1017_47# 0
C41162 net56 net96 0
C41163 clkload2/Y net154 0.00221f
C41164 acc0.A\[2\] net10 0
C41165 pp[10] net3 0.06826f
C41166 _0255_ net148 0.00616f
C41167 _0314_ _1007_/a_193_47# 0.00153f
C41168 _0313_ _1007_/a_27_47# 0
C41169 _0327_ _1010_/a_1059_315# 0
C41170 _1037_/a_634_159# _0176_ 0
C41171 net222 _0261_ 0
C41172 _1034_/a_466_413# _0175_ 0
C41173 pp[9] _0189_ 0
C41174 net31 _1040_/a_891_413# 0
C41175 _0201_ _1042_/a_891_413# 0
C41176 net177 _1022_/a_193_47# 0
C41177 net109 _1022_/a_634_159# 0.0237f
C41178 _1068_/a_27_47# _0166_ 0.13691f
C41179 _1068_/a_1059_315# _1068_/a_1017_47# 0
C41180 net206 _0450_ 0
C41181 _1030_/a_1059_315# _1030_/a_891_413# 0.31086f
C41182 _1030_/a_193_47# _1030_/a_975_413# 0
C41183 _1030_/a_466_413# _1030_/a_381_47# 0.03733f
C41184 clkbuf_1_1__f__0464_/a_110_47# _1044_/a_634_159# 0.01343f
C41185 _1041_/a_891_413# _0176_ 0
C41186 _0712_/a_561_47# _0339_ 0.00173f
C41187 hold5/a_49_47# net127 0
C41188 _0217_ net215 0.22296f
C41189 _0134_ net161 0
C41190 net71 _0448_ 0.00203f
C41191 _0627_/a_215_53# _0255_ 0.12102f
C41192 clkbuf_1_1__f__0465_/a_110_47# _0817_/a_266_47# 0
C41193 net32 net174 0
C41194 hold74/a_391_47# clknet_1_0__leaf__0459_ 0
C41195 hold5/a_285_47# _0543_/a_68_297# 0
C41196 _0995_/a_27_47# net42 0.01089f
C41197 clkbuf_1_1__f__0464_/a_110_47# net184 0.00179f
C41198 net81 _0219_ 0.01484f
C41199 _0461_ _0616_/a_493_297# 0
C41200 net188 input4/a_75_212# 0
C41201 _0312_ _1009_/a_592_47# 0
C41202 VPWR _0570_/a_109_47# 0
C41203 _0571_/a_109_297# net113 0
C41204 _1035_/a_592_47# clknet_1_1__leaf__0463_ 0
C41205 _0601_/a_68_297# _0366_ 0
C41206 _0992_/a_891_413# net37 0.01039f
C41207 _0346_ hold91/a_391_47# 0.0068f
C41208 control0.count\[1\] _0486_ 0
C41209 hold18/a_285_47# _0346_ 0
C41210 clknet_1_1__leaf__0463_ B[15] 0.00902f
C41211 _0251_ pp[7] 0.00124f
C41212 _0598_/a_79_21# _0230_ 0.10671f
C41213 _0598_/a_382_297# _0226_ 0
C41214 VPWR _0517_/a_384_47# 0
C41215 _1015_/a_561_413# _0181_ 0
C41216 _0320_ _0737_/a_285_47# 0
C41217 _0987_/a_193_47# _0987_/a_891_413# 0.19489f
C41218 _0987_/a_27_47# _0987_/a_381_47# 0.06222f
C41219 _0987_/a_634_159# _0987_/a_1059_315# 0
C41220 _0632_/a_113_47# clknet_1_0__leaf__0461_ 0
C41221 _0151_ net15 0
C41222 _0337_ acc0.A\[29\] 0
C41223 _0238_ _0294_ 0.10479f
C41224 _0182_ _0261_ 0
C41225 acc0.A\[1\] _0263_ 0
C41226 net194 _1051_/a_634_159# 0
C41227 _0579_/a_27_297# _0183_ 0.22138f
C41228 _0579_/a_109_47# _0217_ 0.00307f
C41229 clkbuf_1_0__f__0461_/a_110_47# net47 0
C41230 _0695_/a_80_21# _0367_ 0
C41231 _0262_ net218 0
C41232 hold49/a_391_47# _1044_/a_27_47# 0
C41233 _0134_ net26 0.01024f
C41234 acc0.A\[1\] _1047_/a_27_47# 0.00118f
C41235 _1052_/a_193_47# input14/a_75_212# 0
C41236 _0314_ _0328_ 0.00195f
C41237 clknet_0__0459_ hold82/a_285_47# 0
C41238 acc0.A\[20\] _0765_/a_79_21# 0.05433f
C41239 net184 _0186_ 0
C41240 acc0.A\[27\] _1008_/a_1017_47# 0
C41241 hold43/a_391_47# acc0.A\[27\] 0
C41242 _1000_/a_561_413# VPWR 0.00308f
C41243 clknet_1_0__leaf__0465_ _0518_/a_109_297# 0
C41244 _1004_/a_193_47# _1004_/a_634_159# 0.11072f
C41245 _1004_/a_27_47# _1004_/a_466_413# 0.27314f
C41246 VPWR _0155_ 0.20627f
C41247 _0216_ acc0.A\[23\] 0.2102f
C41248 clkbuf_1_0__f__0459_/a_110_47# _0114_ 0.01271f
C41249 hold16/a_391_47# _0339_ 0.02956f
C41250 _0169_ _0466_ 0.12701f
C41251 _0983_/a_1017_47# _0181_ 0
C41252 _0557_/a_51_297# _1035_/a_27_47# 0
C41253 _1072_/a_592_47# _0466_ 0
C41254 _0151_ _1053_/a_1059_315# 0
C41255 pp[27] hold61/a_391_47# 0.00561f
C41256 _0476_ _0958_/a_109_47# 0
C41257 _0403_ _0286_ 0
C41258 _0534_/a_81_21# _0145_ 0.11436f
C41259 _0176_ net147 0
C41260 net9 hold83/a_391_47# 0
C41261 _0154_ acc0.A\[10\] 0.0011f
C41262 _0379_ net50 0.12425f
C41263 _1029_/a_634_159# _1029_/a_1059_315# 0
C41264 _1029_/a_27_47# _1029_/a_381_47# 0.06222f
C41265 _1029_/a_193_47# _1029_/a_891_413# 0.19685f
C41266 VPWR hold50/a_391_47# 0.20093f
C41267 _0479_ _0478_ 0.34934f
C41268 hold21/a_391_47# _0186_ 0
C41269 net211 _0580_/a_27_297# 0
C41270 pp[7] net58 0
C41271 _0856_/a_215_47# _0346_ 0.0548f
C41272 _0218_ pp[14] 0
C41273 hold67/a_285_47# hold35/a_391_47# 0
C41274 VPWR _0565_/a_245_297# 0.00619f
C41275 clkbuf_0__0464_/a_110_47# _0148_ 0
C41276 _0999_/a_1059_315# _0407_ 0
C41277 _0318_ _0321_ 0.09723f
C41278 _0502_/a_27_47# net134 0
C41279 input14/a_75_212# net12 0.03784f
C41280 _0805_/a_27_47# _0091_ 0
C41281 net61 _0271_ 0.2822f
C41282 _0637_/a_139_47# _0450_ 0
C41283 _0343_ _0998_/a_592_47# 0
C41284 net219 _0393_ 0.04396f
C41285 _0275_ acc0.A\[6\] 0
C41286 _0401_ net47 0
C41287 _0346_ _0670_/a_510_47# 0
C41288 _0430_ _0831_/a_285_47# 0.00127f
C41289 clkload0/a_27_47# _1072_/a_466_413# 0.00168f
C41290 hold65/a_391_47# VPWR 0.1661f
C41291 comp0.B\[13\] _1045_/a_891_413# 0.03821f
C41292 _0172_ _0194_ 0
C41293 hold66/a_285_47# _0754_/a_240_47# 0
C41294 acc0.A\[4\] _0987_/a_27_47# 0.03386f
C41295 acc0.A\[12\] _0295_ 0
C41296 _1015_/a_27_47# _0565_/a_240_47# 0
C41297 _1015_/a_1059_315# _0565_/a_51_297# 0.00944f
C41298 _0476_ _0160_ 0.04452f
C41299 hold97/a_391_47# _0345_ 0.1257f
C41300 _0182_ _0509_/a_27_47# 0.17238f
C41301 _0661_/a_27_297# _0289_ 0.20238f
C41302 net168 _0180_ 0.67772f
C41303 _0581_/a_27_297# _0347_ 0
C41304 _0121_ net51 0
C41305 _0998_/a_975_413# acc0.A\[17\] 0
C41306 A[10] _0514_/a_109_297# 0
C41307 acc0.A\[14\] _0347_ 0.0228f
C41308 acc0.A\[27\] _0729_/a_68_297# 0
C41309 net222 net47 0
C41310 _1037_/a_381_47# clknet_1_1__leaf__0463_ 0
C41311 _0998_/a_381_47# clkbuf_1_1__f__0461_/a_110_47# 0
C41312 _1033_/a_1059_315# _0956_/a_32_297# 0
C41313 _0960_/a_109_47# _0976_/a_505_21# 0
C41314 _1028_/a_634_159# _1028_/a_466_413# 0.23992f
C41315 _1028_/a_193_47# _1028_/a_1059_315# 0.03405f
C41316 _1028_/a_27_47# _1028_/a_891_413# 0.03071f
C41317 hold41/a_285_47# hold42/a_285_47# 0.00672f
C41318 acc0.A\[1\] clknet_1_0__leaf__0461_ 0.00111f
C41319 A[12] _0188_ 0.02225f
C41320 _0629_/a_59_75# _0856_/a_215_47# 0
C41321 net216 _0324_ 0
C41322 _0371_ _0359_ 0
C41323 _0369_ _0989_/a_193_47# 0.00577f
C41324 _0399_ net42 0.04919f
C41325 _0837_/a_81_21# _0255_ 0
C41326 _0440_ _0835_/a_78_199# 0
C41327 net58 _0986_/a_381_47# 0.00823f
C41328 _0195_ hold60/a_391_47# 0.02926f
C41329 _0216_ hold60/a_49_47# 0
C41330 net194 clknet_1_0__leaf__0465_ 0.02893f
C41331 _0306_ _1009_/a_891_413# 0
C41332 _1033_/a_381_47# _0131_ 0.12138f
C41333 _1033_/a_466_413# comp0.B\[1\] 0
C41334 _0369_ _0992_/a_193_47# 0.00338f
C41335 _0467_ clknet_0_clk 0.24484f
C41336 _0985_/a_891_413# VPWR 0.1894f
C41337 net63 _0987_/a_561_413# 0
C41338 _0554_/a_68_297# net26 0.00561f
C41339 net125 _0176_ 0.09306f
C41340 VPWR _1018_/a_1059_315# 0.39244f
C41341 net186 comp0.B\[4\] 0
C41342 clknet_1_1__leaf__0460_ _0354_ 0
C41343 clknet_0__0463_ net180 0.00106f
C41344 _0521_/a_299_297# clknet_1_0__leaf__0465_ 0.00597f
C41345 _0197_ acc0.A\[3\] 0.12406f
C41346 VPWR _1049_/a_634_159# 0.18357f
C41347 hold55/a_285_47# _0130_ 0.00324f
C41348 _0647_/a_129_47# clknet_1_1__leaf__0459_ 0.00289f
C41349 hold67/a_285_47# net182 0
C41350 _0123_ _0347_ 0
C41351 _0743_/a_512_297# _0367_ 0
C41352 _0743_/a_149_47# _0315_ 0
C41353 VPWR _0552_/a_150_297# 0.00142f
C41354 acc0.A\[21\] _0761_/a_113_47# 0
C41355 net88 hold93/a_285_47# 0.0103f
C41356 _1041_/a_27_47# net31 0.05467f
C41357 net207 net149 0
C41358 _1009_/a_1017_47# _0219_ 0.0023f
C41359 _0375_ net46 0.45166f
C41360 VPWR _1066_/a_634_159# 0.19448f
C41361 _0538_/a_51_297# clknet_1_1__leaf__0464_ 0
C41362 _0833_/a_215_47# clkbuf_1_1__f__0458_/a_110_47# 0
C41363 _0704_/a_68_297# clknet_1_1__leaf__0462_ 0
C41364 VPWR _1068_/a_634_159# 0.18202f
C41365 pp[28] hold61/a_285_47# 0
C41366 pp[27] clknet_1_1__leaf__0462_ 0
C41367 net49 _0487_ 0
C41368 _0962_/a_109_297# _0480_ 0.0156f
C41369 clknet_1_1__leaf__0459_ _0671_/a_199_47# 0
C41370 net44 clkbuf_1_1__f__0461_/a_110_47# 0
C41371 clknet_0_clk comp0.B\[0\] 0.20469f
C41372 _0741_/a_109_297# _0219_ 0
C41373 _0315_ _0345_ 0.39364f
C41374 _0258_ hold101/a_285_47# 0
C41375 _0626_/a_150_297# net248 0
C41376 _0277_ acc0.A\[15\] 0.04152f
C41377 _0993_/a_27_47# _0419_ 0
C41378 _0993_/a_634_159# _0417_ 0
C41379 _0993_/a_381_47# net79 0
C41380 clknet_0__0457_ hold60/a_285_47# 0.00489f
C41381 net231 comp0.B\[3\] 0
C41382 hold66/a_391_47# _0228_ 0.01283f
C41383 clknet_1_0__leaf__0464_ _0528_/a_384_47# 0
C41384 clknet_1_0__leaf__0465_ _1046_/a_634_159# 0.00216f
C41385 _0107_ _0680_/a_217_297# 0
C41386 clknet_1_1__leaf__0460_ _0693_/a_68_297# 0.00127f
C41387 _0642_/a_215_297# acc0.A\[8\] 0.0849f
C41388 _0697_/a_217_297# _0689_/a_68_297# 0
C41389 _0343_ _0983_/a_891_413# 0.02425f
C41390 _0531_/a_109_297# net175 0.00248f
C41391 net167 _1071_/a_1059_315# 0
C41392 _0170_ _1071_/a_193_47# 0
C41393 _0996_/a_27_47# acc0.A\[13\] 0
C41394 _0174_ _0463_ 0.03776f
C41395 _0699_/a_68_297# _0319_ 0
C41396 acc0.A\[0\] hold2/a_391_47# 0.00285f
C41397 hold19/a_391_47# hold72/a_285_47# 0
C41398 acc0.A\[14\] _1016_/a_891_413# 0
C41399 _1002_/a_381_47# acc0.A\[20\] 0
C41400 _0998_/a_466_413# _0998_/a_561_413# 0.00772f
C41401 _0998_/a_634_159# _0998_/a_975_413# 0
C41402 _1019_/a_193_47# clkbuf_0__0457_/a_110_47# 0.02269f
C41403 pp[17] net60 0.01057f
C41404 _0579_/a_109_297# hold40/a_49_47# 0
C41405 _0579_/a_27_297# hold40/a_285_47# 0.00193f
C41406 _0216_ hold61/a_391_47# 0
C41407 _1009_/a_27_47# _0318_ 0
C41408 _0305_ _0673_/a_253_47# 0.00158f
C41409 _0552_/a_68_297# _0550_/a_51_297# 0
C41410 acc0.A\[11\] _0806_/a_113_297# 0
C41411 _0118_ _0369_ 0
C41412 _0529_/a_109_47# _0186_ 0.00214f
C41413 _0498_/a_245_297# _0465_ 0
C41414 _0779_/a_510_47# _0308_ 0
C41415 hold10/a_285_47# net247 0
C41416 _1003_/a_381_47# _0369_ 0
C41417 net238 _0400_ 0
C41418 _0410_ _0405_ 0.05764f
C41419 _0118_ clknet_0__0457_ 0.17868f
C41420 net110 _1023_/a_891_413# 0
C41421 _0122_ _1023_/a_1059_315# 0
C41422 _1024_/a_193_47# acc0.A\[23\] 0
C41423 _0259_ _0986_/a_193_47# 0
C41424 _0388_ clknet_1_0__leaf__0461_ 0
C41425 clkbuf_1_1__f__0463_/a_110_47# comp0.B\[5\] 0
C41426 _0362_ _0370_ 0.00159f
C41427 _0310_ _0394_ 0.09519f
C41428 hold38/a_285_47# comp0.B\[3\] 0.08312f
C41429 _0496_/a_27_47# _0213_ 0.01599f
C41430 _0191_ acc0.A\[4\] 0
C41431 _0717_/a_303_47# _0221_ 0
C41432 _1019_/a_634_159# _1019_/a_381_47# 0
C41433 _1046_/a_381_47# net132 0
C41434 net77 _0263_ 0
C41435 _1057_/a_193_47# _0188_ 0
C41436 clknet_0__0464_ net10 0.39938f
C41437 clknet_1_0__leaf__0464_ _0180_ 0.46337f
C41438 net133 acc0.A\[1\] 0.0106f
C41439 _0342_ net116 0
C41440 net61 pp[2] 0.00776f
C41441 net72 _0986_/a_634_159# 0
C41442 VPWR _1012_/a_891_413# 0.19934f
C41443 clknet_1_0__leaf__0464_ net218 0
C41444 _0218_ _0408_ 0
C41445 _1004_/a_193_47# net46 0
C41446 _0565_/a_240_47# _0215_ 0
C41447 _0635_/a_27_47# _0264_ 0.03892f
C41448 _0469_ _1063_/a_27_47# 0.00119f
C41449 hold83/a_285_47# _0522_/a_27_297# 0.00108f
C41450 _0473_ _0176_ 0.18717f
C41451 _0343_ pp[18] 0
C41452 _0726_/a_51_297# _0726_/a_245_297# 0.01218f
C41453 _1050_/a_466_413# net131 0
C41454 _1050_/a_634_159# net184 0
C41455 clkbuf_1_0__f__0463_/a_110_47# _0953_/a_32_297# 0
C41456 net108 net49 0.00426f
C41457 _1058_/a_193_47# net67 0.02899f
C41458 _0580_/a_373_47# _0345_ 0
C41459 _0994_/a_1059_315# output40/a_27_47# 0
C41460 net9 _1049_/a_561_413# 0
C41461 net175 _1049_/a_1017_47# 0
C41462 _0243_ _0343_ 0
C41463 hold8/a_391_47# acc0.A\[25\] 0
C41464 _0786_/a_80_21# hold70/a_391_47# 0.00271f
C41465 _0293_ _0426_ 0.00531f
C41466 hold25/a_285_47# _1039_/a_27_47# 0
C41467 net53 net50 0
C41468 pp[27] net242 0
C41469 _0334_ net116 0
C41470 _0291_ _0218_ 0
C41471 _0393_ _0352_ 0.09752f
C41472 net1 _0566_/a_27_47# 0
C41473 acc0.A\[31\] _1031_/a_891_413# 0.00277f
C41474 acc0.A\[1\] _0585_/a_27_297# 0
C41475 _0533_/a_27_297# net149 0
C41476 net162 _1031_/a_466_413# 0
C41477 _0902_/a_27_47# _0610_/a_59_75# 0
C41478 _0342_ hold92/a_285_47# 0
C41479 VPWR _0998_/a_27_47# 0.46026f
C41480 _0982_/a_466_413# net207 0
C41481 hold3/a_49_47# hold3/a_285_47# 0.22264f
C41482 clkbuf_1_1__f__0464_/a_110_47# _0176_ 0
C41483 hold23/a_49_47# _0270_ 0
C41484 _0335_ hold61/a_49_47# 0
C41485 clknet_1_0__leaf__0465_ _0987_/a_193_47# 0.01323f
C41486 net45 net46 0.0135f
C41487 _1021_/a_1059_315# _0578_/a_109_297# 0
C41488 _1021_/a_891_413# _0578_/a_27_297# 0
C41489 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# 1.6339f
C41490 net166 _0218_ 0
C41491 net81 _0799_/a_209_297# 0.00178f
C41492 _0758_/a_79_21# _0352_ 0.21125f
C41493 _1024_/a_891_413# pp[24] 0
C41494 _1024_/a_561_413# net52 0
C41495 _0294_ _0991_/a_466_413# 0
C41496 _0991_/a_634_159# _0218_ 0
C41497 _0380_ net51 0.00116f
C41498 clkload2/Y clknet_0__0464_ 0.00131f
C41499 _0581_/a_373_47# _0116_ 0
C41500 _0990_/a_1059_315# _0990_/a_891_413# 0.31086f
C41501 _0990_/a_193_47# _0990_/a_975_413# 0
C41502 _0990_/a_466_413# _0990_/a_381_47# 0.03733f
C41503 _0463_ _0208_ 0
C41504 net219 net206 0
C41505 net69 net165 0.15805f
C41506 clknet_0__0458_ clkload1/Y 0.00105f
C41507 _0461_ _0771_/a_27_413# 0.00138f
C41508 _0790_/a_35_297# _0219_ 0.06451f
C41509 _1002_/a_466_413# clknet_1_0__leaf__0457_ 0.00117f
C41510 _1002_/a_193_47# _0460_ 0.04524f
C41511 _0322_ clkbuf_1_1__f__0460_/a_110_47# 0.00245f
C41512 _0369_ net142 0
C41513 net64 _0642_/a_215_297# 0
C41514 _0571_/a_109_297# hold8/a_285_47# 0.00197f
C41515 _0571_/a_27_297# hold8/a_391_47# 0
C41516 clkbuf_1_1__f__0465_/a_110_47# _0181_ 0.04721f
C41517 _0984_/a_1017_47# net58 0
C41518 _0327_ clkbuf_1_1__f__0460_/a_110_47# 0.17009f
C41519 clknet_0__0465_ net62 0.21321f
C41520 _0172_ net195 0.00839f
C41521 hold86/a_285_47# _0268_ 0
C41522 net203 _0132_ 0
C41523 _0343_ _0088_ 0.02604f
C41524 _0967_/a_215_297# _0967_/a_487_297# 0.00167f
C41525 hold49/a_49_47# _0176_ 0.00501f
C41526 _0346_ _1014_/a_1017_47# 0
C41527 _0260_ _0626_/a_68_297# 0
C41528 _0343_ _0407_ 0.03383f
C41529 comp0.B\[10\] _0205_ 0.04061f
C41530 hold24/a_49_47# _1039_/a_27_47# 0
C41531 hold53/a_285_47# _1025_/a_1059_315# 0.00108f
C41532 hold53/a_49_47# _1025_/a_891_413# 0.00386f
C41533 _0123_ _1025_/a_27_47# 0
C41534 hold53/a_391_47# _1025_/a_466_413# 0.00388f
C41535 _1049_/a_975_413# acc0.A\[3\] 0
C41536 _0195_ net113 0.18078f
C41537 _0216_ clknet_1_1__leaf__0462_ 0.57796f
C41538 _1034_/a_1059_315# _0955_/a_32_297# 0
C41539 hold52/a_391_47# _0366_ 0
C41540 clknet_1_0__leaf__0459_ _1018_/a_1059_315# 0
C41541 control0.add _0345_ 0.13133f
C41542 _0230_ hold3/a_391_47# 0
C41543 net216 _0104_ 0.00719f
C41544 net243 _0576_/a_373_47# 0
C41545 _0606_/a_297_297# _0236_ 0.00392f
C41546 _0606_/a_215_297# _0238_ 0.1016f
C41547 _0850_/a_68_297# _0264_ 0.02652f
C41548 _0229_ _0352_ 0
C41549 _0469_ _1062_/a_1059_315# 0
C41550 _1070_/a_27_47# _0168_ 0.07442f
C41551 _1070_/a_634_159# VPWR 0.21773f
C41552 _1070_/a_1059_315# _1070_/a_1017_47# 0
C41553 net106 _1033_/a_27_47# 0
C41554 _1045_/a_27_47# _1045_/a_1059_315# 0.04875f
C41555 _1045_/a_193_47# _1045_/a_466_413# 0.08301f
C41556 net44 _1030_/a_592_47# 0
C41557 acc0.A\[12\] _0515_/a_299_297# 0
C41558 net61 clknet_1_0__leaf__0465_ 0.0371f
C41559 _0209_ control0.sh 0.00401f
C41560 _0146_ _0465_ 0.00473f
C41561 _0689_/a_150_297# _0345_ 0
C41562 clknet_1_0__leaf__0462_ hold30/a_49_47# 0.01673f
C41563 comp0.B\[11\] _0541_/a_68_297# 0.17714f
C41564 clknet_0__0459_ _0671_/a_113_297# 0
C41565 _0179_ _0150_ 0.15657f
C41566 _1014_/a_891_413# _0465_ 0
C41567 _1062_/a_891_413# _0468_ 0
C41568 VPWR _1030_/a_891_413# 0.1788f
C41569 _0089_ net47 0.00655f
C41570 _1043_/a_27_47# _1043_/a_1059_315# 0.04875f
C41571 _1043_/a_193_47# _1043_/a_466_413# 0.07482f
C41572 net7 _1040_/a_891_413# 0
C41573 _0465_ _0492_/a_27_47# 0.00441f
C41574 _0183_ net36 0.02087f
C41575 acc0.A\[2\] _0146_ 0
C41576 net21 net128 0
C41577 _0749_/a_299_297# _0219_ 0
C41578 clkbuf_1_1__f__0464_/a_110_47# net130 0.07977f
C41579 _0315_ net52 0.30068f
C41580 _1038_/a_466_413# _0209_ 0
C41581 hold63/a_285_47# net200 0
C41582 _0678_/a_150_297# _0219_ 0
C41583 hold52/a_49_47# _0217_ 0
C41584 _0763_/a_109_47# _0460_ 0
C41585 _1004_/a_634_159# VPWR 0.18379f
C41586 _1021_/a_1059_315# _1002_/a_27_47# 0.011f
C41587 _1021_/a_634_159# _1002_/a_634_159# 0
C41588 _1021_/a_466_413# _1002_/a_193_47# 0
C41589 _1021_/a_193_47# _1002_/a_466_413# 0.00811f
C41590 hold89/a_49_47# _0484_ 0
C41591 _0767_/a_59_75# _0359_ 0
C41592 clkbuf_1_1__f_clk/a_110_47# _0564_/a_68_297# 0
C41593 clknet_1_0__leaf__0462_ _0352_ 0.03297f
C41594 clknet_1_0__leaf__0458_ _1047_/a_1059_315# 0.00546f
C41595 _0785_/a_299_297# _0990_/a_193_47# 0
C41596 acc0.A\[12\] _0091_ 0
C41597 hold65/a_49_47# acc0.A\[6\] 0.0318f
C41598 _1056_/a_1059_315# _1056_/a_891_413# 0.31086f
C41599 _1056_/a_466_413# _1056_/a_381_47# 0.03733f
C41600 _0182_ _0173_ 0
C41601 _1032_/a_975_413# net17 0.00103f
C41602 hold28/a_49_47# _0180_ 0
C41603 hold28/a_285_47# _0182_ 0
C41604 comp0.B\[10\] _1042_/a_193_47# 0
C41605 acc0.A\[4\] clkbuf_1_0__f__0465_/a_110_47# 0
C41606 _0294_ _0401_ 0.16488f
C41607 _0290_ _0218_ 0
C41608 _0271_ _0431_ 0.47782f
C41609 pp[27] _0730_/a_297_297# 0
C41610 hold28/a_49_47# net218 0
C41611 _0987_/a_466_413# _0085_ 0.0306f
C41612 _0987_/a_1059_315# net73 0
C41613 net194 _1044_/a_466_413# 0
C41614 _0704_/a_68_297# hold92/a_49_47# 0.01017f
C41615 net130 _0186_ 0.00331f
C41616 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# 1.65433f
C41617 net194 net137 0.0019f
C41618 _0464_ _0181_ 0
C41619 _0367_ clknet_1_0__leaf__0460_ 0.00146f
C41620 _0655_/a_109_93# _0671_/a_113_297# 0
C41621 _0245_ _0773_/a_117_297# 0.0018f
C41622 _1007_/a_193_47# _0360_ 0
C41623 _0855_/a_299_297# _0456_ 0.00207f
C41624 net185 clknet_1_1__leaf__0463_ 0.00617f
C41625 _0199_ _1047_/a_381_47# 0.00149f
C41626 _0239_ _0394_ 0
C41627 _0145_ hold71/a_391_47# 0
C41628 _1041_/a_1059_315# _0548_/a_51_297# 0.00126f
C41629 _1041_/a_27_47# _0548_/a_240_47# 0
C41630 VPWR hold81/a_49_47# 0.28578f
C41631 _1004_/a_1059_315# _1004_/a_1017_47# 0
C41632 _0216_ net242 0
C41633 net47 _0986_/a_891_413# 0
C41634 output57/a_27_47# hold80/a_49_47# 0.02157f
C41635 net162 _0712_/a_465_47# 0
C41636 _1059_/a_27_47# _0158_ 0
C41637 net145 _1060_/a_193_47# 0
C41638 _0983_/a_27_47# _0983_/a_634_159# 0.13601f
C41639 _0667_/a_113_47# pp[15] 0
C41640 _0854_/a_79_21# _0459_ 0
C41641 clknet_1_0__leaf__0465_ _1045_/a_27_47# 0.00817f
C41642 net36 acc0.A\[15\] 0.14834f
C41643 hold69/a_285_47# clknet_0__0460_ 0
C41644 clknet_1_1__leaf__0464_ net11 0
C41645 _1029_/a_466_413# net191 0
C41646 _1019_/a_891_413# _0352_ 0
C41647 output46/a_27_47# pp[19] 0.15855f
C41648 net24 B[5] 0.00152f
C41649 B[1] net28 0.09556f
C41650 clknet_1_0__leaf__0458_ _0186_ 0.00348f
C41651 _0334_ hold80/a_285_47# 0
C41652 _0257_ _0825_/a_68_297# 0
C41653 output59/a_27_47# net116 0.07335f
C41654 _0217_ clknet_1_0__leaf__0460_ 0.19327f
C41655 comp0.B\[13\] _1044_/a_1059_315# 0
C41656 _0328_ _0360_ 0.29467f
C41657 clknet_1_0__leaf__0462_ _0574_/a_109_297# 0.00675f
C41658 _0497_/a_68_297# _0176_ 0.10193f
C41659 _0462_ _0242_ 0.00905f
C41660 acc0.A\[1\] _0218_ 0
C41661 _0718_/a_285_47# _0221_ 0
C41662 _0747_/a_79_21# _0350_ 0.00174f
C41663 net213 _0377_ 0
C41664 clknet_1_0__leaf__0459_ _0998_/a_27_47# 0.00983f
C41665 hold47/a_391_47# _0180_ 0.00372f
C41666 _1000_/a_1059_315# acc0.A\[18\] 0
C41667 net117 _0218_ 0
C41668 _1020_/a_381_47# _0217_ 0
C41669 _0650_/a_68_297# _0091_ 0
C41670 _1020_/a_1059_315# _0183_ 0
C41671 _0279_ net80 0.01615f
C41672 acc0.A\[29\] _0333_ 0.15563f
C41673 _0806_/a_113_297# _0281_ 0.06591f
C41674 net103 _1016_/a_592_47# 0
C41675 _0289_ _0293_ 0.00117f
C41676 _0116_ _0347_ 0.20078f
C41677 net206 _0352_ 0.00221f
C41678 net162 hold16/a_285_47# 0.01397f
C41679 pp[8] acc0.A\[9\] 0.04312f
C41680 _0854_/a_297_297# clknet_1_0__leaf__0461_ 0
C41681 _1016_/a_193_47# _1016_/a_381_47# 0.09503f
C41682 _1016_/a_634_159# _1016_/a_891_413# 0.03684f
C41683 _1016_/a_27_47# _1016_/a_561_413# 0.00163f
C41684 hold13/a_285_47# _0176_ 0
C41685 net60 _0567_/a_109_297# 0
C41686 VPWR _0726_/a_245_297# 0.00619f
C41687 _0724_/a_113_297# net116 0
C41688 output37/a_27_47# net37 0.22061f
C41689 clknet_1_1__leaf__0459_ clknet_1_1__leaf__0465_ 0.00536f
C41690 hold11/a_49_47# _1061_/a_891_413# 0
C41691 hold11/a_391_47# _1061_/a_466_413# 0
C41692 output59/a_27_47# hold92/a_285_47# 0
C41693 _0613_/a_109_297# _0393_ 0
C41694 _0960_/a_181_47# _0488_ 0.00172f
C41695 _1028_/a_466_413# net114 0.00146f
C41696 hold25/a_391_47# _1041_/a_634_159# 0
C41697 hold25/a_285_47# _1041_/a_466_413# 0
C41698 net9 input9/a_27_47# 0.11083f
C41699 net49 _0760_/a_47_47# 0
C41700 hold41/a_391_47# net189 0.00331f
C41701 _0095_ clknet_1_1__leaf__0461_ 0
C41702 hold17/a_391_47# _1070_/a_193_47# 0
C41703 hold31/a_49_47# _0252_ 0.04982f
C41704 _0343_ _0996_/a_592_47# 0
C41705 hold42/a_285_47# net4 0
C41706 _1067_/a_1059_315# control0.reset 0
C41707 _1057_/a_634_159# _0187_ 0.02087f
C41708 _1057_/a_1059_315# net4 0
C41709 _0812_/a_79_21# _0422_ 0.13238f
C41710 _0385_ clknet_1_0__leaf__0457_ 0.00148f
C41711 VPWR _0990_/a_891_413# 0.19127f
C41712 _0542_/a_51_297# hold51/a_391_47# 0
C41713 _0999_/a_1059_315# _0096_ 0
C41714 _0131_ comp0.B\[1\] 0
C41715 hold57/a_391_47# _0207_ 0
C41716 clknet_0__0462_ _0737_/a_35_297# 0.02853f
C41717 VPWR _0564_/a_68_297# 0.15513f
C41718 _0655_/a_215_53# clkbuf_1_1__f__0459_/a_110_47# 0
C41719 _0110_ net239 0
C41720 acc0.A\[16\] hold19/a_49_47# 0.05387f
C41721 _0557_/a_240_47# _1037_/a_1059_315# 0
C41722 _0557_/a_149_47# _1037_/a_891_413# 0
C41723 VPWR net135 0.4839f
C41724 _0584_/a_27_297# _0584_/a_373_47# 0.01338f
C41725 _1059_/a_27_47# acc0.A\[14\] 0.06668f
C41726 net219 _0774_/a_150_297# 0
C41727 _0475_ _0560_/a_68_297# 0
C41728 _1041_/a_27_47# net7 0.4793f
C41729 hold59/a_285_47# _0181_ 0
C41730 _0211_ input24/a_75_212# 0.00219f
C41731 _0238_ _0371_ 0
C41732 _0179_ net36 0
C41733 hold4/a_49_47# _1022_/a_193_47# 0
C41734 hold4/a_285_47# _1022_/a_27_47# 0.00329f
C41735 net238 clkbuf_0__0459_/a_110_47# 0
C41736 _1017_/a_1059_315# clknet_0__0461_ 0.01005f
C41737 _0460_ _1006_/a_975_413# 0
C41738 _0742_/a_81_21# net52 0.01204f
C41739 _0186_ _0525_/a_299_297# 0
C41740 _0764_/a_81_21# _0346_ 0.19366f
C41741 VPWR clknet_1_1__leaf_clk 2.69097f
C41742 _0532_/a_81_21# _1047_/a_891_413# 0
C41743 _0532_/a_299_297# _1047_/a_1059_315# 0
C41744 _0198_ _1047_/a_27_47# 0
C41745 net53 _0743_/a_245_297# 0
C41746 net63 acc0.A\[8\] 0.02195f
C41747 _0170_ _1072_/a_466_413# 0.00139f
C41748 _0370_ _0324_ 0
C41749 A[11] _0512_/a_27_297# 0.0339f
C41750 hold27/a_49_47# hold27/a_285_47# 0.22264f
C41751 pp[9] net67 0.14832f
C41752 _0562_/a_150_297# _0173_ 0
C41753 output65/a_27_47# output61/a_27_47# 0.0033f
C41754 net81 _0997_/a_891_413# 0
C41755 _0343_ net208 0.0261f
C41756 _0241_ _1006_/a_27_47# 0
C41757 _1054_/a_27_47# VPWR 0.64122f
C41758 _0643_/a_103_199# _0626_/a_68_297# 0.01178f
C41759 pp[27] hold80/a_49_47# 0
C41760 _0305_ _0776_/a_27_47# 0.00125f
C41761 _0149_ _0987_/a_27_47# 0
C41762 net137 _0987_/a_193_47# 0
C41763 _1051_/a_27_47# _0085_ 0
C41764 _1051_/a_193_47# net73 0
C41765 clknet_1_0__leaf__0462_ _1025_/a_466_413# 0.00856f
C41766 _0536_/a_51_297# net10 0
C41767 _1056_/a_891_413# VPWR 0.18554f
C41768 _0993_/a_592_47# _0091_ 0
C41769 _0215_ _0171_ 0
C41770 _0770_/a_79_21# _0389_ 0.09514f
C41771 _0216_ hold92/a_49_47# 0.05973f
C41772 net122 B[4] 0.0055f
C41773 net234 VPWR 0.68946f
C41774 _0292_ clknet_1_1__leaf__0465_ 0.09371f
C41775 _0388_ _0218_ 0
C41776 pp[26] VPWR 0.26221f
C41777 _0742_/a_299_297# clknet_1_0__leaf__0460_ 0
C41778 _1018_/a_193_47# acc0.A\[18\] 0.04947f
C41779 clknet_1_0__leaf__0465_ net132 0.02166f
C41780 acc0.A\[22\] _0576_/a_27_297# 0
C41781 _0217_ _0576_/a_109_297# 0.07433f
C41782 _1028_/a_193_47# _0106_ 0
C41783 hold57/a_391_47# _1039_/a_1059_315# 0
C41784 hold57/a_285_47# _1039_/a_891_413# 0.00101f
C41785 _0996_/a_381_47# _0185_ 0
C41786 _0305_ _0219_ 0.08347f
C41787 clknet_0_clk _1068_/a_381_47# 0.00162f
C41788 _0349_ _0219_ 0.01746f
C41789 net1 clknet_0_clk 0.03303f
C41790 hold56/a_49_47# _0956_/a_32_297# 0
C41791 _0227_ _0382_ 0
C41792 net46 VPWR 1.9931f
C41793 _0342_ _0220_ 0.1116f
C41794 hold1/a_49_47# net148 0
C41795 acc0.A\[12\] net192 0.00356f
C41796 _0416_ net80 0
C41797 _1021_/a_193_47# _0385_ 0
C41798 net178 _1055_/a_891_413# 0
C41799 _0479_ VPWR 0.45124f
C41800 hold30/a_49_47# hold30/a_391_47# 0.00188f
C41801 _0159_ _1061_/a_891_413# 0
C41802 net203 _1033_/a_592_47# 0
C41803 hold56/a_391_47# _0131_ 0
C41804 net224 net95 0
C41805 _0369_ _0988_/a_27_47# 0.00441f
C41806 _0248_ clknet_1_0__leaf__0460_ 0.20586f
C41807 _0984_/a_592_47# net47 0
C41808 _1001_/a_193_47# _0195_ 0
C41809 _1019_/a_193_47# _0350_ 0
C41810 acc0.A\[12\] _0346_ 0.06737f
C41811 _1019_/a_891_413# net207 0
C41812 _1019_/a_381_47# net105 0.00764f
C41813 net35 _1071_/a_193_47# 0.00224f
C41814 _0965_/a_47_47# _0483_ 0.14429f
C41815 _0539_/a_68_297# comp0.B\[12\] 0.17842f
C41816 net51 _1005_/a_891_413# 0.0094f
C41817 _0220_ _0334_ 0.00494f
C41818 _0195_ hold8/a_285_47# 0.00919f
C41819 net155 hold8/a_49_47# 0
C41820 _0271_ _0269_ 0
C41821 _0357_ acc0.A\[27\] 0
C41822 _0172_ _0204_ 0
C41823 _0174_ clkbuf_1_0__f__0463_/a_110_47# 0.27179f
C41824 VPWR _0584_/a_109_47# 0
C41825 _0381_ _0373_ 0.05157f
C41826 net43 _0776_/a_109_297# 0
C41827 hold52/a_391_47# acc0.A\[24\] 0.06411f
C41828 hold83/a_285_47# _0193_ 0
C41829 _0343_ _0995_/a_193_47# 0.03886f
C41830 _1014_/a_634_159# clknet_1_0__leaf__0461_ 0.01316f
C41831 _0575_/a_27_297# net50 0.00527f
C41832 _0726_/a_512_297# net227 0.0018f
C41833 _0726_/a_240_47# _0354_ 0.0148f
C41834 _0726_/a_149_47# _0355_ 0.00984f
C41835 _0673_/a_103_199# acc0.A\[13\] 0
C41836 clkbuf_1_0__f__0461_/a_110_47# _0581_/a_109_297# 0
C41837 _0458_ _0268_ 0.10157f
C41838 _0172_ hold6/a_391_47# 0.02824f
C41839 _0858_/a_27_47# hold71/a_49_47# 0.00862f
C41840 _0393_ hold72/a_285_47# 0
C41841 comp0.B\[14\] net32 0
C41842 _0716_/a_27_47# _0404_ 0
C41843 net242 _1010_/a_561_413# 0
C41844 _0287_ _0655_/a_297_297# 0
C41845 _0800_/a_51_297# clknet_1_1__leaf__0459_ 0.01833f
C41846 net45 _0783_/a_297_297# 0
C41847 net207 net206 0
C41848 control0.state\[0\] _1064_/a_1059_315# 0.00115f
C41849 net34 _1064_/a_634_159# 0.01607f
C41850 control0.state\[1\] _1064_/a_466_413# 0
C41851 _0274_ _0826_/a_27_53# 0.01572f
C41852 _0275_ _0826_/a_219_297# 0
C41853 _0272_ _0826_/a_301_297# 0
C41854 _1033_/a_634_159# clknet_1_1__leaf__0463_ 0
C41855 _1015_/a_891_413# _0584_/a_27_297# 0
C41856 hold86/a_285_47# net222 0
C41857 _1050_/a_193_47# _0148_ 0.25826f
C41858 _0283_ hold81/a_49_47# 0.01188f
C41859 hold46/a_49_47# net10 0.01794f
C41860 _1020_/a_27_47# _0181_ 0
C41861 _1001_/a_466_413# _0247_ 0
C41862 _0951_/a_209_311# hold84/a_391_47# 0.01572f
C41863 net245 _0800_/a_240_47# 0.1103f
C41864 _0199_ net149 0.1177f
C41865 _0200_ _0176_ 0.02862f
C41866 acc0.A\[1\] _0112_ 0
C41867 _0179_ _0515_/a_81_21# 0.00373f
C41868 _0080_ net207 0.00192f
C41869 clknet_0__0457_ _1001_/a_27_47# 0.05233f
C41870 clkbuf_1_0__f__0457_/a_110_47# _1001_/a_466_413# 0
C41871 net46 net48 0
C41872 _1020_/a_1059_315# hold40/a_285_47# 0.0054f
C41873 _0467_ _1065_/a_27_47# 0.44676f
C41874 _0216_ _1047_/a_27_47# 0
C41875 _0346_ _0445_ 0
C41876 _0465_ _1048_/a_381_47# 0
C41877 clknet_1_0__leaf__0465_ _0431_ 0.00582f
C41878 _0402_ net67 0
C41879 _0965_/a_47_47# control0.count\[1\] 0
C41880 hold59/a_49_47# _1018_/a_193_47# 0.00209f
C41881 hold59/a_285_47# _1018_/a_27_47# 0.00178f
C41882 _0838_/a_109_297# _0255_ 0.00304f
C41883 hold100/a_285_47# _0264_ 0
C41884 _0294_ _0089_ 0.02697f
C41885 net77 _0218_ 0.15579f
C41886 _0495_/a_68_297# _0173_ 0.0047f
C41887 _0176_ comp0.B\[8\] 0.78494f
C41888 _0990_/a_381_47# _0088_ 0.13417f
C41889 A[6] net13 0.00473f
C41890 comp0.B\[3\] _1066_/a_634_159# 0
C41891 comp0.B\[5\] _1066_/a_27_47# 0
C41892 _0982_/a_634_159# _0264_ 0
C41893 _0610_/a_145_75# _0345_ 0
C41894 _0100_ clknet_1_0__leaf__0457_ 0.00232f
C41895 _0999_/a_466_413# _0345_ 0
C41896 acc0.A\[2\] _1048_/a_381_47# 0
C41897 _0793_/a_51_297# _0407_ 0.14843f
C41898 _0807_/a_68_297# net246 0.10273f
C41899 hold83/a_49_47# _0150_ 0
C41900 acc0.A\[16\] _1017_/a_193_47# 0.03828f
C41901 _0482_ hold89/a_285_47# 0
C41902 _0461_ _0580_/a_27_297# 0
C41903 _0229_ _0237_ 0.11127f
C41904 _0331_ hold50/a_49_47# 0
C41905 _0228_ _0374_ 0
C41906 hold56/a_49_47# hold56/a_285_47# 0.22264f
C41907 _0313_ _0740_/a_113_47# 0
C41908 hold86/a_285_47# _0182_ 0
C41909 hold86/a_391_47# acc0.A\[1\] 0
C41910 _0539_/a_150_297# _0202_ 0
C41911 VPWR _0996_/a_27_47# 0.70574f
C41912 _0958_/a_303_47# _0468_ 0.00259f
C41913 acc0.A\[11\] A[9] 0
C41914 _0390_ net46 0.28234f
C41915 net66 _0512_/a_27_297# 0
C41916 _0995_/a_27_47# net60 0
C41917 _1065_/a_27_47# comp0.B\[0\] 0.0067f
C41918 comp0.B\[7\] _1039_/a_381_47# 0
C41919 _0856_/a_79_21# _0850_/a_68_297# 0.01992f
C41920 net200 _1025_/a_592_47# 0.00105f
C41921 _1051_/a_27_47# _1044_/a_193_47# 0
C41922 _1051_/a_193_47# _1044_/a_27_47# 0
C41923 _0995_/a_27_47# net5 0
C41924 clknet_1_1__leaf__0460_ hold77/a_49_47# 0.01856f
C41925 _1037_/a_634_159# net28 0.00321f
C41926 _1034_/a_1059_315# _0474_ 0.01764f
C41927 _0777_/a_285_47# clknet_1_1__leaf__0461_ 0.00562f
C41928 _1051_/a_634_159# _1051_/a_592_47# 0
C41929 _1045_/a_193_47# _1044_/a_634_159# 0
C41930 _1045_/a_466_413# _1044_/a_27_47# 0
C41931 _1045_/a_27_47# _1044_/a_466_413# 0.01155f
C41932 _1045_/a_634_159# _1044_/a_193_47# 0
C41933 comp0.B\[14\] _1042_/a_1059_315# 0
C41934 clkbuf_1_0__f__0463_/a_110_47# _0208_ 0
C41935 hold15/a_391_47# hold61/a_391_47# 0
C41936 _0227_ _1005_/a_634_159# 0
C41937 _0576_/a_27_297# _0379_ 0
C41938 acc0.A\[21\] _1005_/a_466_413# 0
C41939 net58 _0841_/a_215_47# 0.01246f
C41940 _1051_/a_27_47# net131 0
C41941 _0656_/a_59_75# _0218_ 0.00119f
C41942 _0294_ _0656_/a_145_75# 0
C41943 net62 _0986_/a_27_47# 0.04321f
C41944 _0501_/a_27_47# _0499_/a_59_75# 0.00235f
C41945 _1045_/a_891_413# _1045_/a_1017_47# 0.00617f
C41946 _1045_/a_193_47# net184 0.2311f
C41947 _1045_/a_634_159# net131 0
C41948 hold56/a_49_47# _1032_/a_193_47# 0
C41949 hold56/a_285_47# _1032_/a_27_47# 0
C41950 net23 _1067_/a_634_159# 0.03749f
C41951 _0680_/a_217_297# _0346_ 0
C41952 _0305_ _0746_/a_81_21# 0.00101f
C41953 _1003_/a_193_47# net213 0
C41954 net157 _0566_/a_27_47# 0.025f
C41955 clknet_1_0__leaf__0462_ _0237_ 0.00261f
C41956 _1072_/a_27_47# clknet_1_0__leaf_clk 0.23118f
C41957 VPWR _1043_/a_975_413# 0.00484f
C41958 _0309_ _0394_ 0.42315f
C41959 _0618_/a_297_297# _0219_ 0.0011f
C41960 hold63/a_285_47# hold63/a_391_47# 0.41909f
C41961 _0837_/a_81_21# hold1/a_49_47# 0
C41962 clknet_1_0__leaf__0458_ hold100/a_49_47# 0.00447f
C41963 _0096_ _0397_ 0
C41964 _0733_/a_79_199# _0322_ 0.00209f
C41965 _1043_/a_891_413# _1043_/a_1017_47# 0.00617f
C41966 _1043_/a_193_47# net196 0.2026f
C41967 _1043_/a_634_159# net129 0
C41968 _1018_/a_381_47# _0399_ 0
C41969 hold32/a_49_47# net16 0.13034f
C41970 VPWR _1015_/a_1059_315# 0.40171f
C41971 comp0.B\[14\] net10 0.27865f
C41972 net193 _0176_ 0.00559f
C41973 net133 _0198_ 0.00127f
C41974 _0314_ _0123_ 0
C41975 net103 hold72/a_391_47# 0.00373f
C41976 _1003_/a_27_47# _0947_/a_109_297# 0
C41977 _0467_ hold12/a_285_47# 0.00175f
C41978 clknet_1_0__leaf__0458_ _0982_/a_193_47# 0
C41979 _0181_ _0776_/a_27_47# 0.0011f
C41980 _0216_ clknet_1_0__leaf__0461_ 0.72693f
C41981 clknet_1_1__leaf__0460_ _0743_/a_51_297# 0
C41982 _0459_ _0240_ 0
C41983 _1034_/a_193_47# _1065_/a_193_47# 0
C41984 _0210_ input24/a_75_212# 0
C41985 _0734_/a_285_47# acc0.A\[27\] 0.02153f
C41986 _0343_ _0096_ 0.00186f
C41987 net120 comp0.B\[4\] 0.00168f
C41988 _1042_/a_634_159# net153 0
C41989 net172 _0209_ 0
C41990 _0369_ _0459_ 0.07561f
C41991 _0104_ _0370_ 0
C41992 VPWR _0630_/a_109_297# 0.00429f
C41993 VPWR _0654_/a_207_413# 0.16491f
C41994 clknet_0__0457_ _0459_ 0.00578f
C41995 clknet_1_1__leaf__0458_ _0825_/a_68_297# 0.01513f
C41996 _1021_/a_634_159# net88 0.00827f
C41997 _1021_/a_193_47# _0100_ 0
C41998 _0119_ _1002_/a_193_47# 0.00102f
C41999 _1032_/a_27_47# _1032_/a_193_47# 0.97453f
C42000 _1054_/a_466_413# _1054_/a_561_413# 0.00772f
C42001 _1054_/a_634_159# _1054_/a_975_413# 0
C42002 _0393_ _0392_ 0.10968f
C42003 _1071_/a_891_413# control0.count\[0\] 0
C42004 _1015_/a_193_47# _1015_/a_381_47# 0.09503f
C42005 _1015_/a_634_159# _1015_/a_891_413# 0.03684f
C42006 _1015_/a_27_47# _1015_/a_561_413# 0.0027f
C42007 comp0.B\[7\] net174 0
C42008 _0983_/a_561_413# VPWR 0.00248f
C42009 _0180_ clkbuf_1_0__f__0464_/a_110_47# 0.07785f
C42010 _0174_ _1042_/a_1017_47# 0.00133f
C42011 _0557_/a_51_297# _0173_ 0.14207f
C42012 _0991_/a_193_47# _0347_ 0
C42013 _0357_ _1010_/a_193_47# 0
C42014 _0399_ acc0.A\[17\] 0.00269f
C42015 _0358_ _1010_/a_27_47# 0
C42016 _0181_ _0219_ 0.46807f
C42017 clkbuf_1_0__f__0464_/a_110_47# net218 0
C42018 _0751_/a_29_53# _0227_ 0.13961f
C42019 net247 _0263_ 0.06429f
C42020 net113 _1027_/a_466_413# 0
C42021 clknet_1_1__leaf__0462_ _1027_/a_891_413# 0.0081f
C42022 _0352_ _0773_/a_35_297# 0.03521f
C42023 net46 clknet_1_0__leaf__0459_ 0
C42024 _0343_ _1031_/a_193_47# 0.01912f
C42025 _0752_/a_300_297# _0228_ 0
C42026 _0234_ _0605_/a_109_297# 0
C42027 _0792_/a_80_21# _0408_ 0.08836f
C42028 _0792_/a_303_47# _0400_ 0.00214f
C42029 VPWR _0550_/a_51_297# 0.48486f
C42030 net247 _1047_/a_27_47# 0
C42031 net53 _0322_ 0
C42032 _0319_ _0686_/a_219_297# 0
C42033 _1038_/a_634_159# _1038_/a_381_47# 0
C42034 _1053_/a_634_159# _0180_ 0
C42035 _0829_/a_27_47# _0435_ 0.105f
C42036 net10 _0543_/a_68_297# 0
C42037 _0082_ _0451_ 0
C42038 _0654_/a_27_413# _0654_/a_207_413# 0.18542f
C42039 _0319_ _1008_/a_1059_315# 0.00151f
C42040 _1067_/a_27_47# clknet_1_0__leaf__0461_ 0.01849f
C42041 net53 _0327_ 0
C42042 _0745_/a_109_47# _0370_ 0.01083f
C42043 net45 _0777_/a_47_47# 0
C42044 output59/a_27_47# _0220_ 0
C42045 pp[30] _0705_/a_59_75# 0.00191f
C42046 clknet_1_0__leaf__0458_ net62 0
C42047 _0446_ _0845_/a_109_47# 0.06155f
C42048 net194 _0148_ 0
C42049 clknet_1_0__leaf__0458_ _0450_ 0.05702f
C42050 net61 _0529_/a_373_47# 0
C42051 net181 acc0.A\[10\] 0
C42052 _0983_/a_381_47# _0983_/a_561_413# 0.00123f
C42053 _0983_/a_27_47# net69 0.23268f
C42054 _0983_/a_891_413# _0983_/a_975_413# 0.00851f
C42055 net214 hold67/a_391_47# 0.132f
C42056 clknet_1_0__leaf__0465_ _1051_/a_592_47# 0
C42057 acc0.A\[21\] net187 0
C42058 hold59/a_391_47# _0242_ 0
C42059 _0995_/a_1059_315# input6/a_75_212# 0
C42060 _0347_ _0380_ 0.00105f
C42061 _0261_ _0844_/a_297_47# 0.05603f
C42062 net40 _0995_/a_891_413# 0.0345f
C42063 net245 _0995_/a_466_413# 0.01639f
C42064 net234 _0453_ 0.04002f
C42065 _0456_ _0452_ 0
C42066 _0346_ net42 0.02332f
C42067 _0290_ net228 0
C42068 clknet_1_0__leaf__0460_ _0755_/a_109_297# 0
C42069 hold89/a_49_47# hold89/a_391_47# 0.00188f
C42070 _0245_ _1006_/a_193_47# 0
C42071 _0985_/a_381_47# net71 0
C42072 _0399_ net5 0.9248f
C42073 _0172_ _0493_/a_27_47# 0
C42074 net21 comp0.B\[11\] 0.00367f
C42075 net183 comp0.B\[12\] 0.00366f
C42076 _0343_ _0093_ 0.02689f
C42077 hold50/a_391_47# _0345_ 0
C42078 _0747_/a_215_47# _1006_/a_27_47# 0
C42079 _0747_/a_79_21# _1006_/a_634_159# 0
C42080 _0087_ pp[5] 0
C42081 _0592_/a_150_297# net51 0
C42082 _0588_/a_113_47# acc0.A\[30\] 0
C42083 _0466_ _1068_/a_1059_315# 0.02725f
C42084 net90 _1007_/a_891_413# 0
C42085 _0318_ _0685_/a_68_297# 0
C42086 _1048_/a_27_47# _1047_/a_466_413# 0
C42087 _1048_/a_193_47# _1047_/a_634_159# 0
C42088 _1048_/a_466_413# _1047_/a_27_47# 0
C42089 _0767_/a_59_75# _0767_/a_145_75# 0.00658f
C42090 _1003_/a_592_47# _0217_ 0
C42091 _1004_/a_1059_315# net50 0.1086f
C42092 _0852_/a_117_297# _0265_ 0.0014f
C42093 _0852_/a_285_47# net47 0.00254f
C42094 clknet_1_0__leaf__0462_ _1005_/a_27_47# 0.00203f
C42095 _1061_/a_27_47# acc0.A\[15\] 0
C42096 hold87/a_285_47# net206 0
C42097 clknet_0__0459_ _0996_/a_381_47# 0.00106f
C42098 _0616_/a_215_47# _0614_/a_29_53# 0
C42099 hold77/a_391_47# net95 0
C42100 net247 clknet_1_0__leaf__0461_ 0
C42101 _0361_ _0743_/a_240_47# 0
C42102 clknet_1_1__leaf__0462_ _1026_/a_975_413# 0
C42103 net113 _1026_/a_381_47# 0
C42104 _0195_ _0336_ 0.08744f
C42105 _0998_/a_193_47# _0096_ 0.44059f
C42106 _0998_/a_634_159# _0399_ 0.00152f
C42107 _0423_ _0347_ 0
C42108 net25 _0176_ 0
C42109 hold17/a_391_47# VPWR 0.17389f
C42110 _0263_ _0841_/a_79_21# 0
C42111 _0337_ hold61/a_391_47# 0.00154f
C42112 _0780_/a_35_297# _0308_ 0.20693f
C42113 _0555_/a_149_47# _0176_ 0
C42114 clknet_1_0__leaf__0459_ _0996_/a_27_47# 0
C42115 hold54/a_285_47# _0956_/a_32_297# 0
C42116 _0502_/a_27_47# _1049_/a_381_47# 0
C42117 _0131_ _0496_/a_27_47# 0.18286f
C42118 _0559_/a_512_297# VPWR 0.00642f
C42119 _0372_ _0346_ 0.02124f
C42120 _0397_ _0395_ 0.00651f
C42121 net39 _0994_/a_1017_47# 0.00168f
C42122 _1008_/a_27_47# hold50/a_49_47# 0.00317f
C42123 net61 output65/a_27_47# 0.02482f
C42124 _0216_ _0585_/a_27_297# 0.09879f
C42125 hold28/a_391_47# _0198_ 0
C42126 _0195_ _0585_/a_109_47# 0.00246f
C42127 _1014_/a_27_47# _0208_ 0
C42128 hold62/a_49_47# net209 0
C42129 _0985_/a_193_47# _0219_ 0
C42130 hold54/a_49_47# comp0.B\[1\] 0.31014f
C42131 net21 _0202_ 0.0411f
C42132 _0201_ net20 0.00357f
C42133 clknet_1_1__leaf__0459_ _1057_/a_381_47# 0
C42134 _0179_ _0527_/a_27_297# 0.01599f
C42135 _0255_ _0834_/a_109_297# 0.00113f
C42136 _1002_/a_891_413# acc0.A\[21\] 0
C42137 _1016_/a_27_47# clknet_0__0461_ 0
C42138 _1048_/a_1059_315# _0509_/a_27_47# 0
C42139 comp0.B\[4\] _1034_/a_466_413# 0
C42140 hold33/a_49_47# net174 0.11744f
C42141 _1056_/a_891_413# net182 0.00116f
C42142 clknet_1_1__leaf__0463_ _0487_ 0
C42143 hold29/a_391_47# net176 0.13055f
C42144 _1046_/a_1059_315# _0139_ 0
C42145 _1004_/a_466_413# net215 0
C42146 _0179_ _0989_/a_634_159# 0
C42147 _0179_ hold1/a_391_47# 0
C42148 _0717_/a_80_21# _0705_/a_59_75# 0
C42149 _0275_ _0626_/a_150_297# 0
C42150 clknet_1_1__leaf__0459_ _0398_ 0
C42151 acc0.A\[5\] _0987_/a_975_413# 0
C42152 VPWR _0569_/a_373_47# 0.00303f
C42153 hold39/a_49_47# _0475_ 0
C42154 _0343_ _0712_/a_297_297# 0.00825f
C42155 B[12] B[10] 0
C42156 clknet_1_0__leaf__0459_ _1015_/a_1059_315# 0
C42157 _0591_/a_109_297# _0352_ 0
C42158 _0174_ _0548_/a_245_297# 0
C42159 _1039_/a_27_47# acc0.A\[15\] 0
C42160 _0195_ _1050_/a_27_47# 0
C42161 _0163_ _1065_/a_381_47# 0.12573f
C42162 _0188_ _0511_/a_81_21# 0
C42163 VPWR _0783_/a_297_297# 0.00929f
C42164 _1038_/a_1017_47# VPWR 0
C42165 net11 net148 0.36577f
C42166 net154 net12 0
C42167 clknet_0__0458_ _0261_ 0
C42168 output64/a_27_47# _0621_/a_285_297# 0
C42169 comp0.B\[10\] clknet_1_1__leaf__0464_ 0.00127f
C42170 VPWR _0286_ 0.8042f
C42171 _0270_ net170 0
C42172 _0387_ _0352_ 0.00436f
C42173 _0257_ _0837_/a_81_21# 0
C42174 _0179_ _1061_/a_27_47# 0
C42175 _0989_/a_193_47# net75 0.00123f
C42176 clknet_0_clk control0.sh 0
C42177 net35 _1072_/a_466_413# 0.00197f
C42178 _1067_/a_381_47# clknet_1_0__leaf__0457_ 0.00504f
C42179 _1067_/a_1059_315# _0460_ 0.0014f
C42180 hold21/a_285_47# A[4] 0.00206f
C42181 _0485_ _0468_ 0
C42182 _0473_ _0954_/a_114_297# 0
C42183 _1059_/a_193_47# net41 0.00161f
C42184 _0241_ _0247_ 0.19601f
C42185 net233 _0264_ 0
C42186 _1020_/a_634_159# net118 0
C42187 _0757_/a_68_297# _0350_ 0.19062f
C42188 _0982_/a_193_47# hold18/a_49_47# 0
C42189 clkbuf_1_0__f__0457_/a_110_47# _0241_ 0
C42190 hold55/a_285_47# net187 0
C42191 net47 net229 0
C42192 _0286_ _0654_/a_27_413# 0
C42193 _0283_ _0654_/a_207_413# 0
C42194 clknet_1_1__leaf__0459_ _0277_ 0.06558f
C42195 _1053_/a_27_47# _0152_ 0
C42196 clkbuf_1_0__f__0463_/a_110_47# comp0.B\[9\] 0
C42197 _1031_/a_381_47# _1030_/a_193_47# 0
C42198 net133 net247 0.02343f
C42199 _0551_/a_27_47# comp0.B\[15\] 0.01618f
C42200 _0457_ _1067_/a_1059_315# 0.00131f
C42201 net205 _0561_/a_51_297# 0.00131f
C42202 VPWR _0794_/a_27_47# 0.01098f
C42203 _0176_ _1045_/a_193_47# 0
C42204 _1012_/a_381_47# _0395_ 0
C42205 _0299_ net5 0.09501f
C42206 _1032_/a_891_413# comp0.B\[15\] 0
C42207 net101 net1 0.19813f
C42208 hold7/a_391_47# net148 0.07662f
C42209 net160 _1037_/a_27_47# 0
C42210 _0712_/a_79_21# net60 0.00156f
C42211 net100 clknet_1_0__leaf__0461_ 0.21633f
C42212 _0458_ _0182_ 0.32599f
C42213 _0382_ _0352_ 0
C42214 _1025_/a_634_159# _1025_/a_381_47# 0
C42215 _0350_ hold95/a_285_47# 0
C42216 _0359_ _1006_/a_1059_315# 0
C42217 net227 _0109_ 0.06258f
C42218 hold64/a_49_47# _0459_ 0.01684f
C42219 _0218_ net83 0
C42220 _1012_/a_891_413# _0345_ 0
C42221 _1012_/a_193_47# _0219_ 0
C42222 net58 _0627_/a_297_297# 0
C42223 hold5/a_49_47# _1042_/a_27_47# 0.00142f
C42224 _0195_ _0208_ 0.47787f
C42225 net119 clknet_1_1__leaf__0463_ 0.23803f
C42226 B[11] _0541_/a_150_297# 0
C42227 _1055_/a_1059_315# _0181_ 0
C42228 _0113_ _0584_/a_109_47# 0
C42229 clkbuf_1_1__f__0463_/a_110_47# control0.reset 0
C42230 net238 hold91/a_391_47# 0.13545f
C42231 net205 _0133_ 0
C42232 _0410_ hold91/a_285_47# 0.0012f
C42233 _0168_ _0976_/a_218_374# 0
C42234 _1070_/a_1059_315# _0466_ 0
C42235 _1070_/a_891_413# _0488_ 0
C42236 VPWR _0976_/a_218_47# 0
C42237 _0800_/a_240_47# VPWR 0.00597f
C42238 _0781_/a_68_297# _0218_ 0.16568f
C42239 _0369_ _0772_/a_79_21# 0.10406f
C42240 _0157_ _0508_/a_299_297# 0.00558f
C42241 net145 _0508_/a_384_47# 0
C42242 hold54/a_391_47# _1032_/a_27_47# 0
C42243 hold54/a_285_47# _1032_/a_193_47# 0
C42244 VPWR _0913_/a_27_47# 0.19948f
C42245 hold49/a_285_47# _0954_/a_32_297# 0
C42246 _1046_/a_561_413# net10 0.00212f
C42247 comp0.B\[3\] _0564_/a_68_297# 0.01408f
C42248 clknet_1_1__leaf__0459_ _0808_/a_81_21# 0.011f
C42249 _0118_ hold40/a_391_47# 0.00832f
C42250 _0982_/a_634_159# _0856_/a_79_21# 0
C42251 _0982_/a_27_47# _0856_/a_215_47# 0
C42252 _0763_/a_109_47# _0373_ 0
C42253 hold17/a_285_47# hold17/a_391_47# 0.41909f
C42254 _0403_ _0994_/a_193_47# 0.00702f
C42255 net61 _0845_/a_109_47# 0.00395f
C42256 _0533_/a_27_297# comp0.B\[15\] 0.01329f
C42257 net31 net153 0.20609f
C42258 hold18/a_285_47# _0446_ 0.0035f
C42259 _1003_/a_891_413# control0.state\[2\] 0
C42260 hold58/a_49_47# _0212_ 0
C42261 _0996_/a_466_413# _0996_/a_561_413# 0.00772f
C42262 _0996_/a_634_159# _0996_/a_975_413# 0
C42263 _1055_/a_193_47# _0517_/a_299_297# 0.00165f
C42264 _1055_/a_634_159# _0517_/a_81_21# 0
C42265 _0458_ _0443_ 0
C42266 _0386_ _0347_ 0
C42267 _0291_ _0090_ 0
C42268 VPWR _0835_/a_215_47# 0.00335f
C42269 _1066_/a_27_47# hold84/a_49_47# 0.00693f
C42270 _0216_ _0105_ 0
C42271 _0753_/a_79_21# acc0.A\[23\] 0
C42272 hold64/a_285_47# clknet_1_0__leaf__0461_ 0.02035f
C42273 _0294_ _0679_/a_68_297# 0.07046f
C42274 comp0.B\[3\] clknet_1_1__leaf_clk 0
C42275 clknet_1_0__leaf__0464_ _1048_/a_891_413# 0
C42276 clknet_1_1__leaf__0457_ _1061_/a_466_413# 0.00395f
C42277 pp[19] net50 0
C42278 net46 pp[22] 0.00654f
C42279 _0234_ net241 0.01413f
C42280 _1060_/a_193_47# net6 0.00101f
C42281 _0732_/a_209_47# _0219_ 0.00139f
C42282 _0559_/a_51_297# _0559_/a_149_47# 0.02487f
C42283 _0211_ net121 0.00126f
C42284 hold57/a_285_47# _0475_ 0
C42285 _0317_ _0686_/a_27_53# 0.12798f
C42286 _0642_/a_215_297# _0369_ 0.00297f
C42287 _1057_/a_634_159# clknet_1_1__leaf__0465_ 0.03762f
C42288 clknet_0__0458_ net47 0
C42289 VPWR _1036_/a_193_47# 0.30962f
C42290 _0430_ clkbuf_1_1__f__0458_/a_110_47# 0.01744f
C42291 _0344_ _0999_/a_1059_315# 0
C42292 hold24/a_49_47# _0174_ 0.02292f
C42293 comp0.B\[7\] _0553_/a_149_47# 0
C42294 _0330_ _1008_/a_466_413# 0
C42295 _1044_/a_27_47# _1044_/a_634_159# 0.14145f
C42296 _0272_ _0640_/a_109_53# 0
C42297 _0274_ _0640_/a_215_297# 0.00978f
C42298 VPWR _0523_/a_299_297# 0.28272f
C42299 _0483_ clknet_0_clk 0.0073f
C42300 _0322_ clkbuf_1_1__f__0462_/a_110_47# 0
C42301 hold24/a_391_47# comp0.B\[10\] 0
C42302 comp0.B\[2\] comp0.B\[6\] 0.01963f
C42303 VPWR _0902_/a_27_47# 0.26779f
C42304 _1051_/a_891_413# acc0.A\[5\] 0.00338f
C42305 hold65/a_391_47# net212 0.13005f
C42306 hold65/a_285_47# _0437_ 0.0012f
C42307 hold64/a_49_47# _0265_ 0
C42308 net131 _1044_/a_193_47# 0
C42309 _1045_/a_193_47# net130 0
C42310 net184 _1044_/a_27_47# 0
C42311 clkbuf_1_1__f__0462_/a_110_47# _0327_ 0.00831f
C42312 A[10] acc0.A\[9\] 0.02833f
C42313 acc0.A\[21\] _0103_ 0
C42314 _0227_ net91 0.30317f
C42315 hold59/a_285_47# _0855_/a_299_297# 0
C42316 _0216_ _0218_ 0.13077f
C42317 _0337_ net242 0
C42318 _0369_ net51 0.00784f
C42319 _0992_/a_975_413# acc0.A\[10\] 0.00183f
C42320 _0440_ _0346_ 0.32872f
C42321 VPWR _0777_/a_47_47# 0.36294f
C42322 clknet_1_1__leaf__0461_ _0219_ 0.49026f
C42323 clknet_1_1__leaf__0459_ _0298_ 0.39736f
C42324 _0736_/a_139_47# VPWR 0
C42325 _0399_ _0990_/a_561_413# 0.00196f
C42326 net46 _1023_/a_27_47# 0.00447f
C42327 control0.state\[0\] hold93/a_285_47# 0
C42328 control0.state\[1\] hold93/a_49_47# 0.29968f
C42329 clknet_1_1__leaf__0458_ net148 0.23614f
C42330 _1011_/a_1059_315# _0723_/a_207_413# 0.00684f
C42331 _0789_/a_201_297# VPWR 0.20863f
C42332 _0440_ net65 0
C42333 hold100/a_391_47# _0449_ 0
C42334 _0274_ _0465_ 0.00949f
C42335 _1002_/a_975_413# net240 0
C42336 _1039_/a_634_159# clknet_0__0463_ 0.01164f
C42337 _0280_ net37 0
C42338 _0402_ _0302_ 0
C42339 _0714_/a_240_47# _1013_/a_27_47# 0
C42340 _0714_/a_149_47# _1013_/a_193_47# 0
C42341 _0271_ clkbuf_0__0458_/a_110_47# 0
C42342 clknet_1_1__leaf__0459_ _0296_ 0.00284f
C42343 clknet_1_1__leaf__0460_ _0308_ 0.003f
C42344 _1003_/a_381_47# _0467_ 0
C42345 input29/a_75_212# B[6] 0.19839f
C42346 VPWR _0673_/a_103_199# 0.45761f
C42347 acc0.A\[20\] _0183_ 0
C42348 net58 _0272_ 0
C42349 VPWR _0672_/a_79_21# 0.4772f
C42350 _0627_/a_215_53# clknet_1_1__leaf__0458_ 0.0019f
C42351 _0972_/a_250_297# _1062_/a_634_159# 0.00118f
C42352 _0972_/a_93_21# _1062_/a_466_413# 0
C42353 hold76/a_391_47# _1000_/a_193_47# 0
C42354 _0858_/a_27_47# _0532_/a_81_21# 0
C42355 _0849_/a_79_21# _0849_/a_215_47# 0.04584f
C42356 control0.count\[1\] clknet_0_clk 0
C42357 hold101/a_285_47# _0987_/a_27_47# 0
C42358 _1032_/a_466_413# _1032_/a_592_47# 0.00553f
C42359 _1032_/a_634_159# _1032_/a_1017_47# 0
C42360 _1054_/a_561_413# net169 0
C42361 _0568_/a_27_297# net208 0.13036f
C42362 output42/a_27_47# net40 0
C42363 pp[15] hold98/a_49_47# 0.01753f
C42364 _1015_/a_1059_315# _0113_ 0.01618f
C42365 clknet_1_1__leaf__0462_ _0319_ 0.00201f
C42366 _0229_ _0222_ 0
C42367 hold31/a_391_47# _0186_ 0
C42368 hold14/a_391_47# net28 0
C42369 _0343_ clknet_1_0__leaf__0460_ 0.57732f
C42370 _1051_/a_1059_315# _0180_ 0
C42371 net113 net156 0.07f
C42372 _0399_ _0303_ 0
C42373 _0820_/a_215_47# _0990_/a_27_47# 0
C42374 net48 _0902_/a_27_47# 0
C42375 A[12] A[9] 0.00159f
C42376 _1014_/a_634_159# _0112_ 0.00106f
C42377 net100 _0585_/a_27_297# 0.01477f
C42378 _0769_/a_299_297# _0773_/a_35_297# 0.07368f
C42379 VPWR _0172_ 1.95427f
C42380 acc0.A\[16\] net219 0
C42381 _0783_/a_79_21# _0783_/a_297_297# 0.01735f
C42382 net139 _0180_ 0
C42383 _1038_/a_381_47# net124 0
C42384 _1038_/a_891_413# net172 0
C42385 _0600_/a_253_47# _0352_ 0
C42386 _0765_/a_215_47# hold3/a_285_47# 0
C42387 net33 _1066_/a_891_413# 0.0436f
C42388 hold21/a_49_47# hold21/a_391_47# 0.00188f
C42389 _0255_ net9 0
C42390 hold46/a_391_47# _0548_/a_240_47# 0
C42391 hold24/a_49_47# _0208_ 0
C42392 _0718_/a_47_47# _0705_/a_59_75# 0.03737f
C42393 _0852_/a_285_297# _0218_ 0
C42394 _0341_ output41/a_27_47# 0
C42395 hold75/a_391_47# VPWR 0.17179f
C42396 _0283_ _0286_ 0.00667f
C42397 _0290_ _0090_ 0
C42398 _0750_/a_109_47# _0383_ 0
C42399 _0642_/a_27_413# _0825_/a_68_297# 0
C42400 control0.count\[2\] _0976_/a_76_199# 0
C42401 clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ 1.67674f
C42402 _0343_ _0221_ 0.45158f
C42403 clknet_1_0__leaf__0465_ _1044_/a_1017_47# 0
C42404 acc0.A\[4\] net10 0
C42405 _0088_ acc0.A\[6\] 0
C42406 net203 net106 0
C42407 hold81/a_49_47# _0345_ 0.00838f
C42408 hold16/a_49_47# _1030_/a_891_413# 0.00267f
C42409 _0129_ _1030_/a_27_47# 0
C42410 hold16/a_391_47# _1030_/a_466_413# 0
C42411 _1020_/a_466_413# net1 0.01108f
C42412 hold12/a_391_47# _1068_/a_891_413# 0
C42413 clknet_1_0__leaf__0462_ _0222_ 0.04597f
C42414 net168 _1052_/a_27_47# 0
C42415 _0997_/a_1059_315# net43 0.04443f
C42416 net198 hold51/a_391_47# 0.14808f
C42417 net18 hold51/a_285_47# 0
C42418 _0352_ _1006_/a_27_47# 0.02858f
C42419 _0732_/a_80_21# acc0.A\[23\] 0
C42420 VPWR _0995_/a_466_413# 0.25333f
C42421 output47/a_27_47# _0988_/a_1059_315# 0.00166f
C42422 _0443_ clkbuf_1_1__f__0458_/a_110_47# 0
C42423 _0285_ _0993_/a_193_47# 0
C42424 _0284_ _0993_/a_27_47# 0.02389f
C42425 _0751_/a_29_53# _0352_ 0
C42426 _0399_ _0281_ 0
C42427 _0304_ hold81/a_285_47# 0
C42428 net45 _0712_/a_465_47# 0
C42429 net188 _0156_ 0
C42430 _0225_ _0754_/a_149_47# 0.00445f
C42431 _1056_/a_27_47# _0820_/a_215_47# 0
C42432 net178 net47 0.02146f
C42433 hold13/a_285_47# net28 0
C42434 _0511_/a_299_297# _0187_ 0.00863f
C42435 _0347_ _0986_/a_466_413# 0
C42436 _0218_ net247 0
C42437 _1051_/a_27_47# _0525_/a_81_21# 0
C42438 hold28/a_285_47# _1048_/a_1059_315# 0.01349f
C42439 net150 clknet_1_0__leaf__0457_ 0.03697f
C42440 hold23/a_49_47# net170 0.04297f
C42441 _0550_/a_245_297# net180 0.00215f
C42442 _0550_/a_51_297# net30 0.15002f
C42443 net190 _1008_/a_466_413# 0
C42444 _0126_ _1008_/a_27_47# 0
C42445 net216 _1006_/a_381_47# 0
C42446 _0240_ _0775_/a_510_47# 0.0021f
C42447 _0104_ _1006_/a_466_413# 0.00875f
C42448 _0371_ _1006_/a_891_413# 0
C42449 _0533_/a_27_297# _0533_/a_109_47# 0.00393f
C42450 net227 _0725_/a_80_21# 0
C42451 _0726_/a_240_47# _0353_ 0
C42452 _0355_ _0725_/a_209_297# 0.02716f
C42453 _0354_ _0725_/a_209_47# 0
C42454 _0229_ net220 0
C42455 clkbuf_1_0__f__0460_/a_110_47# acc0.A\[23\] 0.00662f
C42456 _1048_/a_27_47# _0145_ 0
C42457 _1000_/a_1059_315# _0461_ 0.01053f
C42458 _0186_ _0524_/a_109_47# 0.00486f
C42459 _0762_/a_79_21# _0373_ 0
C42460 _0684_/a_145_75# acc0.A\[27\] 0
C42461 _0276_ _0347_ 0
C42462 _0195_ hold9/a_49_47# 0.03151f
C42463 _0250_ acc0.A\[23\] 0
C42464 _0546_/a_51_297# _0546_/a_240_47# 0.03076f
C42465 VPWR _1023_/a_193_47# 0.30466f
C42466 hold100/a_285_47# _0846_/a_51_297# 0
C42467 A[15] _0547_/a_68_297# 0
C42468 _0163_ hold93/a_391_47# 0
C42469 _0534_/a_384_47# _0180_ 0
C42470 net132 _0148_ 0
C42471 hold101/a_391_47# net63 0.00142f
C42472 net113 acc0.A\[26\] 0.25677f
C42473 _0991_/a_634_159# _0991_/a_466_413# 0.23992f
C42474 _0991_/a_193_47# _0991_/a_1059_315# 0.03405f
C42475 _0991_/a_27_47# _0991_/a_891_413# 0.03224f
C42476 _0534_/a_384_47# net218 0
C42477 net160 _0561_/a_51_297# 0
C42478 VPWR _0516_/a_373_47# 0.00142f
C42479 net84 _0399_ 0.11066f
C42480 _0367_ hold90/a_285_47# 0
C42481 _0315_ hold90/a_391_47# 0.00499f
C42482 _0726_/a_245_297# _0345_ 0
C42483 _0837_/a_81_21# clknet_1_1__leaf__0458_ 0
C42484 B[12] net20 0.00716f
C42485 _0794_/a_110_297# _0794_/a_27_47# 0
C42486 _1041_/a_634_159# net22 0
C42487 _0773_/a_35_297# _0392_ 0.16713f
C42488 _0195_ _1029_/a_27_47# 0
C42489 _0210_ _0957_/a_304_297# 0
C42490 _0554_/a_150_297# _0475_ 0
C42491 net61 hold18/a_285_47# 0
C42492 acc0.A\[19\] hold60/a_285_47# 0
C42493 _0216_ _0112_ 0.00757f
C42494 net10 _1045_/a_891_413# 0
C42495 _0982_/a_381_47# _1014_/a_1059_315# 0
C42496 clknet_1_1__leaf__0459_ _0811_/a_81_21# 0.00326f
C42497 _0502_/a_27_47# control0.sh 0
C42498 net160 _0133_ 0.00128f
C42499 _0573_/a_27_47# _0208_ 0
C42500 _1001_/a_193_47# _0183_ 0.01683f
C42501 _1001_/a_466_413# _0217_ 0.0012f
C42502 hold6/a_49_47# _1040_/a_466_413# 0
C42503 hold6/a_391_47# _1040_/a_193_47# 0
C42504 _0399_ _0996_/a_634_159# 0.03805f
C42505 _0294_ net229 0
C42506 acc0.A\[17\] _0306_ 0.197f
C42507 _0376_ clknet_1_0__leaf__0460_ 0.02644f
C42508 _0574_/a_27_297# acc0.A\[25\] 0.09452f
C42509 net176 net50 0.10783f
C42510 _1021_/a_27_47# _0217_ 0.02724f
C42511 _1021_/a_193_47# net150 0
C42512 hold54/a_285_47# hold54/a_391_47# 0.41909f
C42513 net36 _0171_ 0.10482f
C42514 hold35/a_49_47# _0154_ 0.37066f
C42515 comp0.B\[7\] hold46/a_49_47# 0
C42516 _1041_/a_634_159# clknet_1_0__leaf__0463_ 0.0011f
C42517 _0352_ _0737_/a_35_297# 0
C42518 _0558_/a_68_297# net160 0
C42519 _0854_/a_79_21# _0347_ 0.12365f
C42520 _0731_/a_81_21# _0326_ 0.1927f
C42521 net130 net73 0
C42522 _0125_ hold9/a_285_47# 0.00623f
C42523 _0174_ _0540_/a_240_47# 0.0162f
C42524 acc0.A\[20\] hold40/a_285_47# 0.09205f
C42525 _1058_/a_634_159# acc0.A\[10\] 0.00452f
C42526 hold44/a_285_47# _0354_ 0
C42527 hold44/a_49_47# _0355_ 0
C42528 _0343_ _0344_ 0.0748f
C42529 net48 _1023_/a_193_47# 0
C42530 _0366_ _1007_/a_592_47# 0.00263f
C42531 net223 _0771_/a_27_413# 0
C42532 clknet_0__0457_ _0178_ 0
C42533 _0163_ control0.reset 0
C42534 _0218_ _0841_/a_79_21# 0.00671f
C42535 _0155_ _0156_ 0
C42536 hold32/a_49_47# net142 0
C42537 _0953_/a_32_297# acc0.A\[15\] 0
C42538 _0258_ _0441_ 0
C42539 _0522_/a_27_297# net13 0.18725f
C42540 comp0.B\[2\] net26 0
C42541 _0800_/a_149_47# _0800_/a_240_47# 0.06872f
C42542 VPWR _0601_/a_68_297# 0.16722f
C42543 hold57/a_285_47# _0136_ 0.00359f
C42544 control0.add clknet_1_0__leaf__0457_ 0.68012f
C42545 net224 clkbuf_0__0462_/a_110_47# 0
C42546 net170 _0085_ 0
C42547 net234 _0345_ 0.03664f
C42548 VPWR _0697_/a_217_297# 0.18989f
C42549 _0401_ _0291_ 0.01199f
C42550 _0593_/a_113_47# net109 0
C42551 pp[17] _1031_/a_891_413# 0.00448f
C42552 _1002_/a_1059_315# _0352_ 0.02435f
C42553 net167 _1068_/a_193_47# 0
C42554 acc0.A\[16\] _0352_ 0.03179f
C42555 VPWR _0695_/a_472_297# 0.00853f
C42556 _1011_/a_193_47# _0350_ 0
C42557 hold29/a_285_47# _1023_/a_1059_315# 0
C42558 hold29/a_49_47# _1023_/a_891_413# 0.01541f
C42559 net58 _0181_ 0
C42560 control0.count\[3\] _0466_ 0.05382f
C42561 _0627_/a_369_297# _0254_ 0.00317f
C42562 _1004_/a_634_159# net52 0
C42563 _1033_/a_891_413# _1067_/a_27_47# 0
C42564 VPWR _1031_/a_466_413# 0.25531f
C42565 clkbuf_0__0465_/a_110_47# _0986_/a_466_413# 0.00899f
C42566 _0237_ _0382_ 0.02394f
C42567 _0673_/a_103_199# _0283_ 0
C42568 _0195_ _1019_/a_193_47# 0
C42569 net46 _0345_ 0.05277f
C42570 net178 _0988_/a_592_47# 0
C42571 _0216_ _0099_ 0
C42572 _0401_ _0991_/a_634_159# 0
C42573 _0290_ _0991_/a_466_413# 0
C42574 _0423_ _0991_/a_1059_315# 0
C42575 _0425_ _0991_/a_193_47# 0
C42576 _0325_ _1006_/a_1059_315# 0
C42577 _0176_ _1044_/a_27_47# 0
C42578 _0983_/a_592_47# _0399_ 0.00258f
C42579 hold68/a_49_47# net50 0.05399f
C42580 net167 _0478_ 0.01037f
C42581 net51 _1022_/a_975_413# 0.00109f
C42582 net205 _0208_ 0.06419f
C42583 _0502_/a_27_47# net157 0
C42584 _0835_/a_493_297# _0835_/a_215_47# 0
C42585 _0975_/a_59_75# control0.count\[0\] 0
C42586 _0955_/a_32_297# _0955_/a_220_297# 0.00132f
C42587 hold76/a_285_47# _0242_ 0.02753f
C42588 hold15/a_285_47# _0220_ 0.01285f
C42589 hold15/a_49_47# _0336_ 0
C42590 net247 _0177_ 0.06114f
C42591 _1038_/a_592_47# _0172_ 0
C42592 _0337_ hold80/a_49_47# 0
C42593 _0179_ _0143_ 0
C42594 net143 net37 0
C42595 _0216_ _0359_ 0
C42596 _1004_/a_466_413# clknet_1_0__leaf__0460_ 0.00684f
C42597 _1025_/a_634_159# acc0.A\[25\] 0.02139f
C42598 acc0.A\[13\] _0301_ 0.24207f
C42599 _1020_/a_27_47# _1015_/a_27_47# 0
C42600 _0343_ _0434_ 0.05464f
C42601 _0971_/a_384_47# _0880_/a_27_47# 0
C42602 hold21/a_49_47# _0519_/a_81_21# 0.00138f
C42603 net240 _1067_/a_27_47# 0
C42604 net55 pp[27] 0.00494f
C42605 clk rst 0.10672f
C42606 hold65/a_285_47# _0252_ 0
C42607 _0982_/a_1017_47# _0195_ 0
C42608 hold64/a_285_47# _0218_ 0
C42609 _0112_ net247 0
C42610 net54 _1008_/a_27_47# 0.006f
C42611 hold65/a_391_47# _0989_/a_891_413# 0.00206f
C42612 _0179_ _0988_/a_193_47# 0
C42613 _0180_ acc0.A\[8\] 0.00929f
C42614 hold20/a_391_47# _1072_/a_27_47# 0.0042f
C42615 hold20/a_285_47# _1072_/a_193_47# 0.0148f
C42616 _1001_/a_1059_315# control0.add 0
C42617 clkbuf_1_0__f__0457_/a_110_47# _1019_/a_466_413# 0
C42618 clknet_0__0457_ _1019_/a_27_47# 0.02693f
C42619 _0266_ acc0.A\[18\] 0
C42620 _0559_/a_51_297# comp0.B\[5\] 0.00282f
C42621 _0238_ _1006_/a_1059_315# 0
C42622 net63 _0369_ 0.06392f
C42623 net7 net153 0.00311f
C42624 _1021_/a_193_47# control0.add 0
C42625 _0119_ _1067_/a_1059_315# 0.00933f
C42626 clknet_0__0463_ net147 0
C42627 _0199_ comp0.B\[15\] 0.02596f
C42628 VPWR _0808_/a_585_47# 0
C42629 VPWR net79 0.42845f
C42630 _0473_ _0142_ 0.0264f
C42631 _1036_/a_27_47# _1036_/a_193_47# 0.97441f
C42632 _1055_/a_891_413# _0153_ 0.01248f
C42633 net217 hold70/a_391_47# 0.12951f
C42634 _0422_ hold70/a_285_47# 0.05108f
C42635 _0367_ clknet_0__0462_ 0
C42636 _1047_/a_634_159# acc0.A\[15\] 0
C42637 input3/a_75_212# net37 0
C42638 net77 _0268_ 0
C42639 net219 _0247_ 0.3845f
C42640 net231 clknet_1_0__leaf__0457_ 0
C42641 _0217_ hold19/a_49_47# 0
C42642 _0993_/a_193_47# _0218_ 0.01131f
C42643 _0994_/a_193_47# acc0.A\[13\] 0
C42644 net200 _0216_ 0
C42645 _0224_ clknet_1_0__leaf__0460_ 0.00342f
C42646 _0358_ _0685_/a_150_297# 0
C42647 _0523_/a_81_21# _0523_/a_299_297# 0.08213f
C42648 _0525_/a_299_297# net73 0.00196f
C42649 _0488_ clkbuf_1_0__f_clk/a_110_47# 0.01807f
C42650 _0387_ _0392_ 0.00734f
C42651 _0432_ acc0.A\[8\] 0
C42652 _0662_/a_299_297# _0181_ 0.00655f
C42653 output67/a_27_47# _0179_ 0
C42654 _0274_ _0831_/a_117_297# 0.0016f
C42655 hold101/a_285_47# clkbuf_1_0__f__0465_/a_110_47# 0.02314f
C42656 acc0.A\[16\] _1016_/a_975_413# 0.00171f
C42657 hold24/a_285_47# _0555_/a_51_297# 0
C42658 _0433_ _0826_/a_27_53# 0.13598f
C42659 _1041_/a_466_413# _0544_/a_51_297# 0
C42660 _0333_ clknet_1_1__leaf__0462_ 0.00579f
C42661 clknet_1_0__leaf__0463_ _1039_/a_1017_47# 0
C42662 hold54/a_285_47# _0182_ 0
C42663 _1050_/a_1059_315# _0524_/a_27_297# 0
C42664 A[15] net127 0.01732f
C42665 _1059_/a_634_159# clkbuf_0__0459_/a_110_47# 0.00238f
C42666 _1044_/a_891_413# _1044_/a_975_413# 0.00851f
C42667 _1044_/a_27_47# net130 0.22455f
C42668 _1044_/a_381_47# _1044_/a_561_413# 0.00123f
C42669 _0654_/a_207_413# _0808_/a_266_47# 0
C42670 comp0.B\[13\] _0954_/a_304_297# 0.01447f
C42671 _0274_ _0254_ 0.00335f
C42672 hold46/a_285_47# comp0.B\[12\] 0
C42673 net101 net157 0.0055f
C42674 _0529_/a_27_297# _0529_/a_109_47# 0.00393f
C42675 _0606_/a_215_297# _0383_ 0
C42676 _1038_/a_561_413# comp0.B\[6\] 0
C42677 _0504_/a_27_47# net36 0
C42678 hold52/a_391_47# net199 0.17257f
C42679 hold41/a_285_47# _1058_/a_891_413# 0
C42680 _0343_ acc0.A\[7\] 0
C42681 _0996_/a_27_47# _0345_ 0
C42682 _0343_ _0989_/a_1059_315# 0.00969f
C42683 _0343_ _0997_/a_27_47# 0.00277f
C42684 _0423_ _0425_ 0.11488f
C42685 _0290_ _0401_ 0.74206f
C42686 _0971_/a_299_297# _1062_/a_193_47# 0
C42687 VPWR _0743_/a_240_47# 0.00552f
C42688 _0946_/a_30_53# _0978_/a_27_297# 0
C42689 net173 _0206_ 0
C42690 net36 _1038_/a_634_159# 0.03978f
C42691 pp[0] _1038_/a_27_47# 0.00236f
C42692 clknet_1_1__leaf_clk _1065_/a_1059_315# 0.08177f
C42693 _0343_ hold94/a_285_47# 0
C42694 _0368_ _1007_/a_27_47# 0
C42695 net36 _0456_ 0.02017f
C42696 _0985_/a_634_159# acc0.A\[2\] 0
C42697 _0186_ _0142_ 0.00754f
C42698 _0382_ _1005_/a_27_47# 0
C42699 _0237_ _1005_/a_634_159# 0
C42700 _0216_ _1028_/a_466_413# 0
C42701 _0195_ _1028_/a_891_413# 0.04478f
C42702 hold42/a_49_47# hold42/a_391_47# 0.00188f
C42703 hold42/a_285_47# _1057_/a_1059_315# 0
C42704 _1057_/a_634_159# _1057_/a_381_47# 0
C42705 _0257_ _0838_/a_109_297# 0.00288f
C42706 _0756_/a_47_47# net51 0.00181f
C42707 hold48/a_391_47# hold49/a_391_47# 0
C42708 B[13] _1042_/a_193_47# 0
C42709 net125 clknet_0__0463_ 0
C42710 _0269_ _0986_/a_193_47# 0
C42711 _0984_/a_27_47# _0991_/a_27_47# 0.00131f
C42712 _0812_/a_510_47# _0288_ 0
C42713 net225 _1013_/a_1059_315# 0.00144f
C42714 _0111_ _1013_/a_634_159# 0.05396f
C42715 VPWR _1064_/a_1059_315# 0.44025f
C42716 _0552_/a_68_297# _0207_ 0.00181f
C42717 _0209_ _0549_/a_68_297# 0.00185f
C42718 _0334_ hold95/a_49_47# 0
C42719 net8 _0463_ 0.0221f
C42720 _1059_/a_634_159# _1059_/a_381_47# 0
C42721 _0789_/a_75_199# _0789_/a_201_297# 0.15956f
C42722 hold59/a_49_47# _0266_ 0
C42723 _1004_/a_1059_315# _0576_/a_27_297# 0
C42724 net248 _0271_ 0
C42725 pp[15] clknet_1_1__leaf__0459_ 0
C42726 net231 _1062_/a_466_413# 0
C42727 hold76/a_49_47# _0098_ 0
C42728 _0528_/a_81_21# _0528_/a_299_297# 0.08213f
C42729 _0181_ _0262_ 0
C42730 net208 _0128_ 0.44521f
C42731 _0982_/a_975_413# net247 0
C42732 input21/a_75_212# net10 0
C42733 _0346_ net5 0.34077f
C42734 VPWR hold2/a_285_47# 0.29485f
C42735 _0654_/a_207_413# _0345_ 0.00492f
C42736 _0820_/a_297_297# clknet_1_1__leaf__0465_ 0.00151f
C42737 _1065_/a_891_413# clkbuf_1_1__f_clk/a_110_47# 0.00708f
C42738 clknet_1_0__leaf__0458_ _0849_/a_79_21# 0.01259f
C42739 _0181_ _0582_/a_109_297# 0
C42740 clknet_0__0460_ _0318_ 0.0381f
C42741 net1 hold60/a_285_47# 0
C42742 comp0.B\[13\] _0540_/a_240_47# 0.00499f
C42743 hold46/a_391_47# _0202_ 0.00245f
C42744 net197 _0320_ 0
C42745 net100 _0112_ 0.03292f
C42746 net23 _0181_ 0.68173f
C42747 _0310_ _0246_ 0.07679f
C42748 _0783_/a_215_47# _0096_ 0.00317f
C42749 _0783_/a_510_47# _0399_ 0.00728f
C42750 init control0.sh 0
C42751 _0369_ _0812_/a_79_21# 0.11518f
C42752 _0751_/a_29_53# _0237_ 0
C42753 net242 _0333_ 0
C42754 hold8/a_285_47# acc0.A\[26\] 0.10539f
C42755 net44 _0129_ 0
C42756 _0984_/a_27_47# _0350_ 0
C42757 net233 _0846_/a_51_297# 0.1111f
C42758 _0427_ _0426_ 0
C42759 net61 _0846_/a_512_297# 0
C42760 net55 _0216_ 0
C42761 net64 _0432_ 0
C42762 acc0.A\[27\] _1028_/a_592_47# 0
C42763 hold33/a_49_47# comp0.B\[14\] 0
C42764 hold38/a_285_47# _1062_/a_466_413# 0
C42765 _0138_ _1046_/a_27_47# 0
C42766 hold16/a_285_47# VPWR 0.29965f
C42767 _0679_/a_68_297# _0371_ 0
C42768 control0.count\[2\] _0488_ 0.86489f
C42769 _0195_ _0739_/a_79_21# 0
C42770 _0144_ net7 0.00159f
C42771 _0118_ net1 0.02445f
C42772 net155 _0347_ 0
C42773 _1052_/a_891_413# _0186_ 0
C42774 _0707_/a_75_199# hold62/a_285_47# 0
C42775 net186 _1033_/a_891_413# 0
C42776 _0388_ clkbuf_1_0__f__0461_/a_110_47# 0
C42777 _1056_/a_27_47# _1055_/a_891_413# 0
C42778 _1056_/a_193_47# _1055_/a_1059_315# 0
C42779 _1058_/a_634_159# _0188_ 0
C42780 _0433_ _0087_ 0
C42781 _0501_/a_27_47# clkbuf_0__0463_/a_110_47# 0.01036f
C42782 _0972_/a_256_47# net17 0.00259f
C42783 clkbuf_1_0__f__0464_/a_110_47# _1048_/a_891_413# 0.00189f
C42784 _0612_/a_59_75# acc0.A\[18\] 0.13256f
C42785 _1014_/a_891_413# clkbuf_0__0457_/a_110_47# 0
C42786 _0733_/a_79_199# hold90/a_49_47# 0
C42787 _0107_ hold69/a_285_47# 0
C42788 net30 _0172_ 0.1481f
C42789 acc0.A\[1\] _0182_ 0.40479f
C42790 _0533_/a_109_47# _0199_ 0.00281f
C42791 _1000_/a_27_47# _0459_ 0
C42792 hold66/a_391_47# net51 0.0036f
C42793 _0218_ net148 0
C42794 _0349_ _0108_ 0
C42795 clknet_0__0463_ _0473_ 0.47025f
C42796 _0183_ _1060_/a_561_413# 0
C42797 clkbuf_1_1__f__0463_/a_110_47# _0475_ 0.00247f
C42798 clknet_0__0458_ hold86/a_285_47# 0
C42799 input31/a_75_212# _0546_/a_51_297# 0
C42800 control0.state\[0\] _1063_/a_27_47# 0
C42801 hold47/a_285_47# net12 0
C42802 hold87/a_391_47# _0264_ 0.01376f
C42803 _0217_ _0241_ 0
C42804 _0123_ _1024_/a_466_413# 0
C42805 clknet_1_0__leaf__0462_ _1022_/a_466_413# 0.00604f
C42806 net108 _1022_/a_193_47# 0.01325f
C42807 net192 acc0.A\[11\] 0.03677f
C42808 hold23/a_285_47# _0449_ 0
C42809 _1005_/a_27_47# _1005_/a_634_159# 0.14145f
C42810 _0978_/a_109_297# _0485_ 0
C42811 _0978_/a_27_297# _0487_ 0
C42812 _0383_ hold3/a_49_47# 0.00285f
C42813 _0369_ hold3/a_391_47# 0
C42814 _0240_ _0347_ 0.09856f
C42815 _1031_/a_381_47# _0567_/a_27_297# 0
C42816 _0247_ _0352_ 0.12257f
C42817 _0376_ hold94/a_285_47# 0
C42818 _0604_/a_113_47# _0460_ 0
C42819 _0369_ _0347_ 0.06353f
C42820 net117 _1013_/a_27_47# 0
C42821 _0546_/a_512_297# _0139_ 0
C42822 hold75/a_285_47# hold75/a_391_47# 0.41909f
C42823 _1047_/a_891_413# clknet_1_1__leaf__0457_ 0.01899f
C42824 comp0.B\[4\] _0175_ 0.33245f
C42825 clkbuf_1_0__f__0457_/a_110_47# _0352_ 0.00509f
C42826 _0984_/a_1059_315# _0849_/a_79_21# 0.00195f
C42827 control0.state\[0\] _0974_/a_448_47# 0
C42828 hold45/a_285_47# VPWR 0.27802f
C42829 net149 _0580_/a_109_47# 0.00338f
C42830 _0346_ acc0.A\[11\] 0
C42831 _0991_/a_634_159# _0089_ 0.02375f
C42832 _0991_/a_466_413# net77 0
C42833 net160 _0208_ 0.11562f
C42834 control0.state\[1\] clknet_1_0__leaf__0457_ 0.00308f
C42835 _0354_ _0219_ 0.53281f
C42836 _0536_/a_240_47# net134 0
C42837 _0297_ _0300_ 0.24174f
C42838 net53 hold90/a_49_47# 0.3208f
C42839 hold96/a_285_47# _0347_ 0
C42840 _0817_/a_368_297# _0294_ 0
C42841 clknet_1_1__leaf__0465_ _0219_ 0.05685f
C42842 _0104_ _0369_ 0.04206f
C42843 _0260_ _0256_ 0.02567f
C42844 _0985_/a_27_47# _0261_ 0.00607f
C42845 _0985_/a_193_47# _0262_ 0
C42846 _0461_ net201 0
C42847 _0283_ net79 0
C42848 _0286_ _0808_/a_266_47# 0.00554f
C42849 _0583_/a_27_297# _1060_/a_193_47# 0
C42850 _0216_ _1029_/a_592_47# 0
C42851 hold52/a_391_47# VPWR 0.18714f
C42852 _0728_/a_59_75# _0354_ 0.00361f
C42853 clknet_1_1__leaf__0459_ _0992_/a_634_159# 0.01644f
C42854 _0603_/a_68_297# _0460_ 0.01488f
C42855 _0214_ _0493_/a_27_47# 0
C42856 _0563_/a_149_47# _0171_ 0
C42857 _0730_/a_215_47# _0317_ 0
C42858 _0460_ hold73/a_391_47# 0.00604f
C42859 _0982_/a_975_413# net100 0
C42860 VPWR _1065_/a_891_413# 0.18211f
C42861 _0174_ _0542_/a_512_297# 0
C42862 _0600_/a_253_297# _0600_/a_253_47# 0.00137f
C42863 _0159_ _1046_/a_381_47# 0
C42864 hold6/a_49_47# net174 0
C42865 net14 net138 0
C42866 _1038_/a_1059_315# comp0.B\[4\] 0
C42867 _0995_/a_634_159# _0995_/a_466_413# 0.23992f
C42868 _0995_/a_193_47# _0995_/a_1059_315# 0.03405f
C42869 _0995_/a_27_47# _0995_/a_891_413# 0.03224f
C42870 _0529_/a_109_297# net170 0.00518f
C42871 _0412_ _0300_ 0
C42872 clknet_1_0__leaf__0457_ _0610_/a_145_75# 0
C42873 _0419_ _0418_ 0.09863f
C42874 _0091_ _0281_ 0.15526f
C42875 hold87/a_285_47# clknet_1_0__leaf__0458_ 0.00408f
C42876 _1002_/a_1059_315# _0237_ 0
C42877 _1060_/a_561_413# acc0.A\[15\] 0
C42878 _1002_/a_891_413# _0381_ 0
C42879 net62 _0444_ 0
C42880 output59/a_27_47# hold95/a_49_47# 0
C42881 _0693_/a_68_297# _0219_ 0.00807f
C42882 _0450_ _0444_ 0
C42883 net144 acc0.A\[10\] 0
C42884 clknet_1_0__leaf__0458_ _0529_/a_27_297# 0
C42885 _0174_ acc0.A\[15\] 0
C42886 net36 _0550_/a_149_47# 0
C42887 hold9/a_391_47# _1027_/a_193_47# 0.00107f
C42888 hold9/a_285_47# _1027_/a_634_159# 0
C42889 hold9/a_49_47# _1027_/a_466_413# 0.01453f
C42890 VPWR _0819_/a_299_297# 0.19617f
C42891 _0232_ _0350_ 0
C42892 _0803_/a_68_297# _0399_ 0.00723f
C42893 net152 _1042_/a_27_47# 0
C42894 net53 _1007_/a_381_47# 0
C42895 acc0.A\[21\] hold66/a_49_47# 0
C42896 _1070_/a_1059_315# _1069_/a_1059_315# 0.00819f
C42897 net13 _0193_ 0.02203f
C42898 hold45/a_285_47# input4/a_75_212# 0
C42899 _0183_ _0208_ 0.00447f
C42900 control0.state\[1\] _1062_/a_466_413# 0.01258f
C42901 _0243_ _0611_/a_68_297# 0.10698f
C42902 control0.state\[0\] _1062_/a_1059_315# 0.13368f
C42903 _0982_/a_193_47# _0217_ 0
C42904 VPWR _0836_/a_150_297# 0.002f
C42905 _1034_/a_891_413# _0957_/a_32_297# 0
C42906 net78 acc0.A\[9\] 0
C42907 clknet_0__0465_ acc0.A\[9\] 0.00914f
C42908 net82 net43 0
C42909 net54 _0688_/a_109_297# 0
C42910 hold25/a_285_47# input8/a_75_212# 0
C42911 _1011_/a_634_159# _1011_/a_381_47# 0
C42912 _0286_ _0345_ 0.27419f
C42913 net50 _1023_/a_466_413# 0
C42914 _0985_/a_27_47# _0509_/a_27_47# 0.00808f
C42915 _1016_/a_891_413# _0369_ 0.04337f
C42916 net188 output37/a_27_47# 0
C42917 hold41/a_391_47# pp[10] 0
C42918 VPWR _0437_ 0.25397f
C42919 _0171_ _1061_/a_27_47# 0
C42920 _0133_ _1034_/a_193_47# 0.01704f
C42921 _0343_ output43/a_27_47# 0.02382f
C42922 _0643_/a_253_47# _0446_ 0
C42923 clknet_1_0__leaf__0464_ _0181_ 0
C42924 _1034_/a_891_413# net23 0
C42925 hold85/a_285_47# _0164_ 0.00322f
C42926 clknet_0__0465_ _0986_/a_592_47# 0
C42927 acc0.A\[22\] pp[23] 0.00183f
C42928 _0289_ _0992_/a_193_47# 0
C42929 _0287_ _0992_/a_27_47# 0
C42930 net45 _0997_/a_634_159# 0.00145f
C42931 acc0.A\[12\] _0278_ 0.07245f
C42932 _0290_ _0089_ 0.01966f
C42933 _1021_/a_1059_315# hold73/a_285_47# 0.00341f
C42934 _0195_ _1025_/a_193_47# 0
C42935 _1055_/a_193_47# VPWR 0.35799f
C42936 clknet_1_0__leaf__0462_ net243 0.04776f
C42937 _1020_/a_975_413# VPWR 0.00528f
C42938 VPWR _0791_/a_199_47# 0
C42939 _1001_/a_27_47# acc0.A\[19\] 0
C42940 _1026_/a_1059_315# _0687_/a_59_75# 0
C42941 _1003_/a_27_47# VPWR 0.6929f
C42942 hold65/a_49_47# _0831_/a_35_297# 0.02391f
C42943 _0982_/a_891_413# _0580_/a_27_297# 0
C42944 _0982_/a_1059_315# _0580_/a_109_297# 0
C42945 _0163_ _1063_/a_193_47# 0
C42946 _0181_ _1063_/a_466_413# 0
C42947 _0837_/a_81_21# _0218_ 0.0209f
C42948 _0399_ acc0.A\[18\] 0.03888f
C42949 clk control0.state\[2\] 0.55361f
C42950 _0955_/a_220_297# _0474_ 0
C42951 _0567_/a_27_297# _0219_ 0
C42952 net57 hold95/a_391_47# 0.00227f
C42953 _0195_ hold95/a_285_47# 0.02416f
C42954 hold44/a_49_47# _0127_ 0.31186f
C42955 _0404_ _0297_ 0.38442f
C42956 _0241_ _0248_ 0.20574f
C42957 clkbuf_0__0465_/a_110_47# _0369_ 0
C42958 _0794_/a_27_47# _0345_ 0.00425f
C42959 _0292_ _0428_ 0.00137f
C42960 _0966_/a_27_47# _0488_ 0.00758f
C42961 _0292_ _0660_/a_113_47# 0.01015f
C42962 _1023_/a_27_47# _1023_/a_193_47# 0.97064f
C42963 _0163_ _0460_ 0
C42964 _0217_ _0450_ 0
C42965 net248 clknet_1_0__leaf__0465_ 0.13833f
C42966 _0221_ _0568_/a_27_297# 0
C42967 _1042_/a_27_47# _1042_/a_466_413# 0.26005f
C42968 _1042_/a_193_47# _1042_/a_634_159# 0.11897f
C42969 _0511_/a_299_297# clknet_1_1__leaf__0465_ 0
C42970 acc0.A\[14\] _0790_/a_35_297# 0.00247f
C42971 _0181_ _1060_/a_466_413# 0.04012f
C42972 _0486_ net159 0.09726f
C42973 net44 hold61/a_285_47# 0.00104f
C42974 B[12] B[9] 0.00134f
C42975 clknet_1_1__leaf_clk hold93/a_49_47# 0.00126f
C42976 _0179_ _0174_ 0
C42977 _1037_/a_1059_315# _0552_/a_68_297# 0.00124f
C42978 clkbuf_1_0__f__0457_/a_110_47# net207 0.00102f
C42979 _1010_/a_466_413# _0352_ 0.01904f
C42980 _1010_/a_381_47# _0347_ 0.00416f
C42981 _0401_ _0656_/a_59_75# 0
C42982 _0216_ _0238_ 0.02704f
C42983 _0174_ B[14] 0
C42984 _0459_ _0507_/a_27_297# 0.01609f
C42985 _0531_/a_109_297# _0465_ 0.00179f
C42986 _1051_/a_381_47# clknet_1_1__leaf__0464_ 0.00101f
C42987 hold63/a_49_47# _0124_ 0.04134f
C42988 _0412_ _0404_ 0.03169f
C42989 _0179_ _1050_/a_27_47# 0.02096f
C42990 _0800_/a_51_297# _0219_ 0.25991f
C42991 _0800_/a_240_47# _0345_ 0
C42992 _1045_/a_975_413# clknet_1_1__leaf__0464_ 0
C42993 _0458_ _0844_/a_297_47# 0.00253f
C42994 _1039_/a_27_47# _0171_ 0
C42995 _1036_/a_466_413# _1036_/a_592_47# 0.00553f
C42996 _1036_/a_634_159# _1036_/a_1017_47# 0
C42997 _0714_/a_245_297# _0339_ 0
C42998 _0401_ _0986_/a_1059_315# 0
C42999 _0346_ _0990_/a_561_413# 0
C43000 pp[30] hold62/a_49_47# 0.00658f
C43001 acc0.A\[2\] _0531_/a_109_297# 0
C43002 hold26/a_391_47# _0172_ 0.0063f
C43003 _0459_ net165 0
C43004 _0578_/a_109_47# net187 0
C43005 _0644_/a_377_297# _0276_ 0.00215f
C43006 _0684_/a_59_75# _0315_ 0
C43007 _0767_/a_59_75# _0679_/a_68_297# 0.00598f
C43008 _1003_/a_27_47# net48 0
C43009 _0725_/a_209_47# _0353_ 0.00623f
C43010 VPWR _1040_/a_193_47# 0.30112f
C43011 clknet_0__0463_ _0497_/a_68_297# 0
C43012 hold27/a_49_47# net7 0.03325f
C43013 _0966_/a_109_297# net236 0
C43014 _0997_/a_27_47# _0793_/a_51_297# 0
C43015 _0458_ _1048_/a_1059_315# 0
C43016 _1050_/a_1059_315# _0194_ 0
C43017 _0227_ _0217_ 0.0336f
C43018 net238 net42 0.01897f
C43019 _0366_ _0758_/a_79_21# 0
C43020 A[12] _0515_/a_299_297# 0
C43021 pp[0] B[6] 0.1836f
C43022 output37/a_27_47# _0155_ 0.00752f
C43023 _0350_ _0321_ 0
C43024 _1011_/a_27_47# _0334_ 0
C43025 hold13/a_285_47# clknet_0__0463_ 0.00161f
C43026 hold49/a_285_47# net19 0
C43027 hold49/a_391_47# net195 0
C43028 clkbuf_0__0460_/a_110_47# _0350_ 0
C43029 _1002_/a_27_47# _0765_/a_79_21# 0
C43030 _0305_ _0775_/a_79_21# 0
C43031 _0576_/a_373_47# VPWR 0
C43032 _0163_ _1062_/a_891_413# 0.00139f
C43033 _0992_/a_1059_315# _0282_ 0
C43034 clknet_1_0__leaf__0462_ _1024_/a_381_47# 0
C43035 _0467_ _1063_/a_381_47# 0.00736f
C43036 _1058_/a_891_413# net4 0.04631f
C43037 _1058_/a_466_413# _0187_ 0
C43038 hold59/a_49_47# _0399_ 0.0076f
C43039 _0092_ net39 0.39631f
C43040 _0459_ acc0.A\[19\] 0.10516f
C43041 _0958_/a_27_47# _0164_ 0.00107f
C43042 _0477_ _0972_/a_250_297# 0
C43043 hold32/a_391_47# net47 0
C43044 net58 _0990_/a_193_47# 0
C43045 _0346_ _0303_ 0.03235f
C43046 _1032_/a_27_47# _1067_/a_193_47# 0.00135f
C43047 _1032_/a_193_47# _1067_/a_27_47# 0
C43048 _0467_ _0959_/a_472_297# 0.00404f
C43049 _0777_/a_377_297# _0395_ 0.00188f
C43050 net36 net124 0.10332f
C43051 _0197_ _0261_ 0.00101f
C43052 _1049_/a_1017_47# _0465_ 0
C43053 _0476_ hold39/a_391_47# 0
C43054 _0902_/a_27_47# _0345_ 0
C43055 _0329_ _0109_ 0
C43056 _0428_ _0990_/a_975_413# 0.0014f
C43057 _0216_ _0721_/a_27_47# 0
C43058 _1012_/a_1059_315# net239 0.00414f
C43059 _0381_ _0103_ 0
C43060 _0237_ net91 0.00859f
C43061 _0351_ _0350_ 0.10512f
C43062 _1054_/a_193_47# acc0.A\[7\] 0
C43063 _0179_ _0518_/a_27_297# 0.0078f
C43064 _1054_/a_1059_315# hold1/a_285_47# 0
C43065 _1054_/a_891_413# _0989_/a_27_47# 0
C43066 _1054_/a_1059_315# _0989_/a_193_47# 0
C43067 _0795_/a_81_21# net41 0.02579f
C43068 net197 hold8/a_49_47# 0
C43069 hold42/a_391_47# net189 0.1316f
C43070 clkbuf_1_1__f__0463_/a_110_47# _1033_/a_193_47# 0.01336f
C43071 _0311_ _0614_/a_29_53# 0
C43072 _1057_/a_891_413# net189 0.00258f
C43073 _0626_/a_68_297# VPWR 0.15477f
C43074 hold10/a_391_47# control0.sh 0
C43075 clkbuf_0__0463_/a_110_47# _0498_/a_240_47# 0
C43076 _0463_ _0498_/a_245_297# 0
C43077 _1053_/a_193_47# _1052_/a_193_47# 0
C43078 _1053_/a_27_47# _1052_/a_634_159# 0
C43079 _0579_/a_109_297# net211 0.0015f
C43080 _0550_/a_51_297# _1040_/a_27_47# 0.00841f
C43081 _0789_/a_315_47# _0298_ 0.00567f
C43082 _1059_/a_381_47# net145 0
C43083 _0093_ _0995_/a_1059_315# 0
C43084 VPWR _0301_ 0.35754f
C43085 _0789_/a_201_297# _0345_ 0
C43086 _0754_/a_51_297# _0754_/a_240_47# 0.03076f
C43087 _0640_/a_215_297# _0433_ 0
C43088 _0643_/a_103_199# _0256_ 0
C43089 _0951_/a_209_311# _0161_ 0.07169f
C43090 _0421_ hold81/a_285_47# 0.00315f
C43091 net231 _0160_ 0.03611f
C43092 net165 _0265_ 0.12943f
C43093 _0346_ _0281_ 0.0155f
C43094 _0673_/a_103_199# _0345_ 0.01001f
C43095 _0785_/a_81_21# _0346_ 0
C43096 net167 VPWR 0.30905f
C43097 _0221_ _0109_ 0.00336f
C43098 _1055_/a_1059_315# clknet_1_1__leaf__0465_ 0
C43099 net211 _0399_ 0
C43100 net15 net148 0
C43101 _0672_/a_79_21# _0345_ 0.00402f
C43102 hold11/a_49_47# clknet_1_0__leaf__0465_ 0.04184f
C43103 _0757_/a_68_297# net90 0
C43104 _0562_/a_68_297# _0562_/a_150_297# 0.00477f
C43105 _0710_/a_109_47# _0342_ 0.00414f
C43106 _0176_ _1042_/a_381_47# 0
C43107 _0779_/a_297_297# _0352_ 0.00209f
C43108 _0323_ _0462_ 0.0284f
C43109 net1 clknet_1_0__leaf_clk 0
C43110 _0673_/a_337_297# _0295_ 0.00985f
C43111 _0555_/a_51_297# _0210_ 0.12491f
C43112 _0555_/a_245_297# net160 0
C43113 _0663_/a_27_413# _0288_ 0.23494f
C43114 net14 hold83/a_285_47# 0
C43115 net193 _0142_ 0
C43116 input24/a_75_212# control0.sh 0
C43117 _1051_/a_193_47# _0524_/a_27_297# 0
C43118 _1051_/a_27_47# _0524_/a_109_297# 0
C43119 _0672_/a_510_47# _0296_ 0.00217f
C43120 clkload3/a_268_47# _0459_ 0
C43121 _0455_ _0849_/a_79_21# 0
C43122 _0992_/a_466_413# _0281_ 0
C43123 input20/a_75_212# net198 0
C43124 hold23/a_285_47# _0260_ 0
C43125 _1030_/a_1017_47# clknet_1_1__leaf__0462_ 0
C43126 net8 clkbuf_1_0__f__0463_/a_110_47# 0
C43127 _0971_/a_299_297# net17 0.00102f
C43128 _1053_/a_193_47# net12 0.04156f
C43129 clknet_0__0458_ _0458_ 0.00559f
C43130 _0536_/a_240_47# net22 0.05884f
C43131 net2 _0369_ 0.00193f
C43132 _0265_ acc0.A\[19\] 0
C43133 net47 _0242_ 0
C43134 net34 hold85/a_285_47# 0
C43135 control0.state\[1\] hold85/a_391_47# 0
C43136 A[3] A[2] 0.2436f
C43137 _0197_ _0509_/a_27_47# 0
C43138 _0530_/a_81_21# _0186_ 0.0025f
C43139 VPWR _0994_/a_193_47# 0.31875f
C43140 _0974_/a_448_47# _1068_/a_193_47# 0
C43141 _0125_ acc0.A\[28\] 0
C43142 _0852_/a_285_297# _0268_ 0
C43143 VPWR _1008_/a_1017_47# 0
C43144 net118 clknet_1_0__leaf__0461_ 0.01898f
C43145 _0981_/a_109_297# clknet_0_clk 0
C43146 clknet_1_0__leaf__0462_ _0366_ 0.03419f
C43147 hold43/a_391_47# VPWR 0.19732f
C43148 _0461_ _1015_/a_193_47# 0.03883f
C43149 _1034_/a_1059_315# _0959_/a_80_21# 0
C43150 clkload2/a_268_47# clkload2/Y 0.00587f
C43151 _0576_/a_27_297# net176 0.06821f
C43152 _0338_ hold62/a_285_47# 0
C43153 _0339_ hold62/a_49_47# 0.00253f
C43154 _0278_ net42 0
C43155 _0697_/a_80_21# _0697_/a_217_297# 0.12661f
C43156 clknet_1_0__leaf__0458_ _0199_ 0
C43157 _0785_/a_299_297# _0428_ 0.02209f
C43158 _0785_/a_384_47# _0427_ 0
C43159 _0341_ _1013_/a_891_413# 0
C43160 _0340_ _1013_/a_1059_315# 0
C43161 hold10/a_391_47# net157 0.16434f
C43162 net144 _0188_ 0
C43163 _0961_/a_113_297# clknet_1_0__leaf_clk 0
C43164 clknet_1_0__leaf__0463_ _0536_/a_240_47# 0.00131f
C43165 clknet_0__0463_ _0132_ 0
C43166 _0305_ _0158_ 0
C43167 VPWR hold93/a_285_47# 0.2925f
C43168 comp0.B\[4\] _0955_/a_114_297# 0.01339f
C43169 _0174_ _0544_/a_51_297# 0.13809f
C43170 _0521_/a_81_21# _0179_ 0.00607f
C43171 _0695_/a_217_297# _0695_/a_472_297# 0.00517f
C43172 _0695_/a_80_21# _0695_/a_300_47# 0.00997f
C43173 _0820_/a_79_21# _0399_ 0.20197f
C43174 _1009_/a_27_47# _0350_ 0.00164f
C43175 _0222_ _0600_/a_253_47# 0
C43176 _1010_/a_1059_315# hold95/a_391_47# 0.01554f
C43177 _0268_ net247 0
C43178 _0307_ _0218_ 0.05067f
C43179 comp0.B\[10\] _0544_/a_512_297# 0.00275f
C43180 _1031_/a_634_159# _1031_/a_466_413# 0.23992f
C43181 _1031_/a_193_47# _1031_/a_1059_315# 0.03405f
C43182 _1031_/a_27_47# _1031_/a_891_413# 0.03224f
C43183 _0247_ hold72/a_285_47# 0
C43184 _0227_ _0248_ 0
C43185 VPWR _0214_ 0.5027f
C43186 net31 _0205_ 0
C43187 _0996_/a_634_159# _0346_ 0
C43188 hold30/a_391_47# net243 0
C43189 _0804_/a_297_297# _0403_ 0.00641f
C43190 net105 _1014_/a_1017_47# 0
C43191 _1000_/a_193_47# _0218_ 0
C43192 output42/a_27_47# _0995_/a_27_47# 0
C43193 hold53/a_391_47# acc0.A\[24\] 0
C43194 _0123_ _0122_ 0
C43195 clknet_1_0__leaf__0462_ net151 0.05274f
C43196 _1005_/a_381_47# _1005_/a_561_413# 0.00123f
C43197 _1005_/a_27_47# net91 0.26778f
C43198 _1005_/a_891_413# _1005_/a_975_413# 0.00851f
C43199 clkbuf_0__0458_/a_110_47# _0986_/a_193_47# 0
C43200 _0244_ _0616_/a_493_297# 0
C43201 hold66/a_285_47# net49 0.00486f
C43202 hold55/a_49_47# _0183_ 0
C43203 _0519_/a_299_297# _0152_ 0.00163f
C43204 control0.add _0246_ 0
C43205 VPWR _0729_/a_68_297# 0.17028f
C43206 _0984_/a_891_413# _0082_ 0.0094f
C43207 _0984_/a_975_413# net222 0
C43208 net230 net12 0.00369f
C43209 _1013_/a_466_413# _1013_/a_561_413# 0.00772f
C43210 _1013_/a_634_159# _1013_/a_975_413# 0
C43211 _0200_ clknet_0__0463_ 0
C43212 _0751_/a_29_53# _0222_ 0.06259f
C43213 _0991_/a_1017_47# net67 0
C43214 net77 _0089_ 0.00186f
C43215 _0251_ _0438_ 0.05501f
C43216 VPWR _0853_/a_68_297# 0.14374f
C43217 _1002_/a_193_47# _1002_/a_891_413# 0.19489f
C43218 _1002_/a_27_47# _1002_/a_381_47# 0.06222f
C43219 _1002_/a_634_159# _1002_/a_1059_315# 0
C43220 hold68/a_49_47# _0576_/a_27_297# 0
C43221 _1027_/a_193_47# _0739_/a_215_47# 0
C43222 _1027_/a_466_413# _0739_/a_79_21# 0
C43223 _0985_/a_27_47# hold28/a_285_47# 0
C43224 _0985_/a_193_47# hold28/a_49_47# 0
C43225 _0595_/a_109_297# _0486_ 0
C43226 _0984_/a_634_159# clknet_1_0__leaf__0458_ 0.01043f
C43227 _1027_/a_1059_315# _0347_ 0
C43228 _0462_ net237 0.00256f
C43229 net22 _1046_/a_27_47# 0
C43230 _1017_/a_891_413# net43 0.00126f
C43231 _0118_ net157 0
C43232 net165 _1060_/a_381_47# 0
C43233 _0114_ _1060_/a_193_47# 0
C43234 _0389_ _0461_ 0.00411f
C43235 clknet_0__0463_ comp0.B\[8\] 0.01122f
C43236 _0612_/a_59_75# _0611_/a_150_297# 0
C43237 VPWR _0252_ 1.0308f
C43238 B[7] A[15] 0.14898f
C43239 _0108_ _1012_/a_193_47# 0
C43240 hold35/a_391_47# _1055_/a_193_47# 0
C43241 _0372_ _0245_ 0
C43242 VPWR _0989_/a_381_47# 0.07788f
C43243 VPWR _0997_/a_634_159# 0.19229f
C43244 net36 _0464_ 0
C43245 _0795_/a_384_47# _0405_ 0.01047f
C43246 _0274_ _0273_ 0.01017f
C43247 _0795_/a_299_297# _0400_ 0.00104f
C43248 _0174_ _0141_ 0.00116f
C43249 _1038_/a_891_413# _1040_/a_891_413# 0
C43250 _1059_/a_27_47# _0369_ 0.02476f
C43251 _0217_ _1019_/a_466_413# 0.00842f
C43252 _0183_ _1019_/a_193_47# 0.03301f
C43253 _0690_/a_150_297# _0319_ 0.00157f
C43254 _0153_ net47 0
C43255 _0834_/a_109_297# clknet_1_1__leaf__0458_ 0
C43256 VPWR _0992_/a_381_47# 0.07682f
C43257 B[13] clknet_1_1__leaf__0464_ 0.00618f
C43258 hold56/a_285_47# net186 0
C43259 net203 hold39/a_285_47# 0
C43260 _0734_/a_285_47# _0361_ 0.06861f
C43261 control0.state\[1\] _0958_/a_109_47# 0.00109f
C43262 control0.state\[0\] _0958_/a_197_47# 0
C43263 hold35/a_49_47# net181 0.00296f
C43264 _0154_ _0515_/a_299_297# 0.00152f
C43265 _1035_/a_193_47# _0175_ 0.02573f
C43266 _0765_/a_215_47# _0765_/a_510_47# 0.00529f
C43267 _0503_/a_109_297# clknet_1_0__leaf__0461_ 0
C43268 output56/a_27_47# _1011_/a_466_413# 0
C43269 hold20/a_49_47# _0486_ 0.00124f
C43270 VPWR _1061_/a_1059_315# 0.46203f
C43271 hold23/a_391_47# _0447_ 0
C43272 _0305_ acc0.A\[14\] 0.23086f
C43273 _0580_/a_27_297# clkbuf_0__0457_/a_110_47# 0.00428f
C43274 clknet_1_0__leaf__0463_ _1046_/a_27_47# 0.00115f
C43275 _0201_ _0537_/a_68_297# 0.10723f
C43276 net58 _0438_ 0.02552f
C43277 _0355_ _0703_/a_109_297# 0
C43278 _0636_/a_145_75# _0465_ 0
C43279 _0350_ _0771_/a_27_413# 0
C43280 VPWR _0207_ 0.38048f
C43281 _1034_/a_1059_315# _0173_ 0.00771f
C43282 _1034_/a_193_47# _0208_ 0
C43283 _1034_/a_891_413# _0213_ 0
C43284 acc0.A\[12\] _0512_/a_109_297# 0
C43285 hold87/a_391_47# _0454_ 0
C43286 _1035_/a_634_159# control0.sh 0
C43287 _0217_ net219 0.24353f
C43288 hold9/a_49_47# net156 0
C43289 clknet_0__0458_ clkbuf_1_1__f__0458_/a_110_47# 0.34209f
C43290 net58 _0636_/a_59_75# 0
C43291 _0800_/a_51_297# _0799_/a_209_297# 0
C43292 net32 _1042_/a_1017_47# 0
C43293 net165 _0267_ 0.04851f
C43294 acc0.A\[17\] net221 0
C43295 hold54/a_391_47# _0216_ 0
C43296 A[12] net192 0
C43297 _1018_/a_975_413# _0459_ 0
C43298 control0.count\[1\] _1069_/a_634_159# 0.01301f
C43299 _1070_/a_634_159# control0.count\[0\] 0
C43300 _0168_ _1069_/a_891_413# 0.00208f
C43301 _1070_/a_381_47# clknet_1_0__leaf_clk 0
C43302 VPWR _1069_/a_561_413# 0.0034f
C43303 control0.state\[1\] _0160_ 0
C43304 pp[6] hold31/a_285_47# 0
C43305 hold27/a_391_47# _0138_ 0.04027f
C43306 _0398_ _0219_ 0
C43307 _1056_/a_1059_315# _1058_/a_27_47# 0
C43308 _1056_/a_27_47# _1058_/a_1059_315# 0
C43309 _1011_/a_381_47# net97 0
C43310 _1011_/a_634_159# net57 0
C43311 output50/a_27_47# acc0.A\[23\] 0
C43312 net50 net177 0.00469f
C43313 _0195_ _1011_/a_193_47# 0
C43314 _0985_/a_381_47# _0186_ 0.01243f
C43315 _1000_/a_891_413# _0614_/a_29_53# 0
C43316 _1055_/a_466_413# A[9] 0
C43317 _0399_ _0669_/a_29_53# 0.01406f
C43318 _0216_ clkbuf_1_0__f__0461_/a_110_47# 0.02471f
C43319 _0374_ net51 0.16264f
C43320 _0343_ _0748_/a_81_21# 0.00356f
C43321 net243 _0574_/a_373_47# 0
C43322 _0182_ _0198_ 0.3239f
C43323 _1006_/a_466_413# _1006_/a_381_47# 0.03733f
C43324 _1006_/a_193_47# _1006_/a_975_413# 0
C43325 _1006_/a_1059_315# _1006_/a_891_413# 0.31086f
C43326 _0179_ _0987_/a_27_47# 0
C43327 hold47/a_49_47# _1049_/a_27_47# 0
C43328 _0656_/a_59_75# _0656_/a_145_75# 0.00658f
C43329 _0247_ _0392_ 0
C43330 _1049_/a_466_413# _0186_ 0
C43331 _0476_ _0972_/a_93_21# 0.00134f
C43332 acc0.A\[1\] _1014_/a_466_413# 0
C43333 net182 _1055_/a_193_47# 0
C43334 net206 _0580_/a_109_47# 0.00119f
C43335 _0221_ _0725_/a_80_21# 0.07705f
C43336 _0343_ _0186_ 0.021f
C43337 _1052_/a_634_159# A[5] 0
C43338 _0984_/a_193_47# _0984_/a_891_413# 0.19683f
C43339 _0984_/a_27_47# _0984_/a_381_47# 0.06222f
C43340 _0984_/a_634_159# _0984_/a_1059_315# 0
C43341 net181 A[9] 0
C43342 net21 _1043_/a_466_413# 0
C43343 _0260_ clknet_0__0465_ 0
C43344 clknet_1_0__leaf__0462_ _0378_ 0.00631f
C43345 _0808_/a_266_47# _0808_/a_585_47# 0.0013f
C43346 _0817_/a_81_21# _0347_ 0
C43347 _1018_/a_592_47# clknet_1_0__leaf__0461_ 0
C43348 clkbuf_1_1__f__0461_/a_110_47# _0459_ 0.00377f
C43349 acc0.A\[19\] _0772_/a_79_21# 0
C43350 hold66/a_391_47# hold3/a_391_47# 0.00216f
C43351 net213 _0373_ 0
C43352 _0183_ net49 0.44042f
C43353 _0982_/a_891_413# _0117_ 0
C43354 _0181_ _0161_ 0
C43355 net9 net11 0.64124f
C43356 hold69/a_285_47# _0346_ 0.07685f
C43357 _0727_/a_193_47# _0332_ 0
C43358 _1039_/a_1059_315# VPWR 0.39794f
C43359 _0343_ hold19/a_49_47# 0.01595f
C43360 _0712_/a_297_297# _1031_/a_1059_315# 0
C43361 hold20/a_391_47# _0467_ 0
C43362 _0470_ _0163_ 0
C43363 _0986_/a_466_413# _0986_/a_381_47# 0.03733f
C43364 _0986_/a_193_47# _0986_/a_975_413# 0
C43365 _0986_/a_1059_315# _0986_/a_891_413# 0.31086f
C43366 _0524_/a_109_297# _0085_ 0
C43367 _0277_ _0219_ 0.00186f
C43368 _0856_/a_79_21# _0264_ 0.12885f
C43369 _1023_/a_634_159# _1023_/a_1017_47# 0
C43370 _1023_/a_466_413# _1023_/a_592_47# 0.00553f
C43371 _0990_/a_27_47# net47 0.02291f
C43372 _0400_ net6 0
C43373 hold101/a_391_47# _0432_ 0.00455f
C43374 _0277_ _0669_/a_111_297# 0
C43375 _0221_ _0128_ 0
C43376 _1042_/a_193_47# net128 0.00407f
C43377 _1042_/a_1059_315# _1042_/a_1017_47# 0
C43378 hold57/a_49_47# _0463_ 0
C43379 _0181_ _0158_ 0.27249f
C43380 _0313_ _0195_ 0
C43381 net36 hold59/a_285_47# 0.00124f
C43382 _0731_/a_299_297# clkbuf_0__0460_/a_110_47# 0
C43383 _0362_ _0317_ 0
C43384 _1045_/a_193_47# _0142_ 0
C43385 _1045_/a_1059_315# net20 0.01455f
C43386 _0459_ _0185_ 0.07363f
C43387 acc0.A\[5\] clknet_1_1__leaf__0464_ 0
C43388 _0346_ _0617_/a_68_297# 0.01742f
C43389 hold89/a_285_47# _0972_/a_93_21# 0
C43390 _0347_ _0084_ 0.05868f
C43391 _1036_/a_381_47# comp0.B\[4\] 0
C43392 _0466_ _1064_/a_381_47# 0
C43393 clknet_1_0__leaf__0464_ _0531_/a_27_297# 0
C43394 hold16/a_391_47# _1031_/a_193_47# 0.00283f
C43395 hold16/a_285_47# _1031_/a_634_159# 0.01163f
C43396 _0710_/a_109_297# _0216_ 0
C43397 net9 hold7/a_391_47# 0.01673f
C43398 _0404_ _0417_ 0
C43399 _0808_/a_585_47# _0345_ 0
C43400 _0752_/a_300_297# net51 0.00742f
C43401 hold77/a_49_47# _0219_ 0.00216f
C43402 pp[29] _1011_/a_891_413# 0
C43403 _0578_/a_27_297# _0369_ 0
C43404 _1057_/a_193_47# net192 0
C43405 _1056_/a_27_47# net47 0
C43406 _0981_/a_27_297# _0488_ 0.06252f
C43407 _0359_ _0319_ 0
C43408 net101 _1020_/a_193_47# 0
C43409 _0227_ _0755_/a_109_297# 0
C43410 _0997_/a_466_413# _0407_ 0
C43411 clknet_1_0__leaf__0458_ acc0.A\[9\] 0
C43412 _0732_/a_209_297# net93 0
C43413 _0732_/a_80_21# _0105_ 0.00479f
C43414 acc0.A\[4\] net12 0
C43415 _0425_ _0369_ 0
C43416 _0367_ _0352_ 0
C43417 net178 clkbuf_1_1__f__0458_/a_110_47# 0
C43418 _0743_/a_149_47# _0743_/a_240_47# 0.06872f
C43419 clknet_1_0__leaf__0462_ net112 0.15035f
C43420 _0858_/a_27_47# clknet_1_1__leaf__0457_ 0.20082f
C43421 _1002_/a_1059_315# net220 0
C43422 _0777_/a_47_47# _0394_ 0.38756f
C43423 _0777_/a_285_47# _0308_ 0.0012f
C43424 net58 clknet_1_1__leaf__0465_ 0.00371f
C43425 hold30/a_49_47# _0217_ 0.0675f
C43426 net34 _0481_ 0
C43427 clknet_1_0__leaf__0462_ acc0.A\[24\] 0.1222f
C43428 hold28/a_285_47# _0197_ 0.0054f
C43429 _0477_ _0164_ 0.03076f
C43430 _0216_ _0182_ 0.07322f
C43431 _0353_ _0219_ 0
C43432 _0227_ _0235_ 0
C43433 VPWR _0631_/a_109_297# 0.00717f
C43434 clkload4/a_268_47# VPWR 0
C43435 _0714_/a_51_297# net162 0.00141f
C43436 _1033_/a_27_47# _0565_/a_51_297# 0
C43437 _1057_/a_27_47# _0992_/a_1059_315# 0
C43438 _0743_/a_240_47# _0345_ 0
C43439 _0743_/a_51_297# _0219_ 0.17385f
C43440 _0294_ _0242_ 0.04254f
C43441 net215 pp[24] 0
C43442 hold30/a_391_47# net151 0
C43443 net63 net75 0.00346f
C43444 _0999_/a_975_413# _0218_ 0
C43445 _0445_ _0431_ 0
C43446 _0179_ _0191_ 0.35204f
C43447 _0195_ _1013_/a_634_159# 0.00722f
C43448 _0216_ _1013_/a_27_47# 0
C43449 _0636_/a_59_75# _0262_ 0
C43450 _0236_ _0749_/a_299_297# 0.0124f
C43451 _0249_ net51 0.0032f
C43452 _0728_/a_59_75# _0353_ 0
C43453 _0454_ _0264_ 0.02951f
C43454 input26/a_75_212# B[3] 0.19382f
C43455 _0995_/a_27_47# _0799_/a_80_21# 0.00129f
C43456 _1058_/a_975_413# acc0.A\[11\] 0
C43457 _0274_ _0086_ 0
C43458 _0984_/a_592_47# net77 0
C43459 acc0.A\[14\] _0181_ 0.23711f
C43460 net70 _0991_/a_592_47# 0
C43461 _0250_ _0105_ 0.0032f
C43462 _0130_ clkbuf_1_1__f__0463_/a_110_47# 0
C43463 _1000_/a_1059_315# net223 0
C43464 VPWR _1035_/a_561_413# 0.00345f
C43465 net139 _1052_/a_27_47# 0
C43466 _0172_ _1040_/a_27_47# 0.03606f
C43467 net30 _1040_/a_193_47# 0
C43468 _1001_/a_891_413# net45 0
C43469 _0217_ _0352_ 0.07525f
C43470 _1058_/a_27_47# VPWR 0.62822f
C43471 _0275_ _0271_ 0.00276f
C43472 _0298_ _0219_ 0.00791f
C43473 _0254_ _0433_ 0
C43474 _0754_/a_240_47# _0219_ 0.02773f
C43475 _0982_/a_381_47# _0181_ 0.01154f
C43476 _0814_/a_27_47# _0814_/a_109_47# 0.00517f
C43477 _0434_ acc0.A\[6\] 0.03751f
C43478 clknet_1_0__leaf__0465_ net20 0.00274f
C43479 comp0.B\[13\] _0141_ 0
C43480 _0992_/a_891_413# _0286_ 0
C43481 _0992_/a_381_47# _0283_ 0
C43482 _1056_/a_1059_315# pp[8] 0
C43483 hold38/a_391_47# _0477_ 0.0021f
C43484 _1055_/a_466_413# _0516_/a_27_297# 0
C43485 comp0.B\[7\] _0463_ 0
C43486 _1064_/a_193_47# _1064_/a_381_47# 0.10164f
C43487 _1064_/a_634_159# _1064_/a_891_413# 0.03684f
C43488 _1064_/a_27_47# _1064_/a_561_413# 0.00163f
C43489 _0643_/a_253_47# _0431_ 0
C43490 _1018_/a_466_413# net149 0
C43491 _0604_/a_113_47# _0373_ 0
C43492 _0180_ _0369_ 0
C43493 _1015_/a_27_47# net23 0.00981f
C43494 _1018_/a_891_413# _1017_/a_193_47# 0
C43495 output42/a_27_47# _0299_ 0
C43496 _0440_ _0987_/a_193_47# 0
C43497 _0472_ _0493_/a_27_47# 0
C43498 _0244_ _0771_/a_27_413# 0
C43499 _0111_ net99 0.00177f
C43500 _0712_/a_297_297# _0712_/a_561_47# 0
C43501 net9 clknet_1_1__leaf__0458_ 0.02783f
C43502 _1051_/a_466_413# net12 0
C43503 _1051_/a_193_47# _0194_ 0
C43504 _0343_ _1017_/a_193_47# 0.00194f
C43505 B[1] B[6] 0.00559f
C43506 _0845_/a_193_297# _0449_ 0
C43507 clknet_1_0__leaf__0458_ _0449_ 0
C43508 net1 _0585_/a_109_297# 0.00918f
C43509 comp0.B\[14\] hold6/a_49_47# 0
C43510 hold53/a_391_47# net111 0
C43511 clknet_1_1__leaf_clk clknet_1_0__leaf__0457_ 0.24619f
C43512 _0343_ _1060_/a_592_47# 0
C43513 net159 _1068_/a_975_413# 0
C43514 _0974_/a_222_93# _0166_ 0.00771f
C43515 _0266_ _0465_ 0.00461f
C43516 _0598_/a_79_21# _0374_ 0
C43517 control0.state\[0\] _0484_ 0.20427f
C43518 output35/a_27_47# VPWR 0.26464f
C43519 _0603_/a_68_297# _0373_ 0
C43520 _0348_ hold62/a_285_47# 0
C43521 clkbuf_0__0465_/a_110_47# _0084_ 0.00635f
C43522 _0343_ _0241_ 0.00484f
C43523 _1017_/a_27_47# acc0.A\[17\] 0
C43524 _0432_ _0369_ 0
C43525 net154 _0522_/a_109_47# 0
C43526 _0627_/a_109_93# clkbuf_1_1__f__0458_/a_110_47# 0
C43527 hold25/a_285_47# net8 0.07819f
C43528 _0713_/a_27_47# _0461_ 0.02171f
C43529 _1010_/a_1017_47# _0350_ 0
C43530 _0399_ _0087_ 0
C43531 acc0.A\[5\] _0825_/a_68_297# 0
C43532 _0737_/a_35_297# _0364_ 0.16656f
C43533 _0737_/a_285_47# _0360_ 0.00108f
C43534 _0737_/a_285_297# _0321_ 0.06416f
C43535 net58 _0452_ 0
C43536 hold16/a_285_47# _0345_ 0
C43537 _0330_ _0690_/a_68_297# 0
C43538 _0854_/a_79_21# _0854_/a_510_47# 0.00844f
C43539 _0854_/a_297_297# _0854_/a_215_47# 0
C43540 clknet_1_1__leaf__0464_ _1042_/a_634_159# 0
C43541 _0222_ net91 0
C43542 hold2/a_49_47# hold2/a_285_47# 0.22264f
C43543 hold74/a_391_47# net103 0
C43544 _0697_/a_300_47# _0322_ 0
C43545 _0697_/a_472_297# _0329_ 0
C43546 _0565_/a_240_47# _0208_ 0.02436f
C43547 _0289_ _0420_ 0.002f
C43548 hold74/a_49_47# _1016_/a_27_47# 0
C43549 _0768_/a_109_297# _0387_ 0
C43550 _0601_/a_150_297# clknet_1_0__leaf__0460_ 0
C43551 net234 clknet_1_0__leaf__0457_ 0
C43552 _0961_/a_199_47# clk 0
C43553 acc0.A\[7\] acc0.A\[6\] 0.00402f
C43554 net157 _1061_/a_1017_47# 0
C43555 _0479_ control0.count\[0\] 0.01924f
C43556 _0331_ _0329_ 0.16637f
C43557 _0217_ _0574_/a_109_297# 0.01154f
C43558 _0989_/a_1059_315# acc0.A\[6\] 0
C43559 clkbuf_1_1__f_clk/a_110_47# _1063_/a_27_47# 0.0025f
C43560 acc0.A\[31\] net41 0
C43561 _0697_/a_300_47# _0327_ 0
C43562 VPWR net239 0.25394f
C43563 hold36/a_49_47# net183 0
C43564 _0195_ net10 0.02741f
C43565 _0179_ _0812_/a_297_297# 0.00225f
C43566 _0312_ _0323_ 0.12162f
C43567 _0302_ clkbuf_0__0459_/a_110_47# 0.00153f
C43568 _0251_ _0829_/a_27_47# 0
C43569 clknet_1_0__leaf__0465_ _1052_/a_634_159# 0.002f
C43570 _0643_/a_103_199# clknet_0__0465_ 0.0033f
C43571 _0182_ net247 0.04023f
C43572 _0500_/a_27_47# _0534_/a_81_21# 0
C43573 input33/a_75_212# net33 0.10861f
C43574 B[8] net31 0.03568f
C43575 net46 clknet_1_0__leaf__0457_ 0.29313f
C43576 _1037_/a_1059_315# VPWR 0.40397f
C43577 net61 _0440_ 0
C43578 _0183_ _1016_/a_381_47# 0
C43579 _0700_/a_113_47# acc0.A\[28\] 0
C43580 comp0.B\[10\] _0140_ 0.0992f
C43581 net9 _1047_/a_27_47# 0
C43582 net7 _0205_ 0
C43583 _0255_ hold1/a_49_47# 0.05706f
C43584 net68 clknet_1_1__leaf__0457_ 0.00149f
C43585 hold30/a_391_47# _0378_ 0
C43586 _0121_ _0756_/a_285_47# 0
C43587 _0733_/a_544_297# _0324_ 0.00271f
C43588 _1041_/a_561_413# VPWR 0.0025f
C43589 hold98/a_49_47# A[13] 0
C43590 _0264_ _0846_/a_51_297# 0
C43591 net55 _0319_ 0
C43592 pp[15] _0995_/a_381_47# 0.00176f
C43593 net86 _0294_ 0.41617f
C43594 _0722_/a_510_47# _0351_ 0.00586f
C43595 _1005_/a_1017_47# _0103_ 0.00125f
C43596 _0157_ _0288_ 0
C43597 _0983_/a_193_47# clknet_1_0__leaf__0461_ 0
C43598 net17 _0565_/a_149_47# 0
C43599 _0260_ _0529_/a_109_47# 0
C43600 _0179_ _0512_/a_27_297# 0
C43601 hold24/a_49_47# net8 0.03827f
C43602 _0331_ _0221_ 0.07079f
C43603 _0438_ _0831_/a_285_297# 0.07766f
C43604 _0835_/a_78_199# _0465_ 0
C43605 clkbuf_1_1__f__0465_/a_110_47# _0428_ 0.01532f
C43606 clknet_1_1__leaf_clk _1062_/a_466_413# 0.03176f
C43607 _1018_/a_27_47# _0581_/a_27_297# 0
C43608 _0158_ _0507_/a_373_47# 0
C43609 _1060_/a_381_47# _0185_ 0
C43610 _0482_ _0975_/a_59_75# 0.00378f
C43611 _0401_ _0841_/a_79_21# 0
C43612 _1054_/a_891_413# clknet_1_1__leaf__0458_ 0.01349f
C43613 _1021_/a_193_47# clknet_1_1__leaf_clk 0
C43614 hold16/a_49_47# hold16/a_285_47# 0.22264f
C43615 _1002_/a_1059_315# net88 0
C43616 _1020_/a_193_47# _1020_/a_466_413# 0.07855f
C43617 _1020_/a_27_47# _1020_/a_1059_315# 0.04875f
C43618 _1002_/a_466_413# _0100_ 0.03705f
C43619 _0792_/a_80_21# _0406_ 0.15444f
C43620 net156 _0739_/a_79_21# 0
C43621 _1027_/a_1059_315# _0106_ 0
C43622 _1021_/a_975_413# net1 0
C43623 net70 clknet_1_0__leaf__0458_ 0.11374f
C43624 _1016_/a_27_47# _0583_/a_27_297# 0.00955f
C43625 net63 _0442_ 0.0946f
C43626 net45 hold19/a_391_47# 0
C43627 _0598_/a_79_21# _0752_/a_300_297# 0
C43628 _0248_ _0352_ 0
C43629 _0483_ clknet_1_0__leaf_clk 0.1738f
C43630 _0983_/a_27_47# _0265_ 0
C43631 _0983_/a_634_159# net47 0.01838f
C43632 _0341_ acc0.A\[30\] 0.10499f
C43633 _1016_/a_193_47# net43 0
C43634 _0209_ _0173_ 0
C43635 _0179_ clkbuf_1_0__f__0465_/a_110_47# 0
C43636 hold35/a_49_47# net179 0
C43637 _0183_ _0757_/a_68_297# 0.00107f
C43638 _1058_/a_466_413# clknet_1_1__leaf__0465_ 0.00178f
C43639 _0259_ _0785_/a_81_21# 0.1219f
C43640 _0217_ net207 0.00191f
C43641 _0180_ _1048_/a_634_159# 0.01784f
C43642 net22 hold5/a_49_47# 0
C43643 _0182_ _1048_/a_466_413# 0
C43644 _0998_/a_193_47# _1017_/a_193_47# 0.00148f
C43645 _0147_ _1047_/a_1059_315# 0
C43646 hold10/a_49_47# _0502_/a_27_47# 0.00441f
C43647 _1001_/a_1059_315# net46 0.13703f
C43648 acc0.A\[12\] _0189_ 0
C43649 _0346_ _0672_/a_215_47# 0.00178f
C43650 _0457_ _0584_/a_27_297# 0.00462f
C43651 net34 _0477_ 0.00126f
C43652 _1041_/a_634_159# _0550_/a_240_47# 0
C43653 _0443_ _0825_/a_68_297# 0
C43654 clknet_1_0__leaf__0461_ _0526_/a_27_47# 0.0029f
C43655 _1003_/a_634_159# _0466_ 0
C43656 _0222_ _0762_/a_510_47# 0
C43657 hold88/a_391_47# _0181_ 0
C43658 clkload4/a_268_47# clknet_1_0__leaf__0459_ 0.00208f
C43659 _0231_ net51 0.3599f
C43660 _1039_/a_27_47# _0494_/a_27_47# 0
C43661 net23 _0215_ 0
C43662 clkbuf_1_1__f_clk/a_110_47# _1062_/a_1059_315# 0.00957f
C43663 clknet_0__0458_ _0621_/a_285_297# 0
C43664 pp[8] VPWR 0.9631f
C43665 clknet_0__0459_ _0420_ 0
C43666 _0664_/a_79_21# VPWR 0.27259f
C43667 _0117_ clkbuf_0__0457_/a_110_47# 0.00913f
C43668 _0176_ _0540_/a_51_297# 0.00593f
C43669 _0924_/a_27_47# control0.reset 0
C43670 _1036_/a_193_47# net24 0
C43671 net121 control0.sh 0
C43672 _0098_ _0775_/a_79_21# 0.05031f
C43673 _1000_/a_381_47# _0393_ 0.00699f
C43674 net86 _0775_/a_297_297# 0
C43675 _0580_/a_27_297# _0350_ 0.05995f
C43676 _0413_ _0799_/a_303_47# 0
C43677 _0800_/a_240_47# _0411_ 0
C43678 clknet_0__0459_ _0459_ 0.01123f
C43679 _0343_ _0410_ 0.01749f
C43680 comp0.B\[12\] _1044_/a_891_413# 0.00349f
C43681 _1052_/a_1059_315# A[4] 0
C43682 _0269_ _0445_ 0
C43683 _0464_ _1061_/a_27_47# 0
C43684 _0924_/a_27_47# _1061_/a_891_413# 0.01004f
C43685 _0967_/a_403_297# control0.state\[2\] 0.00672f
C43686 _0486_ _0162_ 0
C43687 control0.count\[1\] clknet_1_0__leaf_clk 0.59945f
C43688 clknet_1_0__leaf__0462_ _0682_/a_150_297# 0
C43689 hold75/a_285_47# _0853_/a_68_297# 0
C43690 clkbuf_0__0459_/a_110_47# net6 0.24706f
C43691 _0343_ net62 0.0328f
C43692 hold57/a_391_47# _0176_ 0.04854f
C43693 _0606_/a_297_297# _0374_ 0
C43694 hold67/a_285_47# net143 0
C43695 _1000_/a_27_47# _0347_ 0.09692f
C43696 _1030_/a_975_413# _0336_ 0
C43697 _0414_ _0994_/a_891_413# 0
C43698 _0312_ net237 0.00371f
C43699 VPWR _1063_/a_27_47# 0.40523f
C43700 _1052_/a_891_413# net73 0
C43701 hold66/a_49_47# _0381_ 0
C43702 _0402_ _0651_/a_113_47# 0
C43703 _0762_/a_79_21# _0103_ 0.0506f
C43704 net97 net57 0
C43705 _1017_/a_381_47# clknet_1_1__leaf__0461_ 0
C43706 _0572_/a_27_297# net155 0.12696f
C43707 _0572_/a_109_47# net210 0
C43708 _0572_/a_109_297# _0195_ 0.02703f
C43709 acc0.A\[14\] _0507_/a_373_47# 0
C43710 clknet_1_1__leaf__0460_ hold9/a_49_47# 0
C43711 net179 A[9] 0.05743f
C43712 _0317_ _0324_ 0
C43713 acc0.A\[9\] _0288_ 0.01225f
C43714 VPWR _0974_/a_448_47# 0.0031f
C43715 _0647_/a_47_47# _0218_ 0
C43716 _0147_ _0186_ 0
C43717 clknet_1_1__leaf__0461_ _0158_ 0
C43718 _0993_/a_1017_47# net246 0
C43719 _0476_ net231 0
C43720 pp[7] _0369_ 0
C43721 _0182_ net100 0
C43722 net234 _0850_/a_68_297# 0
C43723 acc0.A\[26\] _0739_/a_79_21# 0.017f
C43724 _0655_/a_109_93# _0420_ 0.00158f
C43725 pp[8] output62/a_27_47# 0
C43726 _0443_ _0841_/a_79_21# 0.00645f
C43727 net59 _0342_ 0
C43728 clknet_1_0__leaf__0460_ _0377_ 0.01138f
C43729 _0172_ _1061_/a_466_413# 0
C43730 _0643_/a_253_47# _0269_ 0.0331f
C43731 _0579_/a_109_297# _0461_ 0.00422f
C43732 net185 comp0.B\[2\] 0
C43733 VPWR _1060_/a_27_47# 0.73635f
C43734 _1019_/a_27_47# acc0.A\[19\] 0
C43735 clkbuf_1_0__f__0459_/a_110_47# hold19/a_49_47# 0.02203f
C43736 acc0.A\[29\] clknet_1_1__leaf__0462_ 0.07971f
C43737 clkload3/Y _1017_/a_1059_315# 0
C43738 _0417_ _0419_ 0.13375f
C43739 _0714_/a_245_297# _0999_/a_193_47# 0
C43740 _0328_ _0693_/a_68_297# 0.00102f
C43741 clknet_1_0__leaf__0465_ A[8] 0
C43742 _0284_ _0289_ 0
C43743 net30 _0207_ 0
C43744 VPWR _0988_/a_891_413# 0.18681f
C43745 clknet_1_1__leaf__0460_ _1029_/a_27_47# 0
C43746 VPWR _0553_/a_245_297# 0.00576f
C43747 _1044_/a_27_47# _0542_/a_51_297# 0
C43748 A[11] acc0.A\[10\] 0
C43749 _0997_/a_1059_315# _0995_/a_27_47# 0
C43750 _0357_ VPWR 0.24276f
C43751 _1054_/a_193_47# _0186_ 0
C43752 net168 _1054_/a_561_413# 0
C43753 _0520_/a_27_297# net140 0
C43754 _0461_ _0399_ 0
C43755 _0174_ _1043_/a_27_47# 0.03652f
C43756 _1056_/a_381_47# _0186_ 0
C43757 net157 _1047_/a_193_47# 0.01582f
C43758 _0216_ _0616_/a_78_199# 0.01725f
C43759 _1023_/a_592_47# net177 0.00174f
C43760 _1023_/a_381_47# acc0.A\[23\] 0
C43761 hold89/a_285_47# _0975_/a_59_75# 0.00205f
C43762 _0699_/a_68_297# clknet_1_1__leaf__0462_ 0.00136f
C43763 pp[28] output57/a_27_47# 0.00173f
C43764 _0581_/a_109_297# _0242_ 0
C43765 _0094_ acc0.A\[13\] 0
C43766 hold45/a_49_47# hold45/a_285_47# 0.22264f
C43767 net238 net5 0.51011f
C43768 _0476_ hold38/a_285_47# 0.00183f
C43769 net118 net240 0
C43770 _0343_ _0227_ 0.00413f
C43771 _0704_/a_68_297# _0704_/a_150_297# 0.00477f
C43772 _0670_/a_79_21# _0670_/a_215_47# 0.04584f
C43773 _1044_/a_466_413# net20 0
C43774 hold64/a_391_47# acc0.A\[1\] 0
C43775 _0732_/a_80_21# _0359_ 0.04935f
C43776 clknet_1_0__leaf__0462_ net111 0.24413f
C43777 hold48/a_49_47# _1044_/a_1059_315# 0
C43778 pp[30] _0722_/a_215_47# 0
C43779 _0298_ _0799_/a_209_297# 0.065f
C43780 _0404_ _0799_/a_209_47# 0
C43781 _0299_ _0799_/a_80_21# 0.0023f
C43782 net205 clknet_1_1__leaf__0463_ 0.01628f
C43783 hold59/a_49_47# _0346_ 0
C43784 _0457_ _1015_/a_634_159# 0.00555f
C43785 net57 _0707_/a_201_297# 0.04639f
C43786 _0744_/a_27_47# acc0.A\[10\] 0.00411f
C43787 _0195_ _0707_/a_75_199# 0.00141f
C43788 _0329_ _1008_/a_27_47# 0
C43789 _0402_ _0806_/a_199_47# 0
C43790 _1037_/a_1017_47# control0.sh 0
C43791 acc0.A\[21\] _1068_/a_1059_315# 0
C43792 _0349_ hold62/a_391_47# 0
C43793 _0757_/a_150_297# _0379_ 0.00142f
C43794 _0380_ _0756_/a_285_47# 0.00131f
C43795 hold89/a_49_47# _0164_ 0
C43796 _0174_ _0171_ 0
C43797 _1037_/a_634_159# B[6] 0
C43798 hold27/a_391_47# net22 0
C43799 _1001_/a_891_413# VPWR 0.19189f
C43800 _0749_/a_384_47# _0350_ 0
C43801 net133 net9 0
C43802 net84 net221 0
C43803 net163 _1031_/a_561_413# 0
C43804 hold36/a_285_47# clknet_0__0464_ 0.01727f
C43805 net45 _1017_/a_466_413# 0.00447f
C43806 _0988_/a_27_47# pp[4] 0
C43807 VPWR _1062_/a_1059_315# 0.37695f
C43808 _0616_/a_292_297# _0240_ 0
C43809 _1059_/a_592_47# net229 0.00224f
C43810 _0157_ _0506_/a_299_297# 0
C43811 net145 _0506_/a_384_47# 0
C43812 _0780_/a_117_297# _0347_ 0
C43813 _0372_ _0326_ 0
C43814 _1039_/a_193_47# _0137_ 0.56479f
C43815 _1039_/a_891_413# net180 0
C43816 _1039_/a_466_413# _0172_ 0
C43817 _1021_/a_634_159# VPWR 0.18581f
C43818 net124 _1037_/a_27_47# 0.00136f
C43819 net43 net41 0.07759f
C43820 _0257_ _0255_ 0.58231f
C43821 _0170_ _0488_ 0
C43822 hold52/a_285_47# hold52/a_391_47# 0.41909f
C43823 acc0.A\[14\] clknet_1_1__leaf__0461_ 0
C43824 _0585_/a_27_297# _0526_/a_27_47# 0.01118f
C43825 _0574_/a_373_47# acc0.A\[24\] 0
C43826 _0359_ _0250_ 0.0092f
C43827 _0625_/a_59_75# _0433_ 0.04708f
C43828 _0503_/a_109_297# _0112_ 0
C43829 _0984_/a_27_47# clkbuf_1_0__f__0458_/a_110_47# 0.00913f
C43830 _0776_/a_27_47# _0308_ 0.04228f
C43831 _0776_/a_109_297# _0306_ 0
C43832 _0752_/a_27_413# net49 0
C43833 _0441_ clkbuf_1_0__f__0465_/a_110_47# 0.00149f
C43834 _0243_ _0719_/a_27_47# 0.00136f
C43835 net242 acc0.A\[29\] 0.12722f
C43836 _0332_ _0350_ 0.03904f
C43837 clknet_1_0__leaf__0463_ hold27/a_391_47# 0.00605f
C43838 net211 _0346_ 0.0187f
C43839 _0810_/a_113_47# _0296_ 0
C43840 _0606_/a_109_53# clkbuf_1_0__f__0460_/a_110_47# 0
C43841 _0100_ _0385_ 0
C43842 VPWR _0561_/a_240_47# 0.00493f
C43843 _1065_/a_1059_315# _1065_/a_891_413# 0.31086f
C43844 _1065_/a_193_47# _1065_/a_975_413# 0
C43845 _1065_/a_466_413# _1065_/a_381_47# 0.03733f
C43846 hold5/a_285_47# _0544_/a_51_297# 0
C43847 _0217_ _0237_ 0.0348f
C43848 hold85/a_391_47# clknet_1_1__leaf_clk 0.0011f
C43849 _0485_ _1066_/a_27_47# 0
C43850 _0817_/a_81_21# _0991_/a_1059_315# 0
C43851 _0998_/a_891_413# _0218_ 0.00207f
C43852 _1036_/a_1059_315# _1035_/a_466_413# 0.0042f
C43853 _1036_/a_891_413# _1035_/a_634_159# 0.00448f
C43854 _1036_/a_193_47# _1035_/a_381_47# 0
C43855 _0350_ _0685_/a_68_297# 0
C43856 control0.state\[1\] _0482_ 0
C43857 _0985_/a_1059_315# _0256_ 0
C43858 _0111_ acc0.A\[31\] 0.00333f
C43859 net225 net162 0
C43860 _0308_ _0219_ 0.26029f
C43861 B[1] comp0.B\[5\] 0
C43862 net31 _0548_/a_149_47# 0.00405f
C43863 comp0.B\[12\] _1042_/a_27_47# 0
C43864 comp0.B\[11\] _1042_/a_193_47# 0.17949f
C43865 _1014_/a_634_159# _1014_/a_466_413# 0.23992f
C43866 _1014_/a_193_47# _1014_/a_1059_315# 0.03405f
C43867 _1014_/a_27_47# _1014_/a_891_413# 0.03224f
C43868 _0851_/a_113_47# _0265_ 0
C43869 net33 hold84/a_391_47# 0.0128f
C43870 net228 hold82/a_49_47# 0.05864f
C43871 hold52/a_391_47# net52 0.01143f
C43872 VPWR _1047_/a_381_47# 0.07671f
C43873 VPWR _0472_ 1.16175f
C43874 _0181_ _0116_ 0
C43875 net56 _0729_/a_68_297# 0
C43876 clknet_1_0__leaf__0460_ net109 0
C43877 _1052_/a_193_47# _0149_ 0
C43878 hold101/a_49_47# net248 0
C43879 _0985_/a_27_47# _0458_ 0.02128f
C43880 net173 _0139_ 0
C43881 VPWR _1007_/a_592_47# 0.00114f
C43882 _0478_ _0484_ 0.05108f
C43883 _1021_/a_634_159# net48 0
C43884 _0734_/a_285_47# VPWR 0.00376f
C43885 hold87/a_285_47# _0217_ 0
C43886 VPWR _0850_/a_150_297# 0.00122f
C43887 _0171_ _0208_ 0.00564f
C43888 _1039_/a_193_47# comp0.B\[6\] 0
C43889 _0301_ _0345_ 0.0267f
C43890 pp[28] _0704_/a_68_297# 0
C43891 _0399_ _0465_ 0.00588f
C43892 net120 hold56/a_285_47# 0
C43893 _1055_/a_466_413# _0190_ 0
C43894 _1055_/a_891_413# net16 0.02171f
C43895 _0278_ net5 0.03803f
C43896 _0316_ _0317_ 0.55123f
C43897 clknet_1_1__leaf__0465_ _1060_/a_466_413# 0.00639f
C43898 pp[27] pp[28] 0.35321f
C43899 _0830_/a_79_21# _0989_/a_634_159# 0
C43900 _0830_/a_215_47# _0989_/a_27_47# 0
C43901 _0089_ _0841_/a_79_21# 0
C43902 input2/a_75_212# acc0.A\[11\] 0
C43903 _0235_ _0352_ 0
C43904 hold41/a_49_47# net2 0
C43905 clknet_1_1__leaf__0458_ _0840_/a_68_297# 0.00141f
C43906 clkbuf_1_0__f__0459_/a_110_47# _1017_/a_193_47# 0
C43907 _0956_/a_114_297# comp0.B\[0\] 0.01151f
C43908 _1018_/a_1059_315# net103 0.00119f
C43909 net66 acc0.A\[10\] 0.03446f
C43910 pp[15] _0219_ 0
C43911 _0664_/a_79_21# _0283_ 0.01006f
C43912 _0335_ _0334_ 0.24888f
C43913 net112 _1025_/a_891_413# 0
C43914 _1026_/a_193_47# acc0.A\[25\] 0.09716f
C43915 net1 _0178_ 0.00188f
C43916 hold78/a_49_47# hold78/a_391_47# 0.00188f
C43917 _0390_ _1001_/a_891_413# 0
C43918 _0819_/a_81_21# _0819_/a_299_297# 0.08213f
C43919 _0317_ _0347_ 0
C43920 acc0.A\[5\] net148 0.00367f
C43921 _0149_ net12 0.21214f
C43922 _1002_/a_1017_47# _0369_ 0
C43923 net55 _0333_ 0.00685f
C43924 VPWR _0586_/a_27_47# 0.23104f
C43925 VPWR _0748_/a_384_47# 0.00139f
C43926 _0210_ _0496_/a_27_47# 0
C43927 _0376_ _0227_ 0.28528f
C43928 _0585_/a_109_297# control0.sh 0
C43929 _0716_/a_27_47# _0347_ 0.39639f
C43930 _1025_/a_891_413# acc0.A\[24\] 0
C43931 _0183_ _1059_/a_193_47# 0
C43932 comp0.B\[1\] comp0.B\[0\] 0.31214f
C43933 net53 _0574_/a_27_297# 0
C43934 net165 _0347_ 0.0262f
C43935 hold41/a_285_47# net3 0
C43936 _0305_ _0370_ 0
C43937 _0107_ _0318_ 0
C43938 control0.state\[1\] _0476_ 0.24544f
C43939 net120 _1032_/a_193_47# 0
C43940 _0985_/a_561_413# net61 0
C43941 hold49/a_391_47# VPWR 0.21276f
C43942 clknet_1_0__leaf__0459_ _1060_/a_27_47# 0.00263f
C43943 _0284_ _0418_ 0
C43944 comp0.B\[7\] clkbuf_1_0__f__0463_/a_110_47# 0.03767f
C43945 _0216_ _0704_/a_150_297# 0
C43946 _1042_/a_193_47# _0202_ 0
C43947 _0836_/a_68_297# _0836_/a_150_297# 0.00477f
C43948 _0222_ _1022_/a_891_413# 0.05384f
C43949 VPWR hold19/a_391_47# 0.18038f
C43950 _1037_/a_193_47# _1036_/a_466_413# 0
C43951 _1037_/a_27_47# _1036_/a_1059_315# 0
C43952 _1037_/a_466_413# _1036_/a_193_47# 0
C43953 _0481_ _1070_/a_466_413# 0
C43954 _0963_/a_35_297# VPWR 0.19366f
C43955 clknet_1_1__leaf__0464_ net128 0.12605f
C43956 output59/a_27_47# net59 0.16913f
C43957 _0273_ _0828_/a_113_297# 0
C43958 _0836_/a_68_297# _0437_ 0
C43959 _0531_/a_27_297# clkbuf_1_0__f__0464_/a_110_47# 0
C43960 clkbuf_0__0463_/a_110_47# clknet_1_1__leaf__0457_ 0.00168f
C43961 _0817_/a_81_21# _0425_ 0.14266f
C43962 _0817_/a_266_47# _0423_ 0.00431f
C43963 _0300_ _0668_/a_79_21# 0.11183f
C43964 _0297_ _0668_/a_297_47# 0.10967f
C43965 _0225_ net51 0.0678f
C43966 _0999_/a_1059_315# _0352_ 0
C43967 _0983_/a_193_47# _0218_ 0
C43968 hold78/a_391_47# _0129_ 0
C43969 _0255_ net11 0
C43970 _1013_/a_193_47# pp[31] 0
C43971 _0596_/a_59_75# _0596_/a_145_75# 0.00658f
C43972 net212 _0437_ 0.16657f
C43973 _0429_ _0827_/a_109_297# 0
C43974 clknet_0__0458_ net77 0
C43975 _0781_/a_68_297# _0781_/a_150_297# 0.00477f
C43976 _0640_/a_392_297# _0255_ 0.00267f
C43977 _0820_/a_297_297# _0428_ 0.00282f
C43978 _0467_ hold56/a_391_47# 0
C43979 comp0.B\[2\] _1033_/a_634_159# 0.01672f
C43980 _0422_ _0181_ 0
C43981 _0195_ _0146_ 0.00195f
C43982 _0680_/a_80_21# _0392_ 0
C43983 _0217_ _1005_/a_27_47# 0
C43984 net150 _1005_/a_193_47# 0.04053f
C43985 net190 _1028_/a_634_159# 0.04875f
C43986 _0195_ _1014_/a_891_413# 0
C43987 _0216_ _1014_/a_466_413# 0
C43988 acc0.A\[10\] _0350_ 0
C43989 _1038_/a_1059_315# comp0.B\[10\] 0
C43990 _0287_ _0218_ 0
C43991 _0293_ _0294_ 0.01781f
C43992 _0350_ _0738_/a_68_297# 0.17183f
C43993 output67/a_27_47# _1057_/a_634_159# 0
C43994 _0992_/a_193_47# _0417_ 0
C43995 _0845_/a_109_47# _0447_ 0.05914f
C43996 hold33/a_391_47# _0176_ 0
C43997 _0274_ _0350_ 0.00167f
C43998 comp0.B\[13\] _1043_/a_27_47# 0
C43999 _0576_/a_27_297# net177 0
C44000 _0972_/a_256_47# _0468_ 0.00146f
C44001 _1003_/a_193_47# clknet_1_0__leaf__0460_ 0.04147f
C44002 net34 hold89/a_49_47# 0.00181f
C44003 clkbuf_0__0462_/a_110_47# hold90/a_285_47# 0.01903f
C44004 control0.state\[0\] hold89/a_391_47# 0.00224f
C44005 control0.state\[1\] hold89/a_285_47# 0.05177f
C44006 _1059_/a_193_47# acc0.A\[15\] 0.00819f
C44007 _1001_/a_891_413# clknet_1_0__leaf__0459_ 0
C44008 _1019_/a_27_47# net1 0
C44009 _0279_ clknet_1_1__leaf__0459_ 0.54857f
C44010 _0643_/a_103_199# _0986_/a_27_47# 0
C44011 clknet_1_1__leaf_clk _0160_ 0.11716f
C44012 _1018_/a_27_47# _0116_ 0.09897f
C44013 _1018_/a_466_413# net206 0.01413f
C44014 _1018_/a_891_413# net219 0.00274f
C44015 _1008_/a_634_159# _1008_/a_381_47# 0
C44016 _1055_/a_27_47# _1055_/a_193_47# 0.97064f
C44017 input21/a_75_212# _0203_ 0
C44018 _0425_ _0084_ 0
C44019 _0488_ _1069_/a_1017_47# 0
C44020 hold56/a_391_47# comp0.B\[0\] 0
C44021 _0648_/a_109_297# VPWR 0.00219f
C44022 _0129_ net163 0
C44023 _1020_/a_193_47# _0118_ 0.41149f
C44024 _1020_/a_891_413# _1020_/a_1017_47# 0.00617f
C44025 net53 _1025_/a_634_159# 0.00859f
C44026 output53/a_27_47# _1025_/a_891_413# 0
C44027 _0231_ _0324_ 0
C44028 _0791_/a_113_297# _0791_/a_199_47# 0
C44029 _1035_/a_891_413# comp0.B\[5\] 0.00833f
C44030 _1035_/a_561_413# comp0.B\[3\] 0
C44031 _0343_ net219 0.24322f
C44032 A[11] _0188_ 0.01638f
C44033 _1016_/a_27_47# _0114_ 0.00633f
C44034 _0226_ _0234_ 0.00137f
C44035 _0255_ hold7/a_391_47# 0
C44036 pp[30] net57 0
C44037 _0390_ _0586_/a_27_47# 0
C44038 net69 net47 0.04441f
C44039 clknet_0__0458_ _0986_/a_1059_315# 0.00214f
C44040 hold69/a_49_47# _0748_/a_81_21# 0
C44041 clknet_0__0457_ _1014_/a_1059_315# 0
C44042 _0515_/a_299_297# net181 0.05857f
C44043 clknet_0__0463_ _0533_/a_27_297# 0
C44044 _0346_ _0669_/a_29_53# 0
C44045 _0104_ _0249_ 0
C44046 _0180_ net134 0.00275f
C44047 _1054_/a_466_413# _0518_/a_27_297# 0.00138f
C44048 net84 _1017_/a_27_47# 0
C44049 _0388_ _0766_/a_109_297# 0.00279f
C44050 pp[8] net182 0
C44051 net160 clknet_1_1__leaf__0463_ 0.00144f
C44052 _1032_/a_634_159# comp0.B\[0\] 0
C44053 _1041_/a_381_47# _0172_ 0
C44054 VPWR B[4] 0.27076f
C44055 _0997_/a_634_159# _0345_ 0.00212f
C44056 net89 _0466_ 0
C44057 _1004_/a_193_47# _0758_/a_79_21# 0.00204f
C44058 _0462_ _1007_/a_1059_315# 0
C44059 pp[28] _0216_ 0.00239f
C44060 _0846_/a_245_297# _0449_ 0.00109f
C44061 _0992_/a_381_47# _0345_ 0
C44062 acc0.A\[1\] clkbuf_1_1__f__0457_/a_110_47# 0.21162f
C44063 clknet_1_1__leaf__0457_ hold71/a_49_47# 0.00999f
C44064 _0410_ _0793_/a_51_297# 0
C44065 hold94/a_49_47# net241 0.00238f
C44066 hold94/a_285_47# _0377_ 0.01545f
C44067 _0227_ _0224_ 0
C44068 A[7] net11 0
C44069 _0991_/a_891_413# acc0.A\[15\] 0
C44070 net197 _0347_ 0.06729f
C44071 _0984_/a_466_413# _0184_ 0
C44072 _0826_/a_219_297# _0434_ 0.12012f
C44073 _0837_/a_81_21# acc0.A\[5\] 0.00136f
C44074 clknet_1_0__leaf__0462_ _0375_ 0
C44075 _0506_/a_81_21# _0505_/a_27_297# 0
C44076 _0982_/a_634_159# net234 0
C44077 net45 _0393_ 0.02614f
C44078 _0578_/a_109_297# _0183_ 0.00717f
C44079 hold65/a_49_47# clknet_1_0__leaf__0465_ 0
C44080 _0117_ _0350_ 0.00903f
C44081 _0578_/a_373_47# _0217_ 0
C44082 _0404_ _0668_/a_79_21# 0
C44083 _0458_ _0197_ 0.00337f
C44084 pp[9] hold35/a_285_47# 0
C44085 _0218_ _0793_/a_240_47# 0
C44086 _0280_ hold81/a_49_47# 0
C44087 _0179_ _1059_/a_193_47# 0.00565f
C44088 hold26/a_49_47# net174 0
C44089 _1000_/a_975_413# _0352_ 0
C44090 _0701_/a_209_47# _0350_ 0
C44091 _0399_ _0582_/a_27_297# 0
C44092 _0111_ net43 0
C44093 net155 _0124_ 0.01872f
C44094 _0902_/a_27_47# clknet_1_0__leaf__0457_ 0.24127f
C44095 _1016_/a_634_159# clknet_1_1__leaf__0461_ 0.04434f
C44096 VPWR net149 1.41937f
C44097 _0679_/a_150_297# _0240_ 0
C44098 pp[19] pp[23] 0.17884f
C44099 VPWR _1017_/a_466_413# 0.24085f
C44100 _0679_/a_150_297# _0369_ 0
C44101 _0432_ _0084_ 0
C44102 _1037_/a_634_159# comp0.B\[5\] 0
C44103 _0416_ clknet_1_1__leaf__0459_ 0.00327f
C44104 clknet_1_1__leaf__0460_ _0745_/a_193_47# 0
C44105 _0183_ net202 0
C44106 net70 _0506_/a_299_297# 0
C44107 _0370_ _0181_ 0.00355f
C44108 _0563_/a_51_297# _0563_/a_512_297# 0.0116f
C44109 _0548_/a_149_47# _0548_/a_240_47# 0.06872f
C44110 _1057_/a_27_47# _0186_ 0
C44111 _1015_/a_466_413# net149 0
C44112 _0183_ clknet_1_1__leaf__0463_ 0
C44113 acc0.A\[29\] hold80/a_49_47# 0.01371f
C44114 _0804_/a_297_297# VPWR 0.01592f
C44115 _1056_/a_1059_315# A[10] 0
C44116 _1017_/a_193_47# clkbuf_0__0461_/a_110_47# 0
C44117 _0255_ clknet_1_1__leaf__0458_ 0.25651f
C44118 VPWR _1033_/a_27_47# 0.45498f
C44119 _1044_/a_193_47# net19 0
C44120 _0243_ _0614_/a_29_53# 0.25566f
C44121 clknet_1_0__leaf__0465_ _1049_/a_27_47# 0.0035f
C44122 _0732_/a_80_21# _0325_ 0
C44123 _0143_ _0464_ 0.00156f
C44124 acc0.A\[8\] _0181_ 0.1815f
C44125 VPWR _1050_/a_1059_315# 0.39779f
C44126 clknet_1_0__leaf__0459_ hold19/a_391_47# 0.04109f
C44127 clknet_0_clk net159 0.35498f
C44128 _0511_/a_81_21# net192 0.06452f
C44129 comp0.B\[10\] net129 0
C44130 hold45/a_285_47# _0156_ 0.00225f
C44131 _1010_/a_27_47# _1010_/a_1059_315# 0.04875f
C44132 _1010_/a_193_47# _1010_/a_466_413# 0.07482f
C44133 clknet_1_0__leaf__0462_ _1004_/a_193_47# 0.0109f
C44134 _0644_/a_285_47# net42 0.0793f
C44135 _0644_/a_129_47# acc0.A\[15\] 0.00228f
C44136 _0717_/a_80_21# net57 0.00106f
C44137 _0991_/a_193_47# _0181_ 0.04013f
C44138 _0682_/a_68_297# _1025_/a_381_47# 0
C44139 pp[27] _1010_/a_975_413# 0
C44140 _1040_/a_27_47# _1040_/a_193_47# 0.96163f
C44141 _0462_ clkbuf_1_0__f__0462_/a_110_47# 0.00359f
C44142 _0322_ _0318_ 0.29911f
C44143 clkbuf_0__0462_/a_110_47# clknet_0__0462_ 1.69329f
C44144 acc0.A\[14\] clkbuf_1_1__f__0459_/a_110_47# 0.00222f
C44145 _0598_/a_79_21# _0225_ 0
C44146 net57 _0339_ 0.13706f
C44147 _0146_ _1048_/a_193_47# 0.57727f
C44148 _0198_ _1048_/a_1059_315# 0.00602f
C44149 _0195_ _0338_ 0
C44150 _0536_/a_240_47# net157 0.05803f
C44151 _0327_ _0318_ 0.20922f
C44152 _1002_/a_27_47# _0183_ 0.02489f
C44153 _1002_/a_634_159# _0217_ 0.0202f
C44154 _0590_/a_113_47# _0122_ 0
C44155 _0325_ _0250_ 0
C44156 hold54/a_49_47# _0181_ 0.00227f
C44157 _0196_ _0142_ 0
C44158 _1020_/a_891_413# _0461_ 0.00121f
C44159 _1067_/a_27_47# _1067_/a_193_47# 0.96675f
C44160 _0397_ _0352_ 0.04668f
C44161 _0174_ _0550_/a_149_47# 0.0224f
C44162 net191 hold50/a_391_47# 0
C44163 _0343_ _0352_ 0.46548f
C44164 clkbuf_0__0458_/a_110_47# _0445_ 0.00584f
C44165 _0112_ _0526_/a_27_47# 0
C44166 net56 net239 0
C44167 _1009_/a_634_159# _1009_/a_1059_315# 0
C44168 _1009_/a_27_47# _1009_/a_381_47# 0.06222f
C44169 _1009_/a_193_47# _1009_/a_891_413# 0.19497f
C44170 _0330_ net114 0
C44171 _0833_/a_79_21# clknet_1_1__leaf__0465_ 0
C44172 _0645_/a_285_47# _1059_/a_27_47# 0
C44173 clknet_1_0__leaf__0460_ hold93/a_391_47# 0.01447f
C44174 hold100/a_391_47# VPWR 0.18146f
C44175 _0238_ clkbuf_1_0__f__0460_/a_110_47# 0.01305f
C44176 comp0.B\[15\] _0565_/a_51_297# 0.00597f
C44177 hold5/a_391_47# net18 0
C44178 _1065_/a_466_413# control0.reset 0
C44179 acc0.A\[12\] net67 0.05934f
C44180 _0982_/a_466_413# VPWR 0.2527f
C44181 _0476_ _1066_/a_634_159# 0.00426f
C44182 _0399_ _0831_/a_117_297# 0.00325f
C44183 _0446_ _0842_/a_145_75# 0
C44184 _0450_ _0842_/a_59_75# 0.00479f
C44185 _0817_/a_266_297# _0089_ 0
C44186 _1036_/a_891_413# net121 0.00613f
C44187 _1036_/a_1059_315# _0133_ 0
C44188 comp0.B\[4\] _1035_/a_193_47# 0.00199f
C44189 _0602_/a_113_47# acc0.A\[23\] 0
C44190 _0186_ acc0.A\[6\] 0.73915f
C44191 net111 _1025_/a_891_413# 0
C44192 net14 net13 0.27221f
C44193 _1036_/a_592_47# B[15] 0
C44194 _0238_ _0250_ 0
C44195 _0967_/a_487_297# net1 0
C44196 clkbuf_1_1__f__0461_/a_110_47# _0347_ 0.01417f
C44197 net8 acc0.A\[15\] 0
C44198 acc0.A\[27\] _1027_/a_193_47# 0.00111f
C44199 _1032_/a_193_47# net118 0.01393f
C44200 hold79/a_391_47# _0168_ 0.0255f
C44201 _0557_/a_245_297# _0211_ 0
C44202 _0643_/a_253_47# clkbuf_0__0458_/a_110_47# 0
C44203 _1018_/a_1059_315# _0774_/a_68_297# 0.00159f
C44204 _1071_/a_193_47# _1071_/a_592_47# 0
C44205 _1071_/a_466_413# _1071_/a_561_413# 0.00772f
C44206 _1071_/a_634_159# _1071_/a_975_413# 0
C44207 _0254_ _0399_ 0.08732f
C44208 _1014_/a_466_413# net100 0.00793f
C44209 _0996_/a_193_47# _0410_ 0.00242f
C44210 _0996_/a_634_159# net238 0.03192f
C44211 _1015_/a_561_413# _0208_ 0.00173f
C44212 net64 _0181_ 0
C44213 _1000_/a_193_47# clkbuf_1_0__f__0461_/a_110_47# 0.00156f
C44214 B[13] B[11] 0.04134f
C44215 _0235_ _0237_ 0
C44216 hold14/a_285_47# net29 0
C44217 _0558_/a_68_297# _1036_/a_1059_315# 0
C44218 _0426_ _0347_ 0.11251f
C44219 _1013_/a_466_413# net42 0
C44220 net45 _0714_/a_51_297# 0.00681f
C44221 hold10/a_49_47# hold10/a_391_47# 0.00188f
C44222 _0177_ _0175_ 0
C44223 net61 net175 0
C44224 hold53/a_391_47# VPWR 0.18699f
C44225 _0821_/a_113_47# _0437_ 0
C44226 _1035_/a_1059_315# net26 0
C44227 _0423_ _0181_ 0.01155f
C44228 _0836_/a_68_297# _0252_ 0
C44229 net46 _0246_ 0
C44230 _0195_ _1026_/a_27_47# 0
C44231 VPWR _0094_ 0.59841f
C44232 net157 _1046_/a_27_47# 0.00739f
C44233 _0689_/a_68_297# _0737_/a_35_297# 0.00115f
C44234 net179 _0190_ 0.00385f
C44235 clknet_1_1__leaf__0465_ _0158_ 0.2017f
C44236 _0252_ net212 0
C44237 net65 _0087_ 0.07561f
C44238 _0809_/a_384_47# _0345_ 0
C44239 _0437_ _0989_/a_891_413# 0
C44240 _0087_ _0989_/a_466_413# 0
C44241 _0195_ net99 0.00111f
C44242 acc0.A\[24\] _1006_/a_27_47# 0
C44243 _0178_ control0.sh 0.22375f
C44244 net45 net206 0.05917f
C44245 clknet_1_0__leaf__0460_ control0.reset 0
C44246 _1015_/a_381_47# net17 0
C44247 _1020_/a_27_47# acc0.A\[20\] 0.00426f
C44248 _0186_ _0523_/a_384_47# 0
C44249 net168 _0150_ 0
C44250 VPWR A[10] 0.23516f
C44251 net130 _0194_ 0
C44252 net36 _1039_/a_561_413# 0.00218f
C44253 _0330_ _0365_ 0
C44254 _0317_ _0106_ 0
C44255 input25/a_75_212# _0175_ 0.00193f
C44256 net88 _1067_/a_561_413# 0
C44257 _1002_/a_466_413# control0.add 0
C44258 _0195_ _1048_/a_381_47# 0
C44259 _0389_ net223 0
C44260 _1012_/a_381_47# _0352_ 0.00187f
C44261 clknet_1_0__leaf__0459_ net149 0.00132f
C44262 _0328_ _0743_/a_51_297# 0
C44263 output65/a_27_47# A[8] 0
C44264 _0343_ _1016_/a_975_413# 0
C44265 _0984_/a_27_47# acc0.A\[15\] 0.01076f
C44266 clknet_1_0__leaf__0459_ _1017_/a_466_413# 0.00141f
C44267 clknet_1_0__leaf__0462_ net199 0.04642f
C44268 net221 acc0.A\[18\] 0
C44269 _0217_ _0222_ 0.01813f
C44270 hold36/a_285_47# comp0.B\[14\] 0.0886f
C44271 _1069_/a_27_47# _1069_/a_634_159# 0.13646f
C44272 net3 net4 0.05745f
C44273 net162 _0340_ 0.09777f
C44274 _0490_ net167 0.54952f
C44275 _0786_/a_80_21# _0295_ 0.14328f
C44276 _0555_/a_51_297# control0.sh 0.00351f
C44277 _0225_ _0606_/a_297_297# 0
C44278 _0481_ _0168_ 0.24728f
C44279 _0714_/a_51_297# _0587_/a_27_47# 0
C44280 _0135_ _1036_/a_193_47# 0
C44281 hold20/a_391_47# _0483_ 0.00716f
C44282 _0998_/a_1059_315# _0347_ 0
C44283 net15 net9 0
C44284 _0313_ acc0.A\[26\] 0.20896f
C44285 net69 _0848_/a_109_297# 0
C44286 acc0.A\[27\] _1026_/a_1059_315# 0
C44287 comp0.B\[7\] hold25/a_285_47# 0
C44288 _0512_/a_109_297# acc0.A\[11\] 0.0015f
C44289 _0405_ acc0.A\[13\] 0
C44290 _1030_/a_193_47# hold62/a_391_47# 0.00283f
C44291 _1030_/a_634_159# hold62/a_285_47# 0.01163f
C44292 net69 _0294_ 0
C44293 VPWR _0508_/a_299_297# 0.21113f
C44294 _0985_/a_634_159# _0350_ 0
C44295 B[14] net32 0
C44296 _0486_ _0969_/a_109_297# 0.00531f
C44297 net247 net7 0.08822f
C44298 net22 net152 0.06106f
C44299 input22/a_75_212# _0139_ 0
C44300 _0376_ _0352_ 0.02139f
C44301 _0084_ _0986_/a_381_47# 0.12804f
C44302 _0579_/a_109_47# _0457_ 0
C44303 _1018_/a_193_47# _0350_ 0
C44304 hold96/a_285_47# _1024_/a_466_413# 0
C44305 hold96/a_49_47# _1024_/a_1059_315# 0
C44306 _1053_/a_1059_315# net9 0
C44307 _1038_/a_975_413# _0136_ 0
C44308 comp0.B\[2\] net119 0.03951f
C44309 net239 _0345_ 0
C44310 _0891_/a_27_47# _0461_ 0.11003f
C44311 net190 net114 0.06896f
C44312 _0453_ net149 0
C44313 _0462_ _0772_/a_79_21# 0
C44314 _0624_/a_59_75# _0186_ 0
C44315 clknet_1_1__leaf__0462_ _1008_/a_1059_315# 0.0035f
C44316 _1032_/a_1059_315# _0565_/a_149_47# 0
C44317 comp0.B\[3\] _0561_/a_240_47# 0
C44318 _0449_ _0448_ 0.08694f
C44319 VPWR _1046_/a_891_413# 0.17804f
C44320 _1022_/a_634_159# _1022_/a_381_47# 0
C44321 input2/a_75_212# A[12] 0
C44322 _0486_ _0950_/a_75_212# 0
C44323 _0178_ net157 0.05815f
C44324 acc0.A\[14\] clknet_1_1__leaf__0465_ 0.00608f
C44325 hold49/a_285_47# _0172_ 0.06117f
C44326 _0856_/a_215_47# acc0.A\[0\] 0
C44327 _1052_/a_466_413# _0525_/a_299_297# 0
C44328 VPWR _0393_ 0.93114f
C44329 clknet_1_0__leaf__0463_ net152 0
C44330 _0994_/a_27_47# _0994_/a_193_47# 0.97386f
C44331 _0607_/a_27_297# _0307_ 0
C44332 _0357_ net56 0.01572f
C44333 _0275_ _0986_/a_193_47# 0.47267f
C44334 _0272_ _0986_/a_466_413# 0
C44335 _0473_ comp0.B\[5\] 0.04371f
C44336 net211 _1001_/a_634_159# 0.02165f
C44337 _0217_ net220 0
C44338 _0289_ _0812_/a_79_21# 0
C44339 _0292_ _0812_/a_297_297# 0
C44340 _1008_/a_381_47# net94 0
C44341 clkbuf_0_clk/a_110_47# _0466_ 0.00825f
C44342 _1055_/a_466_413# _1055_/a_592_47# 0.00553f
C44343 _1055_/a_634_159# _1055_/a_1017_47# 0
C44344 _0313_ _0733_/a_222_93# 0
C44345 _0505_/a_27_297# _0184_ 0.11879f
C44346 hold43/a_285_47# hold43/a_391_47# 0.41909f
C44347 net36 _0262_ 0
C44348 _0718_/a_47_47# net57 0
C44349 hold24/a_49_47# comp0.B\[7\] 0.29604f
C44350 _0984_/a_27_47# _0179_ 0.00212f
C44351 VPWR _0758_/a_79_21# 0.50341f
C44352 _0608_/a_109_297# _0608_/a_27_47# 0
C44353 _1054_/a_1059_315# net63 0
C44354 hold14/a_49_47# _1036_/a_1059_315# 0
C44355 hold14/a_391_47# _1036_/a_634_159# 0
C44356 hold14/a_285_47# _1036_/a_466_413# 0.0041f
C44357 _1003_/a_634_159# _1003_/a_975_413# 0
C44358 _1003_/a_466_413# _1003_/a_561_413# 0.00772f
C44359 _0218_ _0840_/a_68_297# 0.17489f
C44360 net82 _0399_ 0
C44361 hold59/a_49_47# net221 0
C44362 _0456_ _1019_/a_193_47# 0
C44363 _1036_/a_27_47# B[4] 0
C44364 _0248_ _0763_/a_193_47# 0.00411f
C44365 _0372_ _0763_/a_109_47# 0
C44366 hold64/a_391_47# _0216_ 0.05333f
C44367 hold45/a_49_47# _1058_/a_27_47# 0
C44368 _0207_ _1040_/a_27_47# 0
C44369 net171 _1040_/a_193_47# 0
C44370 _0287_ net228 0.03225f
C44371 comp0.B\[11\] clknet_1_1__leaf__0464_ 0.10617f
C44372 acc0.A\[20\] _0219_ 0
C44373 VPWR _0484_ 0.31985f
C44374 hold33/a_285_47# _0548_/a_51_297# 0
C44375 clknet_0__0463_ _0199_ 0.00222f
C44376 _0212_ _0955_/a_304_297# 0
C44377 net138 _0180_ 0
C44378 hold58/a_285_47# net205 0.01149f
C44379 _0176_ net195 0.02349f
C44380 input7/a_75_212# A[15] 0.2006f
C44381 hold20/a_49_47# clknet_0_clk 0
C44382 net22 _1042_/a_466_413# 0
C44383 _1054_/a_891_413# net15 0.00384f
C44384 net169 _0518_/a_27_297# 0
C44385 _1054_/a_466_413# _0191_ 0.00148f
C44386 _0825_/a_68_297# _0825_/a_150_297# 0.00477f
C44387 _0525_/a_299_297# _0194_ 0.00955f
C44388 _0830_/a_215_47# clknet_1_1__leaf__0458_ 0
C44389 _0343_ _0613_/a_109_297# 0.00243f
C44390 _0257_ _0989_/a_27_47# 0
C44391 _0997_/a_592_47# _0219_ 0.00124f
C44392 _0174_ _0494_/a_27_47# 0.15457f
C44393 _0195_ _0396_ 0
C44394 _0844_/a_382_297# _0844_/a_297_47# 0
C44395 _1004_/a_634_159# _0102_ 0.0515f
C44396 _1004_/a_466_413# _0352_ 0.00387f
C44397 _1004_/a_381_47# _0347_ 0
C44398 clkbuf_1_1__f__0462_/a_110_47# acc0.A\[28\] 0.00642f
C44399 net190 _0365_ 0
C44400 net197 _0106_ 0.00165f
C44401 _0983_/a_27_47# _0347_ 0.03354f
C44402 net23 _1065_/a_193_47# 0.01791f
C44403 _0362_ _0462_ 0
C44404 VPWR _0256_ 0.62159f
C44405 _0506_/a_81_21# _0184_ 0.17506f
C44406 _0179_ net10 0.03001f
C44407 net236 clkbuf_0_clk/a_110_47# 0.00262f
C44408 _0765_/a_79_21# hold73/a_285_47# 0
C44409 _0982_/a_1017_47# _0456_ 0
C44410 net68 net234 0
C44411 _0195_ _0580_/a_27_297# 0.02223f
C44412 B[14] net10 0.01324f
C44413 _0664_/a_79_21# _0345_ 0.01021f
C44414 net90 _1024_/a_1059_315# 0
C44415 _0229_ VPWR 1.09471f
C44416 VPWR _0987_/a_1059_315# 0.4152f
C44417 _1024_/a_27_47# _1024_/a_466_413# 0.27314f
C44418 _1024_/a_193_47# _1024_/a_634_159# 0.12729f
C44419 _1058_/a_381_47# net189 0.00496f
C44420 net245 _0405_ 0
C44421 _0461_ _0346_ 0.03307f
C44422 hold93/a_49_47# hold93/a_285_47# 0.22264f
C44423 hold58/a_49_47# _0211_ 0
C44424 _0222_ _0248_ 0
C44425 input32/a_75_212# _1042_/a_193_47# 0
C44426 _0289_ _0347_ 0.48295f
C44427 clknet_1_0__leaf__0459_ _0094_ 0.00735f
C44428 acc0.A\[14\] _0452_ 0
C44429 _0399_ _0115_ 0
C44430 _1000_/a_1059_315# _0244_ 0.03161f
C44431 _1000_/a_466_413# _0386_ 0
C44432 _1000_/a_634_159# _0388_ 0
C44433 VPWR _1029_/a_1059_315# 0.44235f
C44434 _1055_/a_891_413# net142 0.00976f
C44435 _0540_/a_51_297# _0540_/a_512_297# 0.0116f
C44436 _0982_/a_466_413# _0453_ 0
C44437 _0982_/a_381_47# _0452_ 0
C44438 _1048_/a_193_47# _1048_/a_381_47# 0.09503f
C44439 _1048_/a_634_159# _1048_/a_891_413# 0.03684f
C44440 _1048_/a_27_47# _1048_/a_561_413# 0.0027f
C44441 _1034_/a_193_47# clknet_1_1__leaf__0463_ 0.07561f
C44442 clkbuf_1_1__f__0460_/a_110_47# _1010_/a_27_47# 0.00204f
C44443 clknet_1_1__leaf__0464_ _0202_ 0.03751f
C44444 _0399_ _0796_/a_297_297# 0.00247f
C44445 _0096_ _0796_/a_79_21# 0
C44446 _0398_ _0796_/a_215_47# 0
C44447 _0294_ net102 0.01393f
C44448 clknet_1_0__leaf__0462_ VPWR 3.94272f
C44449 _0846_/a_512_297# _0447_ 0
C44450 _0179_ clkload2/Y 0.02739f
C44451 _0234_ _0350_ 0
C44452 _0385_ control0.add 0
C44453 _0113_ net149 0
C44454 _0981_/a_109_297# clknet_1_0__leaf_clk 0.0049f
C44455 net120 _0562_/a_150_297# 0
C44456 net33 net23 0.02736f
C44457 _0349_ _0334_ 0
C44458 _0223_ _0618_/a_79_21# 0.05489f
C44459 net187 hold73/a_391_47# 0
C44460 net45 _0774_/a_150_297# 0
C44461 _0172_ _0497_/a_150_297# 0
C44462 _0229_ net48 0.02264f
C44463 net152 _0544_/a_245_297# 0
C44464 _0546_/a_149_47# _0204_ 0
C44465 net32 _0544_/a_51_297# 0.0078f
C44466 _0546_/a_51_297# net18 0
C44467 _0357_ _0345_ 0.00252f
C44468 _0521_/a_299_297# net140 0
C44469 _0151_ _1054_/a_381_47# 0
C44470 net45 _0405_ 0
C44471 net59 hold15/a_285_47# 0
C44472 _1010_/a_891_413# _1010_/a_1017_47# 0.00617f
C44473 _1010_/a_634_159# net96 0
C44474 _0248_ net220 0
C44475 _0348_ _0195_ 0
C44476 _0464_ _0174_ 0
C44477 _0130_ _1015_/a_634_159# 0
C44478 clknet_0__0460_ _0350_ 0
C44479 _0956_/a_220_297# _0171_ 0
C44480 _0682_/a_68_297# acc0.A\[25\] 0.18011f
C44481 _1040_/a_634_159# _1040_/a_1017_47# 0
C44482 _1040_/a_466_413# _1040_/a_592_47# 0.00553f
C44483 hold26/a_49_47# _0536_/a_51_297# 0.02522f
C44484 hold74/a_285_47# acc0.A\[16\] 0.08388f
C44485 _0768_/a_27_47# _0310_ 0.03943f
C44486 _1017_/a_27_47# acc0.A\[18\] 0
C44487 _0979_/a_27_297# _0480_ 0.09461f
C44488 _0343_ _0237_ 0
C44489 _0432_ _0442_ 0
C44490 hold88/a_391_47# clknet_1_1__leaf__0465_ 0
C44491 _0642_/a_27_413# _0255_ 0
C44492 _0527_/a_109_297# net154 0.0015f
C44493 _1072_/a_27_47# _1072_/a_466_413# 0.26005f
C44494 _1072_/a_193_47# _1072_/a_634_159# 0.12729f
C44495 _0216_ _1027_/a_381_47# 0.02051f
C44496 clknet_0__0458_ _0825_/a_68_297# 0.00477f
C44497 _0841_/a_79_21# _0841_/a_297_297# 0.01735f
C44498 net88 _0217_ 0.06963f
C44499 _0100_ net150 0.02602f
C44500 VPWR _1019_/a_891_413# 0.17999f
C44501 _0714_/a_51_297# VPWR 0.46821f
C44502 hold88/a_49_47# _0088_ 0
C44503 _0640_/a_215_297# _0346_ 0
C44504 _0532_/a_81_21# clknet_1_1__leaf__0457_ 0.05637f
C44505 _0198_ clkbuf_1_1__f__0457_/a_110_47# 0
C44506 clknet_1_0__leaf__0462_ net48 0.54739f
C44507 _0793_/a_51_297# _0352_ 0
C44508 _0625_/a_59_75# _0399_ 0
C44509 _0537_/a_68_297# _1045_/a_1059_315# 0.01364f
C44510 clknet_0__0459_ _0347_ 0
C44511 _0343_ hold72/a_285_47# 0
C44512 net45 _1016_/a_1017_47# 0
C44513 _1067_/a_466_413# _1067_/a_592_47# 0.00553f
C44514 _1067_/a_634_159# _1067_/a_1017_47# 0
C44515 net9 _0987_/a_592_47# 0
C44516 _0136_ net180 0
C44517 hold36/a_49_47# hold37/a_285_47# 0.00183f
C44518 _0244_ _1018_/a_193_47# 0
C44519 clknet_1_0__leaf__0459_ _0393_ 0.03359f
C44520 _1036_/a_1059_315# _0208_ 0.00999f
C44521 _0429_ _0989_/a_27_47# 0
C44522 _0251_ _0989_/a_634_159# 0.00397f
C44523 _1001_/a_891_413# _0345_ 0
C44524 net205 _0134_ 0
C44525 hold31/a_49_47# hold31/a_391_47# 0.00188f
C44526 clknet_1_1__leaf__0460_ _1011_/a_193_47# 0
C44527 _0239_ _0779_/a_79_21# 0
C44528 hold12/a_391_47# net35 0.02248f
C44529 _0154_ input2/a_75_212# 0.00171f
C44530 hold35/a_391_47# A[10] 0.00373f
C44531 _0346_ _0992_/a_975_413# 0
C44532 _1050_/a_466_413# _0172_ 0
C44533 _1071_/a_466_413# _0169_ 0
C44534 net45 _0773_/a_35_297# 0
C44535 _0476_ _0564_/a_68_297# 0
C44536 net62 acc0.A\[6\] 0
C44537 VPWR net206 0.32042f
C44538 acc0.A\[17\] hold72/a_49_47# 0.28054f
C44539 _0239_ _0310_ 0.00109f
C44540 _0482_ _0479_ 0.10088f
C44541 control0.state\[1\] _1002_/a_466_413# 0
C44542 _0717_/a_209_297# _0717_/a_303_47# 0
C44543 net65 _0989_/a_975_413# 0
C44544 _0252_ _0989_/a_891_413# 0.04172f
C44545 _0343_ hold87/a_285_47# 0
C44546 _0195_ _0332_ 0.03604f
C44547 _0989_/a_634_159# _0989_/a_592_47# 0
C44548 _0346_ _0465_ 0.01445f
C44549 _0997_/a_27_47# _0997_/a_466_413# 0.26005f
C44550 _0997_/a_193_47# _0997_/a_634_159# 0.11072f
C44551 _1020_/a_634_159# clknet_1_0__leaf__0461_ 0
C44552 _0129_ hold92/a_285_47# 0
C44553 _0413_ _0218_ 0.04377f
C44554 _0181_ _0986_/a_466_413# 0
C44555 _0544_/a_240_47# _1042_/a_27_47# 0
C44556 _0544_/a_51_297# _1042_/a_1059_315# 0
C44557 _0544_/a_149_47# _1042_/a_193_47# 0
C44558 net36 clknet_1_0__leaf__0464_ 0
C44559 _0080_ VPWR 0.27643f
C44560 acc0.A\[31\] _0195_ 0
C44561 hold30/a_285_47# net46 0.01593f
C44562 clkbuf_0__0461_/a_110_47# net219 0.00304f
C44563 acc0.A\[16\] _0583_/a_109_297# 0.01058f
C44564 _0476_ clknet_1_1__leaf_clk 0.00344f
C44565 net213 _0103_ 0
C44566 _0331_ clknet_0__0462_ 0
C44567 _0992_/a_634_159# _0992_/a_592_47# 0
C44568 _0749_/a_299_297# _0369_ 0.0089f
C44569 VPWR _1051_/a_193_47# 0.31141f
C44570 acc0.A\[2\] _0346_ 0
C44571 _0312_ clkbuf_1_0__f__0462_/a_110_47# 0
C44572 net24 _0214_ 0
C44573 _0263_ _0843_/a_68_297# 0.00147f
C44574 _0570_/a_27_297# acc0.A\[25\] 0
C44575 VPWR _1045_/a_466_413# 0.25079f
C44576 _0402_ _0808_/a_368_297# 0.00191f
C44577 VPWR _1053_/a_1017_47# 0
C44578 _0125_ _1027_/a_592_47# 0
C44579 net216 _0693_/a_68_297# 0
C44580 _0280_ _0286_ 0.18666f
C44581 clknet_0__0458_ _0841_/a_79_21# 0.0066f
C44582 _0354_ _1029_/a_561_413# 0
C44583 _1014_/a_1017_47# acc0.A\[0\] 0
C44584 hold13/a_285_47# comp0.B\[5\] 0.08152f
C44585 hold13/a_49_47# comp0.B\[6\] 0.00282f
C44586 _0655_/a_109_93# _0347_ 0
C44587 _0793_/a_240_47# _0792_/a_80_21# 0
C44588 _0255_ _0218_ 0.02458f
C44589 _0274_ hold101/a_285_47# 0
C44590 hold46/a_49_47# hold26/a_49_47# 0.00377f
C44591 _0935_/a_27_47# _0465_ 0.11008f
C44592 _0963_/a_285_297# _0466_ 0
C44593 net10 _0544_/a_51_297# 0.00398f
C44594 _0465_ _1061_/a_193_47# 0.00394f
C44595 net45 net225 0.00919f
C44596 _1061_/a_193_47# _1061_/a_381_47# 0.10164f
C44597 _1061_/a_27_47# _1061_/a_561_413# 0.0027f
C44598 _1061_/a_634_159# _1061_/a_891_413# 0.03684f
C44599 input5/a_75_212# _0300_ 0
C44600 _0680_/a_472_297# _1009_/a_27_47# 0
C44601 net46 _0102_ 0
C44602 net51 _0754_/a_245_297# 0
C44603 net66 _0990_/a_634_159# 0.03435f
C44604 _0291_ _0990_/a_27_47# 0.00203f
C44605 acc0.A\[8\] _0990_/a_193_47# 0.0251f
C44606 net203 _0493_/a_27_47# 0
C44607 net160 input28/a_75_212# 0
C44608 _0313_ clknet_1_1__leaf__0460_ 0.28009f
C44609 _0629_/a_59_75# _0465_ 0.00232f
C44610 _0216_ _1026_/a_592_47# 0
C44611 _1054_/a_27_47# A[4] 0
C44612 _1007_/a_891_413# _0219_ 0.00104f
C44613 _0216_ net110 0.00108f
C44614 _0180_ hold83/a_285_47# 0.03227f
C44615 _0571_/a_27_297# _0570_/a_27_297# 0
C44616 _1035_/a_27_47# _1035_/a_634_159# 0.14145f
C44617 net182 A[10] 0.00117f
C44618 _0424_ acc0.A\[9\] 0.17941f
C44619 net171 _0207_ 0.18367f
C44620 pp[18] _0714_/a_245_297# 0
C44621 _0629_/a_59_75# acc0.A\[2\] 0.08219f
C44622 _0850_/a_150_297# _0345_ 0
C44623 _0558_/a_150_297# net26 0
C44624 _0959_/a_80_21# _1065_/a_27_47# 0
C44625 _0956_/a_32_297# _0175_ 0
C44626 net58 _0428_ 0
C44627 hold2/a_391_47# _1047_/a_1059_315# 0
C44628 _0183_ _1014_/a_891_413# 0.0012f
C44629 _0787_/a_209_297# _0091_ 0.01203f
C44630 _0787_/a_303_47# _0419_ 0.00306f
C44631 _0100_ control0.add 0
C44632 _0489_ _1069_/a_634_159# 0.0295f
C44633 _0260_ _0448_ 0.00369f
C44634 hold15/a_49_47# _0338_ 0
C44635 _1065_/a_891_413# clknet_1_0__leaf__0457_ 0
C44636 acc0.A\[1\] _0197_ 0
C44637 _0661_/a_27_297# _0290_ 0
C44638 acc0.A\[12\] _0302_ 0
C44639 VPWR _0637_/a_139_47# 0
C44640 hold58/a_49_47# _0210_ 0
C44641 _0131_ _0215_ 0
C44642 _0397_ _0392_ 0
C44643 _0222_ _0755_/a_109_297# 0.00349f
C44644 _0216_ clkbuf_1_1__f__0457_/a_110_47# 0.00392f
C44645 net76 _0990_/a_466_413# 0
C44646 _0343_ _0991_/a_561_413# 0
C44647 net24 _0207_ 0
C44648 _0586_/a_27_47# _0345_ 0.00276f
C44649 _0376_ _0237_ 0
C44650 VPWR _1028_/a_592_47# 0
C44651 _1069_/a_891_413# _1069_/a_975_413# 0.00851f
C44652 _1069_/a_27_47# clknet_1_0__leaf_clk 0.35436f
C44653 _1069_/a_381_47# _1069_/a_561_413# 0.00123f
C44654 _1056_/a_634_159# net66 0
C44655 _0189_ acc0.A\[11\] 0
C44656 _0402_ _0304_ 0
C44657 _0854_/a_79_21# _0181_ 0.05623f
C44658 _0343_ _0392_ 0.03171f
C44659 net117 _1030_/a_27_47# 0
C44660 B[13] _0140_ 0
C44661 comp0.B\[14\] _0545_/a_68_297# 0
C44662 _0349_ output59/a_27_47# 0
C44663 VPWR input30/a_75_212# 0.27084f
C44664 _0552_/a_68_297# _0176_ 0.14619f
C44665 _1059_/a_891_413# acc0.A\[13\] 0.03192f
C44666 clknet_0__0465_ _0990_/a_1059_315# 0.01731f
C44667 _1059_/a_27_47# _0185_ 0.03562f
C44668 pp[8] _1055_/a_27_47# 0.00144f
C44669 _0662_/a_81_21# _0346_ 0.00164f
C44670 comp0.B\[1\] control0.sh 0
C44671 _0753_/a_297_297# _0223_ 0.00113f
C44672 _1062_/a_27_47# hold84/a_391_47# 0.00816f
C44673 net22 _0498_/a_51_297# 0
C44674 net225 _0587_/a_27_47# 0
C44675 _1041_/a_1059_315# _1040_/a_466_413# 0.00365f
C44676 _1041_/a_891_413# _1040_/a_634_159# 0.0012f
C44677 _0997_/a_634_159# _0411_ 0
C44678 _0096_ _1017_/a_1059_315# 0
C44679 _0399_ _1017_/a_891_413# 0
C44680 _0443_ _0838_/a_109_297# 0.01202f
C44681 hold55/a_391_47# net87 0
C44682 pp[15] pp[16] 0.25399f
C44683 pp[20] pp[21] 0.17884f
C44684 hold64/a_285_47# hold64/a_391_47# 0.41909f
C44685 _0624_/a_59_75# net62 0.22053f
C44686 hold23/a_285_47# VPWR 0.34101f
C44687 clknet_1_0__leaf__0460_ _1063_/a_193_47# 0
C44688 _0577_/a_27_297# _0577_/a_109_297# 0.17136f
C44689 B[12] hold51/a_391_47# 0
C44690 _1030_/a_561_413# net209 0
C44691 _0388_ _0242_ 0
C44692 _0556_/a_68_297# net160 0
C44693 hold26/a_49_47# comp0.B\[14\] 0
C44694 _1039_/a_1059_315# net171 0.00155f
C44695 _0176_ _0204_ 0.01056f
C44696 _0172_ _0206_ 0.02344f
C44697 _0337_ pp[28] 0.00216f
C44698 hold89/a_285_47# _0479_ 0
C44699 hold96/a_391_47# net110 0
C44700 _0645_/a_47_47# _0670_/a_79_21# 0.00364f
C44701 acc0.A\[22\] _1022_/a_634_159# 0.00111f
C44702 _0183_ _1022_/a_193_47# 0
C44703 _0217_ _1022_/a_466_413# 0
C44704 _0260_ _0444_ 0
C44705 _0221_ _0705_/a_59_75# 0
C44706 _0620_/a_113_47# clknet_1_1__leaf__0458_ 0
C44707 clknet_1_1__leaf__0458_ _0989_/a_27_47# 0
C44708 hold1/a_49_47# clknet_1_1__leaf__0458_ 0.00501f
C44709 clknet_1_0__leaf__0460_ _0460_ 0.11056f
C44710 _0538_/a_240_47# _0201_ 0
C44711 hold6/a_391_47# _0176_ 0
C44712 clknet_1_0__leaf__0463_ _0498_/a_51_297# 0.00685f
C44713 hold30/a_391_47# VPWR 0.17841f
C44714 comp0.B\[5\] _0132_ 0
C44715 _0146_ acc0.A\[15\] 0
C44716 hold67/a_391_47# acc0.A\[9\] 0.00753f
C44717 _0524_/a_27_297# _0524_/a_109_47# 0.00393f
C44718 _1014_/a_891_413# acc0.A\[15\] 0
C44719 _1022_/a_891_413# net151 0
C44720 _0646_/a_129_47# _0218_ 0
C44721 pp[25] _0572_/a_27_297# 0
C44722 _1065_/a_466_413# _1062_/a_891_413# 0
C44723 hold22/a_49_47# _0191_ 0.03035f
C44724 hold22/a_391_47# net15 0.02501f
C44725 net64 _0990_/a_193_47# 0
C44726 clknet_1_0__leaf__0459_ _1019_/a_891_413# 0.00991f
C44727 net87 _1019_/a_466_413# 0
C44728 _0492_/a_27_47# acc0.A\[15\] 0.04701f
C44729 acc0.A\[17\] clknet_0__0461_ 0.17914f
C44730 _1003_/a_193_47# _0974_/a_222_93# 0
C44731 hold12/a_285_47# net159 0.01021f
C44732 net199 _1025_/a_891_413# 0
C44733 acc0.A\[26\] _0321_ 0.00167f
C44734 _0994_/a_466_413# _0994_/a_592_47# 0.00553f
C44735 _0994_/a_634_159# _0994_/a_1017_47# 0
C44736 _1020_/a_975_413# clknet_1_0__leaf__0457_ 0
C44737 _0284_ _0417_ 0
C44738 _0579_/a_109_297# net223 0
C44739 net211 _0772_/a_215_47# 0
C44740 _0779_/a_510_47# _0396_ 0.00122f
C44741 _0779_/a_297_297# _0097_ 0.00204f
C44742 _0287_ _0090_ 0
C44743 _0462_ _0324_ 0.09109f
C44744 _1055_/a_592_47# net179 0.00301f
C44745 _0500_/a_27_47# _1048_/a_27_47# 0
C44746 _1023_/a_891_413# net51 0.00191f
C44747 _0457_ clknet_1_0__leaf__0460_ 0.00138f
C44748 hold56/a_285_47# _0175_ 0
C44749 _0290_ _0990_/a_27_47# 0
C44750 _0835_/a_215_47# _0270_ 0
C44751 _0464_ _1046_/a_193_47# 0
C44752 hold22/a_391_47# _1053_/a_1059_315# 0.01554f
C44753 _0855_/a_384_47# _0350_ 0
C44754 hold14/a_285_47# net161 0.0102f
C44755 net36 _1047_/a_592_47# 0
C44756 net161 input27/a_75_212# 0
C44757 _0399_ net223 0
C44758 _0503_/a_109_297# _0182_ 0.01263f
C44759 _0993_/a_27_47# _0993_/a_466_413# 0.27314f
C44760 _0993_/a_193_47# _0993_/a_634_159# 0.12729f
C44761 _1058_/a_27_47# _0156_ 0.104f
C44762 _0647_/a_285_47# net80 0
C44763 clknet_1_0__leaf__0459_ net206 0
C44764 _1065_/a_27_47# _0173_ 0
C44765 _0721_/a_27_47# _0526_/a_27_47# 0
C44766 comp0.B\[1\] net157 0
C44767 _1039_/a_193_47# _1039_/a_381_47# 0.09503f
C44768 _1039_/a_634_159# _1039_/a_891_413# 0.03684f
C44769 _1039_/a_27_47# _1039_/a_561_413# 0.00163f
C44770 _0251_ _0258_ 0.00103f
C44771 clkbuf_0__0461_/a_110_47# _0352_ 0.08893f
C44772 _0258_ _0640_/a_109_53# 0
C44773 _0557_/a_240_47# clknet_0__0463_ 0
C44774 _1020_/a_381_47# _0457_ 0.00396f
C44775 acc0.A\[12\] net6 0
C44776 _0578_/a_27_297# net1 0.01632f
C44777 _0280_ _0672_/a_79_21# 0.09562f
C44778 _0279_ _0672_/a_510_47# 0
C44779 net169 _0191_ 0.00566f
C44780 _0985_/a_891_413# net170 0
C44781 A[12] _0512_/a_109_297# 0.00177f
C44782 _1056_/a_193_47# net64 0
C44783 net247 clkbuf_1_1__f__0457_/a_110_47# 0
C44784 _0498_/a_240_47# clknet_1_1__leaf__0457_ 0
C44785 _1010_/a_891_413# _0332_ 0
C44786 _0172_ _1046_/a_1059_315# 0
C44787 hold14/a_285_47# net26 0.00463f
C44788 _1049_/a_27_47# _0148_ 0
C44789 net242 clknet_1_1__leaf__0462_ 0.03679f
C44790 net26 input27/a_75_212# 0
C44791 _1026_/a_634_159# _1026_/a_1059_315# 0
C44792 _1026_/a_27_47# _1026_/a_381_47# 0.06222f
C44793 _1026_/a_193_47# _1026_/a_891_413# 0.19685f
C44794 _0305_ _0240_ 0.0216f
C44795 _0733_/a_222_93# _0321_ 0.00729f
C44796 _0733_/a_544_297# _0360_ 0.00275f
C44797 net188 net37 0.02331f
C44798 _0646_/a_47_47# A[13] 0.00182f
C44799 _0646_/a_285_47# input5/a_75_212# 0
C44800 _0985_/a_1059_315# clknet_1_0__leaf__0458_ 0
C44801 _1021_/a_466_413# clknet_1_0__leaf__0460_ 0.00101f
C44802 _0305_ _0369_ 1.61824f
C44803 hold10/a_285_47# _1047_/a_27_47# 0
C44804 _0234_ _1005_/a_1059_315# 0.00518f
C44805 _0273_ _0399_ 0
C44806 VPWR _0774_/a_150_297# 0.00115f
C44807 net140 _1053_/a_561_413# 0
C44808 net169 _1053_/a_381_47# 0
C44809 _0982_/a_891_413# _0399_ 0
C44810 _0195_ _0117_ 0.03257f
C44811 _0786_/a_80_21# _0346_ 0
C44812 _0179_ _0146_ 0.02957f
C44813 VPWR _0405_ 0.93393f
C44814 _0217_ _1067_/a_891_413# 0
C44815 hold97/a_49_47# clkbuf_1_1__f__0460_/a_110_47# 0
C44816 _1024_/a_27_47# _0122_ 0.08151f
C44817 _1024_/a_193_47# net110 0.00544f
C44818 _1024_/a_1059_315# _1024_/a_1017_47# 0
C44819 _0854_/a_79_21# _1018_/a_27_47# 0
C44820 hold45/a_391_47# _0186_ 0
C44821 _0595_/a_109_297# _0228_ 0
C44822 _0216_ _0692_/a_113_47# 0
C44823 _0245_ acc0.A\[18\] 0.05023f
C44824 _0134_ net160 0
C44825 _0426_ _0425_ 0.10177f
C44826 _0625_/a_59_75# _0619_/a_68_297# 0
C44827 _0195_ net43 0.07562f
C44828 net58 _0258_ 0
C44829 net203 clkbuf_1_1__f_clk/a_110_47# 0
C44830 _1014_/a_193_47# _0181_ 0
C44831 _0121_ hold29/a_285_47# 0
C44832 _0453_ net206 0
C44833 VPWR _0356_ 0.44745f
C44834 _1036_/a_466_413# B[2] 0
C44835 _1036_/a_634_159# net25 0
C44836 _0336_ _0219_ 0.00136f
C44837 _0355_ hold62/a_285_47# 0
C44838 _0438_ acc0.A\[8\] 0.01333f
C44839 acc0.A\[5\] _0834_/a_109_297# 0
C44840 _0835_/a_78_199# acc0.A\[4\] 0.00341f
C44841 _0422_ clknet_1_1__leaf__0465_ 0.00129f
C44842 _0098_ _0386_ 0
C44843 _0574_/a_373_47# VPWR 0
C44844 hold89/a_391_47# VPWR 0.16451f
C44845 _0786_/a_80_21# _0992_/a_466_413# 0
C44846 _0540_/a_51_297# _0142_ 0.10333f
C44847 _0540_/a_149_47# net20 0
C44848 _0953_/a_32_297# _1040_/a_1059_315# 0
C44849 _0080_ _0453_ 0
C44850 clk _1064_/a_592_47# 0
C44851 net243 _0217_ 0.06915f
C44852 _1048_/a_891_413# net134 0
C44853 _0402_ _0811_/a_384_47# 0.01047f
C44854 acc0.A\[14\] _0277_ 0.00487f
C44855 _0831_/a_35_297# _0434_ 0.2556f
C44856 _0253_ _0826_/a_27_53# 0
C44857 _0195_ _0999_/a_27_47# 0
C44858 VPWR comp0.B\[15\] 0.5067f
C44859 _1020_/a_27_47# _0208_ 0
C44860 _1068_/a_1059_315# _0468_ 0.09016f
C44861 net149 _0345_ 0.14341f
C44862 _1041_/a_27_47# _1041_/a_634_159# 0.13601f
C44863 _0343_ _1013_/a_1059_315# 0.0353f
C44864 net1 _0180_ 0
C44865 hold99/a_49_47# _0993_/a_27_47# 0
C44866 _0234_ _0751_/a_183_297# 0
C44867 _0375_ _0751_/a_29_53# 0.1132f
C44868 _0416_ _0803_/a_150_297# 0
C44869 _1059_/a_27_47# _0289_ 0
C44870 _0172_ _0270_ 0
C44871 VPWR _0773_/a_35_297# 0.16256f
C44872 _1015_/a_466_413# comp0.B\[15\] 0
C44873 input33/a_75_212# B[0] 0
C44874 init input17/a_75_212# 0.0072f
C44875 _0302_ net42 0.01176f
C44876 _0372_ _0771_/a_215_297# 0
C44877 _0248_ _0771_/a_298_297# 0
C44878 hold39/a_391_47# net231 0
C44879 _1057_/a_27_47# _0514_/a_109_297# 0
C44880 hold76/a_285_47# _1001_/a_27_47# 0
C44881 _0855_/a_81_21# acc0.A\[1\] 0
C44882 _0212_ net33 0
C44883 _0607_/a_373_47# acc0.A\[17\] 0.00157f
C44884 hold2/a_49_47# net149 0.00129f
C44885 _0596_/a_59_75# _0486_ 0
C44886 _0310_ _0309_ 0.03494f
C44887 clknet_0__0465_ _0439_ 0.00114f
C44888 B[11] net128 0.00224f
C44889 net78 VPWR 0.33925f
C44890 _0129_ _0220_ 0.44263f
C44891 VPWR clknet_0__0465_ 2.37236f
C44892 _1056_/a_561_413# _0189_ 0
C44893 _0830_/a_215_47# _0218_ 0
C44894 clknet_1_0__leaf__0465_ _1054_/a_592_47# 0
C44895 hold44/a_49_47# _1029_/a_193_47# 0
C44896 hold44/a_285_47# _1029_/a_27_47# 0.00329f
C44897 clkbuf_1_0__f__0457_/a_110_47# _0610_/a_59_75# 0
C44898 net226 _0488_ 0.0018f
C44899 clknet_0__0458_ _0627_/a_215_53# 0.00629f
C44900 _0480_ _0169_ 0
C44901 _0293_ _0291_ 0
C44902 _0623_/a_109_297# _0150_ 0
C44903 _0249_ _1006_/a_381_47# 0
C44904 _0250_ _1006_/a_891_413# 0
C44905 _1072_/a_1059_315# _1072_/a_1017_47# 0
C44906 _0841_/a_215_47# _0084_ 0.00406f
C44907 _0155_ net37 0.00117f
C44908 net225 VPWR 0.14782f
C44909 _0317_ _0360_ 0
C44910 _0713_/a_27_47# clkbuf_0__0457_/a_110_47# 0.02101f
C44911 _0254_ _0346_ 0.10094f
C44912 clknet_1_0__leaf__0461_ hold60/a_49_47# 0.00857f
C44913 hold38/a_391_47# hold39/a_285_47# 0.0043f
C44914 hold38/a_285_47# hold39/a_391_47# 0.0043f
C44915 _0554_/a_68_297# net160 0.18754f
C44916 net100 clkbuf_1_1__f__0457_/a_110_47# 0.00351f
C44917 _1013_/a_466_413# net60 0
C44918 _0471_ _1062_/a_634_159# 0.00148f
C44919 hold36/a_391_47# clknet_1_0__leaf__0465_ 0.00569f
C44920 VPWR _1025_/a_891_413# 0.21155f
C44921 _0946_/a_30_53# _0466_ 0.19458f
C44922 _1055_/a_634_159# _0186_ 0
C44923 _0257_ clknet_1_1__leaf__0458_ 0.01667f
C44924 net61 _0624_/a_145_75# 0
C44925 clknet_1_1__leaf__0462_ hold92/a_49_47# 0.02568f
C44926 _0254_ net65 0
C44927 net105 _1015_/a_381_47# 0
C44928 _1012_/a_466_413# _0722_/a_215_47# 0.00141f
C44929 net64 _0438_ 0.1397f
C44930 _0427_ net47 0
C44931 _0476_ _0559_/a_512_297# 0.00149f
C44932 _0822_/a_109_297# VPWR 0.0071f
C44933 net55 acc0.A\[29\] 0.20068f
C44934 control0.state\[1\] _0100_ 0
C44935 net87 _0352_ 0.01115f
C44936 _0363_ _0359_ 0
C44937 clknet_1_0__leaf__0462_ pp[22] 0
C44938 hold75/a_391_47# net233 0
C44939 _0997_/a_1059_315# _0997_/a_1017_47# 0
C44940 _1053_/a_634_159# _0150_ 0
C44941 _1037_/a_1059_315# net24 0
C44942 net203 VPWR 0.29541f
C44943 _0664_/a_297_47# _0346_ 0.00603f
C44944 _0104_ _0462_ 0.00489f
C44945 net18 _1042_/a_891_413# 0.00999f
C44946 net198 _1042_/a_381_47# 0
C44947 _0140_ _1042_/a_634_159# 0.00527f
C44948 clknet_1_0__leaf__0457_ hold93/a_285_47# 0.00427f
C44949 VPWR _1044_/a_634_159# 0.18504f
C44950 clknet_1_0__leaf__0464_ _0527_/a_27_297# 0.00263f
C44951 VPWR _0815_/a_199_47# 0
C44952 hold100/a_391_47# _0345_ 0.00101f
C44953 clkbuf_1_0__f__0459_/a_110_47# _1059_/a_466_413# 0
C44954 clknet_0__0459_ _1059_/a_27_47# 0.001f
C44955 _0349_ _1010_/a_381_47# 0
C44956 hold7/a_391_47# net11 0.00303f
C44957 VPWR net184 0.22698f
C44958 hold88/a_285_47# _0399_ 0.00156f
C44959 _0783_/a_215_47# _0352_ 0.00336f
C44960 _0661_/a_27_297# _0656_/a_59_75# 0
C44961 _0243_ _0773_/a_117_297# 0.0011f
C44962 _0390_ _0773_/a_35_297# 0
C44963 _0756_/a_47_47# _0756_/a_285_47# 0.01755f
C44964 _0407_ _0400_ 0.08847f
C44965 _1001_/a_634_159# _0461_ 0.00586f
C44966 _0342_ clknet_1_1__leaf__0461_ 0
C44967 _1027_/a_634_159# _1027_/a_592_47# 0
C44968 _0643_/a_103_199# _0643_/a_337_297# 0.01015f
C44969 hold87/a_391_47# net234 0.13055f
C44970 _0181_ _0240_ 0.0226f
C44971 _0241_ _0611_/a_68_297# 0.16768f
C44972 _0366_ _0367_ 0.11733f
C44973 _0253_ _0087_ 0
C44974 VPWR _0849_/a_215_47# 0.00449f
C44975 net42 net6 0.03899f
C44976 acc0.A\[8\] clknet_1_1__leaf__0465_ 0.00349f
C44977 VPWR _1032_/a_561_413# 0.00323f
C44978 _0369_ _0181_ 1.67739f
C44979 _0343_ _0222_ 0.22508f
C44980 _1061_/a_891_413# net147 0
C44981 clknet_1_0__leaf__0465_ _0522_/a_373_47# 0
C44982 clkbuf_0__0461_/a_110_47# _0613_/a_109_297# 0
C44983 comp0.B\[5\] net25 0.1914f
C44984 clknet_0__0457_ _0181_ 0.07704f
C44985 clknet_1_0__leaf__0462_ _1023_/a_27_47# 0.00549f
C44986 net15 A[7] 0
C44987 _0555_/a_149_47# comp0.B\[5\] 0.00108f
C44988 _0462_ _0745_/a_109_47# 0
C44989 net248 _0440_ 0
C44990 hold21/a_391_47# VPWR 0.18127f
C44991 hold10/a_285_47# net133 0
C44992 clknet_1_0__leaf__0464_ _1061_/a_27_47# 0
C44993 net126 net124 0
C44994 net26 net17 0
C44995 hold29/a_285_47# _0380_ 0
C44996 _1065_/a_193_47# _0161_ 0
C44997 _0991_/a_193_47# clknet_1_1__leaf__0465_ 0
C44998 _0571_/a_27_297# _0126_ 0
C44999 _0125_ _0570_/a_27_297# 0
C45000 _1035_/a_891_413# _1035_/a_975_413# 0.00851f
C45001 _1035_/a_27_47# net121 0.23156f
C45002 _1035_/a_381_47# _1035_/a_561_413# 0.00123f
C45003 _0668_/a_79_21# _0668_/a_297_47# 0.03259f
C45004 _0399_ _0086_ 0.02194f
C45005 _1012_/a_27_47# _0704_/a_68_297# 0
C45006 _0389_ _0350_ 0.01406f
C45007 hold39/a_49_47# _1034_/a_27_47# 0
C45008 hold76/a_391_47# clknet_1_0__leaf__0461_ 0
C45009 _0946_/a_30_53# _1064_/a_193_47# 0
C45010 clkbuf_1_1__f__0462_/a_110_47# net97 0.00121f
C45011 _1051_/a_27_47# _0172_ 0.07447f
C45012 clkbuf_0__0464_/a_110_47# net174 0
C45013 _0591_/a_109_297# VPWR 0.00563f
C45014 net44 net117 0
C45015 _0489_ clknet_1_0__leaf_clk 0.08148f
C45016 _0217_ _0366_ 0
C45017 net124 input8/a_75_212# 0
C45018 _0809_/a_299_297# _0809_/a_384_47# 0
C45019 VPWR _0533_/a_109_47# 0
C45020 _0172_ _1045_/a_634_159# 0.02169f
C45021 _0287_ _0401_ 0.06573f
C45022 _0293_ _0290_ 0.06186f
C45023 _0289_ _0425_ 0.00333f
C45024 hold69/a_285_47# _0326_ 0
C45025 _1062_/a_1059_315# hold93/a_49_47# 0
C45026 VPWR hold71/a_285_47# 0.32053f
C45027 _1030_/a_193_47# _0334_ 0
C45028 VPWR _0387_ 1.12978f
C45029 clknet_1_1__leaf__0459_ _1013_/a_634_159# 0
C45030 _0460_ hold94/a_285_47# 0.00145f
C45031 VPWR _0546_/a_149_47# 0.00124f
C45032 net76 _0088_ 0.00178f
C45033 clknet_1_1__leaf__0463_ _0171_ 0
C45034 acc0.A\[29\] _1029_/a_592_47# 0
C45035 _1011_/a_193_47# _0726_/a_240_47# 0.00146f
C45036 _1011_/a_634_159# _0726_/a_149_47# 0
C45037 _1011_/a_891_413# _0726_/a_51_297# 0.00143f
C45038 _1033_/a_27_47# _1065_/a_1059_315# 0
C45039 clknet_1_1__leaf__0460_ _0321_ 0.03094f
C45040 net32 _1043_/a_27_47# 0
C45041 net152 _1043_/a_193_47# 0
C45042 clknet_1_1__leaf__0460_ clkbuf_0__0460_/a_110_47# 0.03389f
C45043 _0233_ _0232_ 0.02655f
C45044 hold78/a_285_47# _0218_ 0
C45045 control0.sh _0496_/a_27_47# 0
C45046 clknet_1_0__leaf__0459_ _0773_/a_35_297# 0
C45047 _1041_/a_1059_315# net174 0
C45048 net45 _0340_ 0.00401f
C45049 net125 _1061_/a_891_413# 0.00416f
C45050 _0734_/a_47_47# _0318_ 0.05978f
C45051 _0399_ _1016_/a_193_47# 0
C45052 _0239_ _0309_ 0.04298f
C45053 _0967_/a_109_93# _0466_ 0
C45054 clknet_1_1__leaf__0458_ net11 0.02355f
C45055 control0.state\[1\] hold39/a_391_47# 0
C45056 _0466_ _0487_ 0.37127f
C45057 _0577_/a_373_47# _0183_ 0.00301f
C45058 _0577_/a_109_297# _0120_ 0.0037f
C45059 _0429_ clknet_1_1__leaf__0458_ 0
C45060 _0195_ _1018_/a_193_47# 0.04625f
C45061 net156 _1026_/a_27_47# 0
C45062 net33 _0161_ 0
C45063 net47 net142 0
C45064 _0553_/a_245_297# net171 0
C45065 net58 _0988_/a_193_47# 0.01907f
C45066 _0640_/a_392_297# clknet_1_1__leaf__0458_ 0
C45067 net8 _0171_ 0.0432f
C45068 _0467_ _1067_/a_634_159# 0
C45069 acc0.A\[5\] net9 0.01986f
C45070 _0568_/a_109_297# net209 0.00234f
C45071 net208 hold62/a_49_47# 0.12843f
C45072 _0481_ _1064_/a_891_413# 0
C45073 hold15/a_49_47# acc0.A\[31\] 0.30383f
C45074 _0990_/a_27_47# _0986_/a_1059_315# 0
C45075 _0645_/a_377_297# _0302_ 0.00299f
C45076 _0217_ net151 0.0442f
C45077 _0508_/a_299_297# _0345_ 0
C45078 _0563_/a_512_297# _0173_ 0
C45079 _0579_/a_109_297# clkbuf_0__0457_/a_110_47# 0
C45080 _0343_ acc0.A\[9\] 0
C45081 _0132_ hold84/a_49_47# 0
C45082 net183 _0143_ 0.32419f
C45083 hold58/a_285_47# _1034_/a_193_47# 0
C45084 hold58/a_391_47# _1034_/a_27_47# 0
C45085 _0227_ _0377_ 0
C45086 VPWR _0382_ 0.40069f
C45087 net106 _1015_/a_891_413# 0
C45088 net64 clknet_1_1__leaf__0465_ 0.05749f
C45089 net9 _0528_/a_299_297# 0.01574f
C45090 input18/a_75_212# B[11] 0.002f
C45091 pp[11] _0993_/a_891_413# 0
C45092 pp[25] _0124_ 0
C45093 _1065_/a_891_413# _0160_ 0
C45094 net36 acc0.A\[14\] 0
C45095 net87 net207 0
C45096 _0399_ clkbuf_0__0457_/a_110_47# 0.00145f
C45097 net73 acc0.A\[6\] 0
C45098 net89 _0974_/a_79_199# 0
C45099 _0995_/a_27_47# net41 0
C45100 net211 _1019_/a_634_159# 0
C45101 _0217_ _0580_/a_109_47# 0.00217f
C45102 _0183_ _0580_/a_27_297# 0.19867f
C45103 _0298_ _0798_/a_199_47# 0.01105f
C45104 net30 input30/a_75_212# 0.10876f
C45105 _0299_ _0798_/a_113_297# 0
C45106 _0982_/a_381_47# net36 0.0161f
C45107 net55 _0363_ 0
C45108 net78 _0283_ 0
C45109 _0343_ _0670_/a_79_21# 0
C45110 _0476_ _1036_/a_193_47# 0
C45111 _0423_ clknet_1_1__leaf__0465_ 0.02323f
C45112 net45 _1013_/a_381_47# 0.00631f
C45113 _0461_ _0782_/a_27_47# 0
C45114 hold91/a_285_47# acc0.A\[13\] 0
C45115 _0179_ _1048_/a_381_47# 0.00928f
C45116 hold35/a_49_47# net66 0
C45117 _0220_ hold61/a_285_47# 0.03239f
C45118 _0972_/a_93_21# net231 0.01546f
C45119 net177 pp[23] 0.00191f
C45120 net58 net72 0.00364f
C45121 _0538_/a_51_297# comp0.B\[10\] 0
C45122 _1043_/a_27_47# _1042_/a_1059_315# 0.01576f
C45123 _1043_/a_634_159# _1042_/a_634_159# 0
C45124 _1043_/a_1059_315# _1042_/a_27_47# 0.01576f
C45125 _1043_/a_193_47# _1042_/a_466_413# 0
C45126 _1043_/a_466_413# _1042_/a_193_47# 0
C45127 net45 acc0.A\[16\] 0.12372f
C45128 _1055_/a_466_413# net74 0
C45129 net236 _0487_ 0.03301f
C45130 _0376_ _0222_ 0.43449f
C45131 hold7/a_391_47# clknet_1_1__leaf__0458_ 0.0585f
C45132 _0182_ _0526_/a_27_47# 0
C45133 clkbuf_0__0461_/a_110_47# hold72/a_285_47# 0.02454f
C45134 clknet_1_0__leaf__0463_ A[15] 0.02828f
C45135 _1030_/a_27_47# _0704_/a_68_297# 0
C45136 _0642_/a_27_413# _0989_/a_27_47# 0
C45137 net17 hold84/a_285_47# 0
C45138 _0993_/a_1059_315# _0993_/a_1017_47# 0
C45139 net144 net192 0.0751f
C45140 _0268_ _0840_/a_68_297# 0
C45141 pp[27] _1030_/a_27_47# 0.00111f
C45142 _0627_/a_215_53# _0627_/a_109_93# 0.13675f
C45143 hold85/a_285_47# _0471_ 0
C45144 _1039_/a_1059_315# _0553_/a_51_297# 0.00114f
C45145 _1039_/a_891_413# net125 0
C45146 _0742_/a_299_297# _0366_ 0.08607f
C45147 _0742_/a_81_21# _0315_ 0.057f
C45148 _0182_ net9 0.0019f
C45149 net54 acc0.A\[25\] 0.01351f
C45150 _0278_ _0669_/a_29_53# 0
C45151 _0730_/a_79_21# _0730_/a_215_47# 0.04584f
C45152 _0535_/a_68_297# _1040_/a_1059_315# 0
C45153 net178 pp[1] 0
C45154 _0677_/a_377_297# _0240_ 0.00249f
C45155 _0343_ _0707_/a_544_297# 0
C45156 pp[28] _0333_ 0.05171f
C45157 clkbuf_0__0464_/a_110_47# clknet_0__0464_ 1.67181f
C45158 _0195_ _0708_/a_68_297# 0
C45159 net10 _1043_/a_27_47# 0.00405f
C45160 net234 _0264_ 0.05385f
C45161 _0266_ _0350_ 0.00917f
C45162 _0473_ control0.reset 0
C45163 _0714_/a_51_297# _1031_/a_634_159# 0
C45164 net48 _0382_ 0
C45165 net63 _0830_/a_297_297# 0.0038f
C45166 _0147_ _0196_ 0
C45167 _0485_ _1064_/a_634_159# 0.00209f
C45168 _0487_ _1064_/a_193_47# 0
C45169 net135 net170 0.0019f
C45170 _0747_/a_79_21# _0219_ 0.00312f
C45171 _1026_/a_1059_315# net112 0
C45172 _1026_/a_27_47# acc0.A\[26\] 0
C45173 _1059_/a_891_413# VPWR 0.19115f
C45174 _1054_/a_891_413# acc0.A\[5\] 0
C45175 _0985_/a_381_47# _0449_ 0
C45176 _0465_ _1047_/a_466_413# 0.00463f
C45177 _0119_ clknet_1_0__leaf__0460_ 0.01271f
C45178 _0472_ _1061_/a_466_413# 0
C45179 _0111_ _0567_/a_109_297# 0
C45180 _0216_ _0330_ 0
C45181 _0817_/a_81_21# _0817_/a_266_47# 0.04342f
C45182 clknet_1_1__leaf__0460_ _1009_/a_27_47# 0.03552f
C45183 _0181_ _1009_/a_561_413# 0
C45184 _0312_ _0324_ 0.03313f
C45185 net150 control0.add 0.02285f
C45186 _0542_/a_245_297# net20 0
C45187 net54 _0571_/a_27_297# 0.00286f
C45188 net66 A[9] 0
C45189 _0256_ _0345_ 0
C45190 hold47/a_49_47# _0527_/a_109_47# 0
C45191 hold66/a_49_47# net213 0
C45192 _0230_ _0754_/a_240_47# 0.04355f
C45193 _0598_/a_382_297# _0219_ 0.00163f
C45194 _0229_ _0345_ 0
C45195 _0789_/a_75_199# _0405_ 0.11073f
C45196 _0662_/a_81_21# _0259_ 0.06841f
C45197 clknet_1_1__leaf__0459_ hold70/a_391_47# 0.01736f
C45198 _0536_/a_51_297# _1061_/a_193_47# 0
C45199 net161 B[2] 0
C45200 hold99/a_391_47# pp[11] 0.00123f
C45201 _0182_ _0175_ 0
C45202 _0174_ _1040_/a_1059_315# 0.00365f
C45203 _1037_/a_193_47# _1037_/a_381_47# 0.09503f
C45204 _1037_/a_634_159# _1037_/a_891_413# 0.03684f
C45205 _1037_/a_27_47# _1037_/a_561_413# 0.0027f
C45206 pp[16] _0997_/a_592_47# 0
C45207 _0218_ _0989_/a_27_47# 0
C45208 hold53/a_391_47# net52 0
C45209 _0180_ acc0.A\[3\] 0.08233f
C45210 _0199_ _0147_ 0
C45211 _0402_ _0992_/a_1059_315# 0
C45212 _0217_ _0378_ 0
C45213 _1008_/a_27_47# _0687_/a_59_75# 0
C45214 acc0.A\[3\] net218 0
C45215 comp0.B\[10\] _1040_/a_381_47# 0
C45216 _0369_ _0507_/a_373_47# 0
C45217 _0472_ net24 0.3449f
C45218 _1029_/a_27_47# _0219_ 0
C45219 _0216_ _0242_ 1.08584f
C45220 _0180_ control0.sh 0.23949f
C45221 _0227_ net109 0
C45222 VPWR _1005_/a_634_159# 0.19177f
C45223 net67 acc0.A\[11\] 0.0246f
C45224 _0790_/a_285_297# net42 0.07614f
C45225 _0369_ hold82/a_391_47# 0.01286f
C45226 _0201_ _0473_ 0.07349f
C45227 _1041_/a_891_413# _1041_/a_975_413# 0.00851f
C45228 _1041_/a_381_47# _1041_/a_561_413# 0.00123f
C45229 VPWR _0519_/a_81_21# 0.1999f
C45230 _0228_ hold3/a_49_47# 0
C45231 VPWR _0991_/a_592_47# 0
C45232 _0690_/a_68_297# _1008_/a_891_413# 0
C45233 _0399_ net41 0.08271f
C45234 B[2] net26 0
C45235 net22 comp0.B\[12\] 0
C45236 _1054_/a_1059_315# _0180_ 0.00589f
C45237 clkbuf_1_1__f__0462_/a_110_47# _1010_/a_27_47# 0
C45238 hold30/a_285_47# _1023_/a_193_47# 0
C45239 hold30/a_391_47# _1023_/a_27_47# 0
C45240 clknet_1_0__leaf__0462_ _0345_ 0.11718f
C45241 clkbuf_0__0463_/a_110_47# _0913_/a_27_47# 0
C45242 _0555_/a_512_297# net26 0
C45243 _0389_ _0244_ 0.00243f
C45244 VPWR _0176_ 1.97237f
C45245 hold64/a_49_47# _0181_ 0
C45246 _0113_ comp0.B\[15\] 0.0013f
C45247 _0172_ _0085_ 0.07596f
C45248 _1002_/a_1017_47# net1 0.0012f
C45249 _1003_/a_1059_315# net51 0
C45250 VPWR _0600_/a_253_47# 0.00165f
C45251 _1057_/a_466_413# net2 0
C45252 _1038_/a_634_159# net8 0
C45253 _1039_/a_891_413# _0473_ 0.00361f
C45254 _0625_/a_59_75# net65 0
C45255 _0625_/a_59_75# _0989_/a_466_413# 0
C45256 _0467_ _1072_/a_466_413# 0
C45257 _0201_ clkbuf_1_1__f__0464_/a_110_47# 0
C45258 clkbuf_0__0461_/a_110_47# _0392_ 0.00479f
C45259 _0958_/a_27_47# _0471_ 0.13964f
C45260 _1051_/a_891_413# _0193_ 0
C45261 _0399_ net217 0.00104f
C45262 hold42/a_285_47# net3 0
C45263 _1049_/a_27_47# _1048_/a_27_47# 0.00331f
C45264 _0276_ clkbuf_1_1__f__0459_/a_110_47# 0.02484f
C45265 _0367_ acc0.A\[24\] 0.02864f
C45266 _0224_ _0222_ 0.19767f
C45267 _1058_/a_27_47# output37/a_27_47# 0
C45268 net64 _0829_/a_27_47# 0
C45269 _0461_ _0585_/a_373_47# 0
C45270 _0287_ hold70/a_49_47# 0
C45271 _0289_ hold70/a_285_47# 0.00184f
C45272 hold59/a_391_47# _0347_ 0
C45273 VPWR _1011_/a_891_413# 0.20311f
C45274 hold88/a_285_47# _0190_ 0
C45275 net53 _1024_/a_891_413# 0
C45276 VPWR _1006_/a_27_47# 0.68195f
C45277 _1029_/a_193_47# _1008_/a_193_47# 0.00173f
C45278 _0857_/a_27_47# net23 0
C45279 _0343_ net70 0.01813f
C45280 _0995_/a_193_47# _0400_ 0
C45281 _0751_/a_29_53# VPWR 0.12846f
C45282 net37 hold81/a_49_47# 0
C45283 _0963_/a_285_297# _1069_/a_1059_315# 0
C45284 _1055_/a_27_47# A[10] 0
C45285 _1030_/a_466_413# net57 0
C45286 _0195_ _1030_/a_634_159# 0.02543f
C45287 _0216_ _1030_/a_27_47# 0.02213f
C45288 net48 _1005_/a_634_159# 0.01128f
C45289 _0644_/a_47_47# _0996_/a_891_413# 0
C45290 _0135_ _0207_ 0
C45291 VPWR _0986_/a_27_47# 0.66094f
C45292 input2/a_75_212# net181 0.00109f
C45293 _0287_ _0089_ 0
C45294 _0603_/a_68_297# _0764_/a_81_21# 0.00582f
C45295 _0714_/a_51_297# _0345_ 0.12275f
C45296 hold21/a_49_47# acc0.A\[6\] 0
C45297 _1019_/a_891_413# _0345_ 0.04672f
C45298 output67/a_27_47# _1058_/a_466_413# 0
C45299 net141 _0186_ 0
C45300 _0804_/a_79_21# _0994_/a_193_47# 0
C45301 net67 hold81/a_391_47# 0.01167f
C45302 _1031_/a_27_47# hold62/a_285_47# 0
C45303 _0180_ net157 0.01933f
C45304 _0240_ clknet_1_1__leaf__0461_ 0
C45305 _1012_/a_381_47# _0110_ 0.13795f
C45306 net39 _0403_ 0.0935f
C45307 _0369_ clknet_1_1__leaf__0461_ 0.15625f
C45308 _0217_ acc0.A\[24\] 0.03462f
C45309 _0275_ _0445_ 0.03741f
C45310 _0272_ _0084_ 0
C45311 control0.state\[0\] _0972_/a_250_297# 0.00812f
C45312 control0.state\[1\] _0972_/a_93_21# 0.08592f
C45313 _0218_ _0799_/a_303_47# 0.0013f
C45314 _0216_ net190 0.19598f
C45315 net23 _1062_/a_27_47# 0
C45316 net206 _0345_ 0
C45317 _0140_ net128 0.00918f
C45318 VPWR net130 0.40731f
C45319 _0146_ _1049_/a_891_413# 0
C45320 _0650_/a_150_297# acc0.A\[10\] 0
C45321 clkbuf_1_0__f__0459_/a_110_47# _0157_ 0
C45322 _0957_/a_32_297# _0561_/a_51_297# 0
C45323 net95 _1009_/a_634_159# 0
C45324 _0154_ _0189_ 0.01255f
C45325 comp0.B\[11\] B[11] 0.00267f
C45326 _0080_ _0345_ 0
C45327 control0.count\[3\] _0468_ 0
C45328 _0960_/a_109_47# _0480_ 0
C45329 _0960_/a_27_47# net164 0
C45330 _0175_ _0562_/a_150_297# 0
C45331 _0461_ _0772_/a_215_47# 0.00109f
C45332 _0402_ _0421_ 0.22427f
C45333 _0643_/a_253_47# _0275_ 0.00137f
C45334 _0606_/a_392_297# _0219_ 0
C45335 _0830_/a_79_21# clkbuf_1_0__f__0465_/a_110_47# 0.00153f
C45336 _0601_/a_68_297# _0102_ 0
C45337 _0255_ _0268_ 0
C45338 comp0.B\[8\] _1040_/a_634_159# 0.03593f
C45339 _0206_ _1040_/a_193_47# 0.04976f
C45340 _0516_/a_27_297# net66 0
C45341 _1059_/a_891_413# clknet_1_0__leaf__0459_ 0
C45342 hold76/a_391_47# _0218_ 0
C45343 net25 hold84/a_49_47# 0
C45344 _0172_ clkbuf_0__0463_/a_110_47# 0.00642f
C45345 _0340_ VPWR 0.55923f
C45346 net47 _0988_/a_27_47# 0
C45347 clknet_1_0__leaf__0460_ _0373_ 0
C45348 _0331_ _0352_ 0.00242f
C45349 hold98/a_285_47# net81 0
C45350 clknet_1_0__leaf__0460_ _0758_/a_297_297# 0.00118f
C45351 _0133_ _0957_/a_32_297# 0.00142f
C45352 hold82/a_49_47# net229 0
C45353 VPWR _0845_/a_193_297# 0.00313f
C45354 _0582_/a_27_297# net221 0.13291f
C45355 _0350_ net50 0.10134f
C45356 clknet_1_0__leaf__0458_ VPWR 3.23243f
C45357 _0080_ hold2/a_49_47# 0.09192f
C45358 net68 hold2/a_285_47# 0.00371f
C45359 _0855_/a_299_297# _1014_/a_193_47# 0
C45360 hold23/a_391_47# net71 0
C45361 _1052_/a_634_159# _1052_/a_381_47# 0
C45362 _0478_ _1071_/a_381_47# 0
C45363 _1007_/a_193_47# _1007_/a_891_413# 0.1937f
C45364 _1007_/a_27_47# _1007_/a_381_47# 0.06222f
C45365 _1007_/a_634_159# _1007_/a_1059_315# 0
C45366 _0125_ _0126_ 0.08326f
C45367 _1035_/a_1017_47# _0133_ 0.00125f
C45368 VPWR _0737_/a_35_297# 0.2035f
C45369 _1012_/a_193_47# _1010_/a_381_47# 0
C45370 _1012_/a_381_47# _1010_/a_193_47# 0
C45371 _0967_/a_215_297# net33 0
C45372 hold10/a_285_47# _0177_ 0
C45373 _0243_ _1006_/a_193_47# 0
C45374 _0346_ net146 0
C45375 _0133_ net23 0
C45376 _1012_/a_891_413# acc0.A\[30\] 0
C45377 _0837_/a_81_21# _0837_/a_266_297# 0.01575f
C45378 _1058_/a_634_159# _1058_/a_975_413# 0
C45379 _1058_/a_466_413# _1058_/a_561_413# 0.00772f
C45380 net186 _1034_/a_1059_315# 0
C45381 _0973_/a_109_297# hold93/a_391_47# 0
C45382 _0172_ _1044_/a_193_47# 0.28324f
C45383 _0179_ _1052_/a_193_47# 0.01758f
C45384 _0552_/a_68_297# net28 0
C45385 _0098_ _0240_ 0
C45386 net45 _0247_ 0.64757f
C45387 hold10/a_49_47# _0178_ 0
C45388 _0197_ net247 0
C45389 clknet_1_0__leaf__0462_ hold52/a_285_47# 0.00958f
C45390 _0312_ _0104_ 0
C45391 clkload1/Y net63 0
C45392 _0172_ net131 0.04394f
C45393 net185 _1035_/a_1059_315# 0
C45394 _1050_/a_193_47# net154 0.02762f
C45395 _0558_/a_68_297# net23 0
C45396 _0680_/a_217_297# _0311_ 0.01327f
C45397 VPWR _0722_/a_297_297# 0.01207f
C45398 acc0.A\[12\] _0510_/a_109_47# 0
C45399 _0353_ hold62/a_391_47# 0
C45400 input20/a_75_212# B[12] 0.20097f
C45401 net97 _0726_/a_149_47# 0.00119f
C45402 _1011_/a_466_413# _0109_ 0.03064f
C45403 _1011_/a_381_47# net227 0
C45404 VPWR _1013_/a_381_47# 0.07542f
C45405 _0257_ _0218_ 0.08263f
C45406 _0131_ _1065_/a_193_47# 0
C45407 net166 net102 0.00103f
C45408 net119 _1065_/a_634_159# 0
C45409 _1002_/a_1059_315# VPWR 0.40005f
C45410 input19/a_75_212# net20 0
C45411 _0399_ net66 0.04188f
C45412 acc0.A\[16\] VPWR 0.97255f
C45413 _0143_ clknet_1_0__leaf__0464_ 0.00143f
C45414 _1052_/a_561_413# net12 0
C45415 _0402_ _0809_/a_81_21# 0
C45416 _0329_ _0727_/a_109_47# 0.00869f
C45417 _0259_ _0254_ 0.00685f
C45418 _0742_/a_299_297# acc0.A\[24\] 0.00678f
C45419 _0516_/a_27_297# _0350_ 0
C45420 _0538_/a_149_47# comp0.B\[14\] 0
C45421 _0461_ net17 0
C45422 clknet_1_0__leaf__0462_ net52 0.0422f
C45423 _0312_ _0745_/a_109_47# 0
C45424 net219 _0611_/a_68_297# 0
C45425 _0328_ _1007_/a_891_413# 0
C45426 _1058_/a_193_47# _0186_ 0
C45427 _0179_ net12 0.02228f
C45428 net56 _0356_ 0
C45429 clkbuf_0_clk/a_110_47# _0974_/a_79_199# 0.00659f
C45430 _0327_ _0727_/a_193_47# 0.00924f
C45431 _0555_/a_51_297# _0549_/a_68_297# 0
C45432 _0346_ net223 0
C45433 net65 pp[3] 0.00662f
C45434 net217 _0295_ 0
C45435 _0399_ _0991_/a_27_47# 0
C45436 _0788_/a_68_297# _0788_/a_150_297# 0.00477f
C45437 _0422_ _0296_ 0
C45438 _0218_ clknet_1_1__leaf__0462_ 0
C45439 pp[30] net60 0
C45440 _1038_/a_592_47# _0176_ 0
C45441 _0359_ acc0.A\[23\] 0
C45442 hold70/a_285_47# _0418_ 0
C45443 clknet_0_clk _0950_/a_75_212# 0.00843f
C45444 VPWR _0525_/a_299_297# 0.27463f
C45445 _0974_/a_544_297# _0974_/a_448_47# 0.00203f
C45446 _0536_/a_51_297# clkbuf_0__0464_/a_110_47# 0
C45447 _0984_/a_1059_315# VPWR 0.39446f
C45448 _0172_ _0546_/a_512_297# 0.00116f
C45449 _0550_/a_149_47# net32 0
C45450 _0746_/a_384_47# _0359_ 0.0094f
C45451 _0994_/a_381_47# _0218_ 0.00939f
C45452 _0495_/a_68_297# _0175_ 0.10679f
C45453 output63/a_27_47# pp[5] 0.33669f
C45454 net44 _0704_/a_68_297# 0
C45455 net138 _1052_/a_27_47# 0.22281f
C45456 clkbuf_1_0__f__0464_/a_110_47# _0527_/a_27_297# 0
C45457 pp[27] net44 0
C45458 net67 _0281_ 0.02968f
C45459 _0995_/a_592_47# pp[14] 0
C45460 hold13/a_391_47# _1039_/a_1059_315# 0
C45461 net211 net105 0
C45462 net111 _1026_/a_1059_315# 0
C45463 _0183_ _0117_ 0.1359f
C45464 _0093_ _0400_ 0
C45465 _0570_/a_27_297# _1026_/a_891_413# 0
C45466 _0570_/a_109_297# _1026_/a_1059_315# 0
C45467 _0369_ _0990_/a_193_47# 0
C45468 _0217_ _0583_/a_109_297# 0.01131f
C45469 net183 _0174_ 0.10746f
C45470 clkbuf_1_0__f__0462_/a_110_47# _1007_/a_634_159# 0.01083f
C45471 _0251_ _0642_/a_298_297# 0.00473f
C45472 _1002_/a_1059_315# net48 0.09055f
C45473 _0429_ _0642_/a_27_413# 0.00902f
C45474 VPWR _1042_/a_975_413# 0.00433f
C45475 _0343_ _0795_/a_384_47# 0
C45476 net61 _0087_ 0
C45477 _1056_/a_381_47# acc0.A\[9\] 0.0022f
C45478 net198 _0540_/a_51_297# 0
C45479 _0982_/a_891_413# _0346_ 0
C45480 _1070_/a_27_47# _0979_/a_27_297# 0.02456f
C45481 _0518_/a_373_47# _0252_ 0
C45482 hold98/a_391_47# _0797_/a_27_413# 0
C45483 _0216_ _0855_/a_81_21# 0
C45484 _0195_ _0855_/a_384_47# 0
C45485 control0.sh _0495_/a_150_297# 0
C45486 _0691_/a_150_297# _0315_ 0
C45487 _0783_/a_510_47# clknet_0__0461_ 0
C45488 _0578_/a_27_297# _0462_ 0
C45489 output54/a_27_47# _0216_ 0.00344f
C45490 _0399_ _0350_ 0.89903f
C45491 net179 net74 0
C45492 _0181_ net134 0
C45493 _1030_/a_891_413# acc0.A\[30\] 0.04133f
C45494 _0273_ net65 0
C45495 _0273_ _0989_/a_466_413# 0
C45496 _0343_ hold31/a_49_47# 0
C45497 _0988_/a_1059_315# _0988_/a_891_413# 0.31086f
C45498 _0988_/a_193_47# _0988_/a_975_413# 0
C45499 _0988_/a_466_413# _0988_/a_381_47# 0.03733f
C45500 _0553_/a_51_297# _0553_/a_245_297# 0.01218f
C45501 _0314_ _0462_ 0
C45502 _0352_ _0377_ 0.03393f
C45503 _0459_ net47 0
C45504 _1053_/a_27_47# acc0.A\[7\] 0.00387f
C45505 hold60/a_49_47# _0099_ 0
C45506 clkbuf_0_clk/a_110_47# _1062_/a_193_47# 0
C45507 _0280_ _0301_ 0.13786f
C45508 _0217_ _0610_/a_59_75# 0
C45509 VPWR _0532_/a_299_297# 0.24225f
C45510 _0982_/a_27_47# _0465_ 0.00198f
C45511 _1020_/a_891_413# clkbuf_0__0457_/a_110_47# 0
C45512 _0343_ net243 0
C45513 _0111_ _1031_/a_27_47# 0
C45514 net225 _1031_/a_634_159# 0
C45515 _0181_ _0084_ 0
C45516 _0354_ _0334_ 0.08543f
C45517 _0542_/a_51_297# net195 0.0804f
C45518 _0621_/a_35_297# _0399_ 0
C45519 _1056_/a_193_47# _0369_ 0
C45520 _0399_ net80 0
C45521 A[13] _0994_/a_1059_315# 0
C45522 hold38/a_285_47# net231 0
C45523 _0982_/a_891_413# _0629_/a_59_75# 0
C45524 _0443_ _0840_/a_68_297# 0.01635f
C45525 clkload1/a_110_47# clknet_1_0__leaf__0465_ 0
C45526 _1001_/a_891_413# clknet_1_0__leaf__0457_ 0.01951f
C45527 _0465_ _0145_ 0.01711f
C45528 B[10] net18 0.0079f
C45529 _0999_/a_381_47# _0396_ 0.00142f
C45530 _0999_/a_1059_315# _0097_ 0.00111f
C45531 net89 _0973_/a_27_297# 0
C45532 _0460_ _1062_/a_634_159# 0
C45533 clknet_1_0__leaf__0457_ _1062_/a_1059_315# 0
C45534 _1021_/a_27_47# _0460_ 0.00977f
C45535 _1021_/a_634_159# clknet_1_0__leaf__0457_ 0.00578f
C45536 _1035_/a_891_413# net27 0.01232f
C45537 _0490_ _0484_ 0.00368f
C45538 _0316_ _1008_/a_466_413# 0
C45539 _0179_ acc0.A\[10\] 0.23622f
C45540 _0343_ output60/a_27_47# 0.00267f
C45541 _0244_ _0612_/a_59_75# 0.11044f
C45542 net133 _1047_/a_27_47# 0.23589f
C45543 _0769_/a_81_21# acc0.A\[18\] 0
C45544 input23/a_75_212# B[4] 0.04076f
C45545 B[15] input27/a_75_212# 0
C45546 hold22/a_285_47# _0180_ 0.00125f
C45547 _0831_/a_35_297# _0186_ 0
C45548 _0982_/a_381_47# hold60/a_391_47# 0
C45549 net54 _0125_ 0.23851f
C45550 _0429_ _0218_ 0
C45551 comp0.B\[9\] _1040_/a_1059_315# 0.00186f
C45552 hold48/a_49_47# _0141_ 0
C45553 _0626_/a_68_297# _0270_ 0
C45554 hold87/a_49_47# acc0.A\[18\] 0
C45555 _0302_ net5 0
C45556 net178 hold32/a_285_47# 0
C45557 net194 net154 0
C45558 _1059_/a_1059_315# _0673_/a_103_199# 0
C45559 _0279_ _0994_/a_1059_315# 0
C45560 _0795_/a_299_297# net5 0.00848f
C45561 _0461_ _0245_ 0.02496f
C45562 _0405_ _0345_ 0.16063f
C45563 _0792_/a_209_47# _0219_ 0.0037f
C45564 _0557_/a_51_297# _0175_ 0.11156f
C45565 _0311_ _0372_ 0.00218f
C45566 net43 acc0.A\[15\] 0.00358f
C45567 _0347_ _1008_/a_466_413# 0.01442f
C45568 _0378_ _0755_/a_109_297# 0.01129f
C45569 _1037_/a_1059_315# _0135_ 0.04861f
C45570 _0745_/a_193_47# _0219_ 0
C45571 _0531_/a_109_297# _1048_/a_193_47# 0
C45572 _0531_/a_27_297# _1048_/a_634_159# 0
C45573 _0996_/a_27_47# hold91/a_49_47# 0
C45574 hold97/a_49_47# clkbuf_1_1__f__0462_/a_110_47# 0
C45575 _0195_ _0998_/a_975_413# 0
C45576 _0356_ _0345_ 0.03378f
C45577 hold38/a_49_47# hold38/a_391_47# 0.00188f
C45578 _0171_ _0492_/a_27_47# 0.16459f
C45579 clknet_1_0__leaf__0462_ _0576_/a_109_47# 0.00105f
C45580 _0465_ _0446_ 0.04383f
C45581 pp[30] _1030_/a_561_413# 0
C45582 hold34/a_49_47# hold34/a_285_47# 0.22264f
C45583 _0557_/a_245_297# control0.sh 0.00216f
C45584 net47 _0265_ 0.13524f
C45585 net60 _0339_ 0.00373f
C45586 VPWR net91 0.46759f
C45587 _0513_/a_81_21# acc0.A\[10\] 0
C45588 acc0.A\[2\] _0446_ 0.00304f
C45589 _0999_/a_193_47# net42 0
C45590 _0207_ _0206_ 0
C45591 output56/a_27_47# VPWR 0.24443f
C45592 VPWR hold91/a_285_47# 0.29293f
C45593 _0985_/a_1059_315# _0448_ 0
C45594 hold18/a_49_47# VPWR 0.29728f
C45595 net234 _0454_ 0
C45596 _0959_/a_300_47# net23 0.00293f
C45597 _0218_ _0668_/a_382_297# 0
C45598 _1001_/a_466_413# _1001_/a_381_47# 0.03733f
C45599 _1001_/a_193_47# _1001_/a_975_413# 0
C45600 _1001_/a_1059_315# _1001_/a_891_413# 0.31086f
C45601 _0422_ _0811_/a_81_21# 0.11556f
C45602 _0855_/a_81_21# net247 0
C45603 acc0.A\[16\] clknet_1_0__leaf__0459_ 0.5304f
C45604 net189 net2 0.0044f
C45605 net124 net8 0.16698f
C45606 _0174_ _0957_/a_32_297# 0
C45607 _1062_/a_193_47# _1062_/a_381_47# 0.09799f
C45608 _1062_/a_634_159# _1062_/a_891_413# 0.03684f
C45609 _1062_/a_27_47# _1062_/a_561_413# 0.0027f
C45610 _0179_ pp[5] 0
C45611 _0342_ _0567_/a_27_297# 0.11408f
C45612 clknet_1_0__leaf__0458_ _0453_ 0.0059f
C45613 _1011_/a_466_413# _0725_/a_80_21# 0.00311f
C45614 _0992_/a_27_47# net228 0
C45615 _0477_ _0471_ 0.00145f
C45616 _0472_ _0953_/a_304_297# 0
C45617 _1021_/a_193_47# _1021_/a_634_159# 0.12126f
C45618 _1021_/a_27_47# _1021_/a_466_413# 0.27314f
C45619 _0831_/a_117_297# _0253_ 0
C45620 _1003_/a_466_413# net49 0
C45621 net44 _0216_ 0.02747f
C45622 pp[17] _0195_ 0
C45623 hold41/a_285_47# hold41/a_391_47# 0.41909f
C45624 _0481_ _0977_/a_75_212# 0.00112f
C45625 _0430_ _0827_/a_109_297# 0
C45626 _0091_ _0807_/a_68_297# 0
C45627 _0430_ _0255_ 0.00847f
C45628 hold14/a_285_47# _1037_/a_381_47# 0
C45629 _0642_/a_27_413# clknet_1_1__leaf__0458_ 0
C45630 net78 _0345_ 0.00151f
C45631 control0.state\[0\] _0971_/a_81_21# 0.00271f
C45632 _0254_ _0253_ 0.08829f
C45633 net141 net62 0.00139f
C45634 comp0.B\[14\] clkbuf_0__0464_/a_110_47# 0.0037f
C45635 hold15/a_49_47# _0708_/a_68_297# 0
C45636 _0271_ _0434_ 0
C45637 clknet_0__0465_ _0345_ 0.0011f
C45638 _0459_ _1060_/a_1059_315# 0.02639f
C45639 VPWR _0288_ 0.99391f
C45640 net115 _1008_/a_27_47# 0
C45641 _1029_/a_27_47# net94 0
C45642 _1000_/a_1059_315# _0183_ 0
C45643 _0267_ _0261_ 0
C45644 _0586_/a_27_47# clknet_1_0__leaf__0457_ 0.00213f
C45645 _0963_/a_35_297# control0.count\[0\] 0.2062f
C45646 hold88/a_285_47# _0346_ 0
C45647 hold47/a_391_47# _0143_ 0.00192f
C45648 _0839_/a_109_297# _0399_ 0
C45649 acc0.A\[5\] _0255_ 0.54882f
C45650 _0241_ _0869_/a_27_47# 0
C45651 _0107_ _0350_ 0.112f
C45652 _0856_/a_297_297# VPWR 0.00839f
C45653 clknet_1_1__leaf__0463_ _0494_/a_27_47# 0
C45654 control0.state\[0\] _0975_/a_145_75# 0.00257f
C45655 control0.state\[1\] _0975_/a_59_75# 0.00236f
C45656 net48 net91 0.00236f
C45657 _0826_/a_27_53# _0431_ 0
C45658 clknet_1_1__leaf__0464_ _1043_/a_466_413# 0.03867f
C45659 _0195_ _1015_/a_193_47# 0
C45660 _0749_/a_299_297# acc0.A\[19\] 0
C45661 clknet_1_1__leaf__0459_ _0795_/a_81_21# 0
C45662 net30 _0176_ 0.01588f
C45663 net157 _0498_/a_51_297# 0.00143f
C45664 net225 _0345_ 0
C45665 _0083_ _0846_/a_512_297# 0
C45666 net45 _0779_/a_297_297# 0
C45667 _0585_/a_27_297# clknet_1_0__leaf__0461_ 0
C45668 VPWR _0670_/a_215_47# 0.00535f
C45669 _1034_/a_27_47# clkbuf_1_1__f__0463_/a_110_47# 0.01321f
C45670 net5 net6 0.02018f
C45671 _0092_ _0994_/a_634_159# 0
C45672 hold55/a_285_47# _0461_ 0.00111f
C45673 _1020_/a_634_159# _0721_/a_27_47# 0.00838f
C45674 _0951_/a_209_311# comp0.B\[0\] 0.23039f
C45675 A[12] net67 0.00607f
C45676 _0225_ _1022_/a_27_47# 0
C45677 _0224_ _1022_/a_466_413# 0
C45678 _0714_/a_245_297# _0344_ 0.0019f
C45679 _0438_ _0369_ 0.01632f
C45680 control0.state\[0\] _0164_ 0.00522f
C45681 _0561_/a_149_47# _0561_/a_240_47# 0.06872f
C45682 _0561_/a_51_297# _0213_ 0.10481f
C45683 control0.state\[1\] net231 0.22051f
C45684 VPWR _0247_ 0.63833f
C45685 net8 _0494_/a_27_47# 0
C45686 _0219_ hold95/a_285_47# 0
C45687 clkbuf_1_0__f__0457_/a_110_47# VPWR 1.45072f
C45688 _0180_ net13 0.12645f
C45689 hold13/a_391_47# _1037_/a_1059_315# 0
C45690 net39 acc0.A\[13\] 0
C45691 net181 _0514_/a_27_297# 0
C45692 _0221_ hold62/a_49_47# 0
C45693 output44/a_27_47# _0338_ 0
C45694 clknet_0__0461_ acc0.A\[18\] 0.18263f
C45695 _0179_ _0510_/a_109_297# 0
C45696 hold41/a_49_47# _0181_ 0.0023f
C45697 comp0.B\[13\] net183 0.00486f
C45698 net193 _0201_ 0
C45699 _0957_/a_32_297# _0208_ 0.01137f
C45700 _0957_/a_304_297# _0173_ 0
C45701 _0252_ net235 0
C45702 net65 _0086_ 0
C45703 _1036_/a_1059_315# clknet_1_1__leaf__0463_ 0.01808f
C45704 _1036_/a_634_159# net122 0
C45705 _0226_ _0346_ 0.02346f
C45706 _1052_/a_193_47# hold83/a_49_47# 0.00284f
C45707 _1052_/a_27_47# hold83/a_285_47# 0
C45708 _1050_/a_193_47# clknet_0__0464_ 0
C45709 _0343_ _0366_ 0.00255f
C45710 _0738_/a_150_297# net244 0
C45711 _0461_ _1019_/a_634_159# 0.00407f
C45712 net89 acc0.A\[21\] 0
C45713 _0218_ clknet_1_1__leaf__0458_ 0.01116f
C45714 pp[9] _0186_ 0.01063f
C45715 _0749_/a_299_297# _0249_ 0
C45716 net121 _0173_ 0.00203f
C45717 _0133_ _0213_ 0.59332f
C45718 _1035_/a_1017_47# _0208_ 0
C45719 hold67/a_49_47# hold67/a_391_47# 0.00188f
C45720 _1041_/a_634_159# net153 0.00898f
C45721 _1041_/a_466_413# net127 0
C45722 _1047_/a_634_159# _1047_/a_592_47# 0
C45723 net23 _0208_ 0.02724f
C45724 _1030_/a_561_413# _0339_ 0
C45725 _0307_ _0675_/a_68_297# 0.12296f
C45726 _0190_ net66 0
C45727 _0305_ _0780_/a_117_297# 0.002f
C45728 _0473_ _0475_ 0.13652f
C45729 hold39/a_391_47# clknet_1_1__leaf_clk 0
C45730 _0714_/a_240_47# net163 0
C45731 control0.state\[1\] hold38/a_285_47# 0
C45732 _0131_ _0563_/a_149_47# 0.02989f
C45733 comp0.B\[1\] _0563_/a_51_297# 0
C45734 _1041_/a_891_413# _0136_ 0
C45735 net185 _0561_/a_245_297# 0.0019f
C45736 input9/a_27_47# input18/a_75_212# 0
C45737 _0212_ _0561_/a_51_297# 0.00309f
C45738 _0226_ hold94/a_49_47# 0
C45739 net221 _0115_ 0.05714f
C45740 _0343_ _0718_/a_377_297# 0
C45741 _0474_ _0496_/a_27_47# 0
C45742 _0216_ _0566_/a_27_47# 0.3674f
C45743 acc0.A\[7\] A[5] 0
C45744 _0217_ _1018_/a_466_413# 0.00332f
C45745 _0183_ _1018_/a_193_47# 0
C45746 _0456_ _1014_/a_891_413# 0
C45747 _0855_/a_81_21# net100 0
C45748 _0354_ _0724_/a_113_297# 0.09503f
C45749 _1007_/a_466_413# _0105_ 0.00388f
C45750 net243 _1004_/a_466_413# 0.00217f
C45751 VPWR _0455_ 0.19347f
C45752 net12 hold83/a_49_47# 0.01492f
C45753 _0837_/a_266_47# _0441_ 0.04052f
C45754 _0443_ _0255_ 0.18134f
C45755 net168 _0518_/a_27_297# 0
C45756 _0502_/a_27_47# acc0.A\[1\] 0
C45757 _1020_/a_592_47# _0352_ 0
C45758 _0126_ _1027_/a_634_159# 0
C45759 net190 _1027_/a_891_413# 0
C45760 _0848_/a_27_47# _0263_ 0
C45761 net48 _0762_/a_510_47# 0
C45762 _0667_/a_113_47# net40 0
C45763 clkbuf_1_0__f__0457_/a_110_47# net48 0.00185f
C45764 hold7/a_49_47# _0987_/a_27_47# 0.01011f
C45765 _0397_ _0097_ 0
C45766 hold98/a_49_47# acc0.A\[31\] 0
C45767 _0218_ _0263_ 0.04493f
C45768 _0212_ _0133_ 0.02588f
C45769 _0234_ hold66/a_285_47# 0.00171f
C45770 _0268_ _0843_/a_68_297# 0.11941f
C45771 _0267_ net47 0
C45772 _0850_/a_68_297# _0850_/a_150_297# 0.00477f
C45773 hold32/a_391_47# pp[1] 0
C45774 acc0.A\[4\] _0346_ 0
C45775 _0266_ _1014_/a_27_47# 0
C45776 net44 _0608_/a_109_297# 0.01111f
C45777 comp0.B\[11\] _0140_ 0.19911f
C45778 net57 net227 0.24511f
C45779 VPWR _0505_/a_109_297# 0.19311f
C45780 clknet_1_1__leaf__0460_ _0332_ 0.00431f
C45781 _0558_/a_68_297# _0212_ 0.10608f
C45782 _1061_/a_561_413# comp0.B\[9\] 0
C45783 _0346_ clkbuf_0__0457_/a_110_47# 0.01424f
C45784 _1057_/a_193_47# net67 0.0287f
C45785 net61 _0989_/a_975_413# 0
C45786 _0780_/a_35_297# net43 0
C45787 _0286_ net37 0.00239f
C45788 _0983_/a_1059_315# _0081_ 0
C45789 _0983_/a_381_47# _0455_ 0
C45790 _0190_ _0350_ 0
C45791 pp[2] _0434_ 0.00507f
C45792 _1059_/a_975_413# _0277_ 0
C45793 clknet_1_1__leaf__0460_ _0685_/a_68_297# 0.00293f
C45794 _1063_/a_466_413# _1063_/a_561_413# 0.00772f
C45795 _1063_/a_634_159# _1063_/a_975_413# 0
C45796 input13/a_75_212# net12 0
C45797 _0833_/a_79_21# _0988_/a_193_47# 0
C45798 _0390_ clkbuf_1_0__f__0457_/a_110_47# 0.00108f
C45799 hold58/a_49_47# control0.sh 0.02671f
C45800 _0477_ control0.reset 0
C45801 control0.state\[2\] _0486_ 0.24386f
C45802 _0965_/a_47_47# _1072_/a_193_47# 0
C45803 net61 _0465_ 0.01289f
C45804 clknet_1_1__leaf__0459_ net99 0.00241f
C45805 _1019_/a_561_413# _0346_ 0
C45806 _0179_ _0188_ 0.35482f
C45807 hold75/a_285_47# clknet_1_0__leaf__0458_ 0.00187f
C45808 _0305_ _0507_/a_27_297# 0.0143f
C45809 _0405_ _0791_/a_113_297# 0.1179f
C45810 _0959_/a_80_21# _0959_/a_472_297# 0.01636f
C45811 _0294_ _0459_ 0.03057f
C45812 acc0.A\[20\] _0391_ 0.00202f
C45813 _0462_ _1006_/a_381_47# 0.00104f
C45814 net61 acc0.A\[2\] 0
C45815 net46 _1022_/a_1059_315# 0.00117f
C45816 clknet_1_0__leaf__0464_ _1050_/a_27_47# 0.00943f
C45817 _0748_/a_299_297# _0748_/a_384_47# 0
C45818 net149 clknet_1_0__leaf__0457_ 0
C45819 _0544_/a_51_297# _0203_ 0
C45820 _0716_/a_27_47# _0305_ 0
C45821 _0204_ _0542_/a_51_297# 0
C45822 net205 comp0.B\[2\] 0.01582f
C45823 _0343_ _0790_/a_285_47# 0
C45824 _1028_/a_193_47# net113 0
C45825 _1028_/a_466_413# clknet_1_1__leaf__0462_ 0.02155f
C45826 hold11/a_391_47# net135 0
C45827 hold11/a_285_47# _0147_ 0
C45828 _0663_/a_297_47# _0345_ 0
C45829 _0172_ _0139_ 0.27065f
C45830 VPWR _0506_/a_299_297# 0.21647f
C45831 net15 net11 0.00515f
C45832 control0.count\[3\] _1071_/a_466_413# 0
C45833 _0483_ _1071_/a_193_47# 0
C45834 _0369_ clknet_1_1__leaf__0465_ 0.2625f
C45835 _0733_/a_222_93# _0368_ 0
C45836 _0251_ _0191_ 0
C45837 _0346_ _0807_/a_68_297# 0
C45838 _0819_/a_81_21# clknet_0__0465_ 0.05336f
C45839 hold47/a_49_47# _0186_ 0.00311f
C45840 net167 _0482_ 0
C45841 _0515_/a_299_297# net66 0.01022f
C45842 _0238_ acc0.A\[23\] 0
C45843 _1011_/a_1017_47# acc0.A\[29\] 0
C45844 _0833_/a_215_47# clknet_1_1__leaf__0458_ 0
C45845 _0195_ _0569_/a_27_297# 0.16421f
C45846 hold18/a_391_47# _0266_ 0
C45847 hold101/a_285_47# _0835_/a_78_199# 0.01622f
C45848 net16 _0290_ 0
C45849 VPWR _1010_/a_466_413# 0.26758f
C45850 clkbuf_1_0__f__0462_/a_110_47# net93 0
C45851 _1000_/a_193_47# _1000_/a_634_159# 0.11715f
C45852 _1000_/a_27_47# _1000_/a_466_413# 0.26957f
C45853 net18 net20 0.02161f
C45854 _1060_/a_466_413# _1060_/a_561_413# 0.00772f
C45855 _1060_/a_634_159# _1060_/a_975_413# 0
C45856 _0251_ output58/a_27_47# 0
C45857 _0204_ _0142_ 0
C45858 _0140_ _0202_ 0
C45859 _0513_/a_81_21# _0188_ 0.1825f
C45860 _1051_/a_1059_315# _0527_/a_27_297# 0
C45861 acc0.A\[28\] _1008_/a_193_47# 0
C45862 _0218_ clknet_1_0__leaf__0461_ 0.42349f
C45863 _1070_/a_27_47# _0169_ 0
C45864 hold48/a_285_47# net18 0.00164f
C45865 hold49/a_285_47# hold49/a_391_47# 0.41909f
C45866 _0192_ _0520_/a_109_297# 0.00169f
C45867 net230 _0520_/a_27_297# 0.16269f
C45868 _0462_ _0616_/a_292_297# 0
C45869 _1053_/a_1059_315# net11 0.01442f
C45870 _1039_/a_561_413# comp0.B\[9\] 0
C45871 net194 clknet_0__0464_ 0.26311f
C45872 _0288_ _0283_ 0
C45873 hold69/a_391_47# clkbuf_0__0460_/a_110_47# 0
C45874 net122 comp0.B\[5\] 0
C45875 VPWR _0846_/a_245_297# 0.00558f
C45876 hold26/a_391_47# _0176_ 0.01314f
C45877 _0467_ _0181_ 0.09375f
C45878 _0553_/a_240_47# _0174_ 0.01664f
C45879 _1067_/a_381_47# clknet_1_1__leaf_clk 0.00142f
C45880 _0399_ _0986_/a_634_159# 0.017f
C45881 clknet_1_0__leaf__0459_ _0247_ 0.03142f
C45882 _0352_ _0688_/a_109_297# 0.00516f
C45883 pp[29] _0109_ 0.00285f
C45884 _0973_/a_109_297# _1063_/a_193_47# 0
C45885 _0322_ _0350_ 0
C45886 net53 _0682_/a_68_297# 0.13022f
C45887 control0.state\[0\] net34 0.75519f
C45888 acc0.A\[27\] clkbuf_0__0462_/a_110_47# 0.00457f
C45889 VPWR _1009_/a_1059_315# 0.40205f
C45890 _0303_ _0302_ 0.19175f
C45891 _0579_/a_109_47# net187 0
C45892 _0172_ _0525_/a_81_21# 0
C45893 clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0459_ 0
C45894 hold19/a_285_47# hold19/a_391_47# 0.41909f
C45895 _0582_/a_27_297# _0245_ 0
C45896 _0327_ _0350_ 0.04434f
C45897 _0235_ _0603_/a_150_297# 0
C45898 _0423_ _0811_/a_81_21# 0
C45899 _0195_ _0266_ 0.0032f
C45900 _0343_ _0378_ 0.00151f
C45901 _0234_ _0183_ 0
C45902 _0161_ _1062_/a_27_47# 0
C45903 net55 clknet_1_1__leaf__0462_ 0.01979f
C45904 _1071_/a_193_47# control0.count\[1\] 0
C45905 _1071_/a_381_47# VPWR 0.07645f
C45906 _0973_/a_109_297# _0460_ 0.00476f
C45907 _1001_/a_1059_315# net149 0
C45908 _0191_ hold7/a_49_47# 0
C45909 _0195_ _0567_/a_109_297# 0.01586f
C45910 clknet_1_0__leaf__0465_ _0434_ 0
C45911 _0985_/a_634_159# _0179_ 0.0206f
C45912 net58 output58/a_27_47# 0.23927f
C45913 _0984_/a_1059_315# hold75/a_285_47# 0.0054f
C45914 _0464_ net10 0.03157f
C45915 _0181_ comp0.B\[0\] 0
C45916 _0346_ net41 0.31874f
C45917 _0592_/a_68_297# net50 0.10426f
C45918 _0780_/a_117_297# _0181_ 0.00181f
C45919 _1059_/a_193_47# _0219_ 0
C45920 _0515_/a_299_297# _0350_ 0
C45921 _0701_/a_80_21# _0333_ 0.07731f
C45922 _0573_/a_27_47# _1015_/a_193_47# 0
C45923 _0462_ _0360_ 0
C45924 clkbuf_0__0462_/a_110_47# _0364_ 0
C45925 VPWR pp[13] 0.2642f
C45926 clknet_0__0464_ _1046_/a_634_159# 0.04256f
C45927 clknet_1_1__leaf__0460_ _0738_/a_68_297# 0.05722f
C45928 _1071_/a_634_159# clkbuf_1_0__f_clk/a_110_47# 0.00695f
C45929 net226 _0167_ 0
C45930 pp[26] _1027_/a_27_47# 0
C45931 net54 _1027_/a_634_159# 0.01084f
C45932 _1008_/a_891_413# _0365_ 0
C45933 _1008_/a_466_413# _0106_ 0.0405f
C45934 _0177_ _1047_/a_27_47# 0
C45935 VPWR _0954_/a_114_297# 0.01788f
C45936 net185 input27/a_75_212# 0
C45937 _0337_ _1030_/a_27_47# 0
C45938 _0314_ _0312_ 0
C45939 hold89/a_49_47# _0471_ 0
C45940 comp0.B\[12\] _1043_/a_193_47# 0
C45941 comp0.B\[11\] _1043_/a_634_159# 0
C45942 VPWR net28 1.09682f
C45943 _0346_ net217 0
C45944 _0343_ net162 0.24535f
C45945 _1020_/a_27_47# _0578_/a_109_297# 0
C45946 _1020_/a_193_47# _0578_/a_27_297# 0
C45947 _1000_/a_27_47# _1018_/a_27_47# 0
C45948 _0276_ _0277_ 0.56613f
C45949 _0201_ _1045_/a_193_47# 0
C45950 _0998_/a_1059_315# _0790_/a_35_297# 0
C45951 net149 _1047_/a_891_413# 0.01339f
C45952 clknet_1_0__leaf__0465_ _0527_/a_109_47# 0
C45953 hold13/a_285_47# _0475_ 0
C45954 VPWR _1022_/a_891_413# 0.18846f
C45955 clkbuf_0_clk/a_110_47# net17 0
C45956 pp[30] _0568_/a_109_297# 0.00149f
C45957 _0133_ _0161_ 0
C45958 _1034_/a_27_47# _0163_ 0
C45959 pp[1] _0153_ 0
C45960 clkload2/Y _0464_ 0
C45961 VPWR _0779_/a_297_297# 0.00963f
C45962 _0553_/a_240_47# _0208_ 0.02334f
C45963 clknet_1_1__leaf__0459_ _0993_/a_1059_315# 0
C45964 _0285_ _0218_ 0.0016f
C45965 _0852_/a_35_297# _0266_ 0.00618f
C45966 _0174_ _0213_ 0.00134f
C45967 _0993_/a_381_47# net38 0
C45968 B[14] hold6/a_49_47# 0
C45969 _0999_/a_634_159# _0999_/a_1059_315# 0
C45970 _0999_/a_27_47# _0999_/a_381_47# 0.05658f
C45971 _0999_/a_193_47# _0999_/a_891_413# 0.19489f
C45972 net17 _1063_/a_634_159# 0.03812f
C45973 _0992_/a_27_47# _0090_ 0.12794f
C45974 _0992_/a_634_159# _0422_ 0
C45975 _1017_/a_27_47# _0115_ 0.07889f
C45976 _1017_/a_891_413# net221 0
C45977 _0972_/a_93_21# clknet_1_1__leaf_clk 0.06484f
C45978 _0330_ _0319_ 0.00911f
C45979 clknet_1_0__leaf__0465_ acc0.A\[7\] 0
C45980 hold26/a_49_47# clkbuf_1_0__f__0463_/a_110_47# 0
C45981 _1001_/a_634_159# net223 0
C45982 _0340_ _1031_/a_634_159# 0
C45983 _0341_ _1031_/a_466_413# 0
C45984 _1001_/a_193_47# _0391_ 0.00185f
C45985 clknet_1_0__leaf__0465_ _0989_/a_1059_315# 0
C45986 _0385_ _0902_/a_27_47# 0
C45987 _1004_/a_193_47# _0217_ 0
C45988 net120 _1034_/a_1059_315# 0
C45989 _0850_/a_68_297# net149 0
C45990 acc0.A\[12\] _0651_/a_113_47# 0
C45991 hold86/a_391_47# _0263_ 0
C45992 _0136_ _0473_ 0
C45993 control0.count\[3\] _0978_/a_109_297# 0
C45994 _1062_/a_1059_315# _0160_ 0
C45995 clknet_0__0458_ _0622_/a_193_47# 0
C45996 B[15] B[2] 0.45189f
C45997 net55 net242 0.08603f
C45998 _1020_/a_27_47# net202 0.05039f
C45999 _0118_ _1032_/a_27_47# 0
C46000 hold87/a_285_47# _0611_/a_68_297# 0
C46001 net132 net154 0
C46002 clkbuf_1_1__f__0459_/a_110_47# _0409_ 0
C46003 _0232_ _0754_/a_51_297# 0
C46004 _0634_/a_113_47# net206 0
C46005 _0343_ acc0.A\[24\] 0
C46006 clknet_1_0__leaf__0465_ _1061_/a_634_159# 0.00373f
C46007 _1021_/a_1059_315# _1021_/a_1017_47# 0
C46008 _1021_/a_27_47# _0119_ 0.11161f
C46009 _0101_ net49 0.20911f
C46010 _0181_ _0507_/a_27_297# 0.15479f
C46011 hold24/a_391_47# _1038_/a_891_413# 0.00406f
C46012 _0575_/a_109_47# _0122_ 0
C46013 net15 clknet_1_1__leaf__0458_ 0
C46014 _0081_ _0266_ 0
C46015 _0455_ _0453_ 0
C46016 _1017_/a_561_413# _0459_ 0
C46017 _0306_ _0350_ 0
C46018 _1049_/a_592_47# net134 0.00121f
C46019 acc0.A\[3\] _1048_/a_891_413# 0
C46020 _0576_/a_27_297# _0350_ 0
C46021 hold41/a_49_47# _0187_ 0
C46022 hold55/a_49_47# net23 0.027f
C46023 _0251_ clkbuf_1_0__f__0465_/a_110_47# 0
C46024 _0174_ _0536_/a_245_297# 0
C46025 _0648_/a_27_297# _0648_/a_109_297# 0.00691f
C46026 VPWR _0540_/a_512_297# 0.00705f
C46027 _0996_/a_634_159# _0302_ 0
C46028 comp0.B\[5\] _0560_/a_150_297# 0
C46029 net45 _0217_ 0.09388f
C46030 _1056_/a_466_413# acc0.A\[12\] 0
C46031 _0369_ _0829_/a_27_47# 0
C46032 net62 _0988_/a_381_47# 0
C46033 _0181_ net165 0.27842f
C46034 _1011_/a_193_47# _0219_ 0.02143f
C46035 _0294_ _1060_/a_381_47# 0
C46036 _1031_/a_466_413# _1013_/a_891_413# 0
C46037 net54 clkbuf_1_1__f__0460_/a_110_47# 0
C46038 clknet_1_1__leaf__0464_ net196 0.11257f
C46039 _0751_/a_29_53# _0345_ 0
C46040 _0376_ _0378_ 0.03643f
C46041 acc0.A\[22\] _0593_/a_113_47# 0
C46042 _0817_/a_266_47# _0426_ 0.03443f
C46043 _0112_ clknet_1_0__leaf__0461_ 0.00999f
C46044 _0168_ _0978_/a_109_47# 0
C46045 _0986_/a_27_47# _0345_ 0
C46046 hold46/a_285_47# _0535_/a_68_297# 0
C46047 clknet_1_0__leaf__0465_ _0538_/a_240_47# 0
C46048 control0.count\[2\] _1071_/a_634_159# 0.03919f
C46049 hold37/a_285_47# _0143_ 0.00662f
C46050 _0467_ _1034_/a_891_413# 0
C46051 _0213_ _0208_ 0.02267f
C46052 VPWR _1067_/a_561_413# 0.00308f
C46053 _0181_ acc0.A\[19\] 0
C46054 _0280_ _0664_/a_79_21# 0
C46055 acc0.A\[12\] _0806_/a_199_47# 0
C46056 _1050_/a_891_413# _0186_ 0
C46057 hold31/a_391_47# VPWR 0.18485f
C46058 _0618_/a_79_21# clkbuf_1_0__f__0460_/a_110_47# 0.01151f
C46059 _1033_/a_891_413# clknet_1_0__leaf__0461_ 0
C46060 net181 _0189_ 0.08837f
C46061 _0227_ _0460_ 0.00125f
C46062 _0276_ _0298_ 0
C46063 net1 _0951_/a_209_311# 0
C46064 _0753_/a_79_21# _0753_/a_297_297# 0.05317f
C46065 hold34/a_49_47# _0153_ 0
C46066 _0618_/a_297_297# _0249_ 0
C46067 _0618_/a_79_21# _0250_ 0.05502f
C46068 _0348_ _1030_/a_975_413# 0
C46069 net180 _0548_/a_51_297# 0.00999f
C46070 hold14/a_391_47# net27 0
C46071 _0461_ net105 0.00848f
C46072 VPWR _1027_/a_193_47# 0.32653f
C46073 _0555_/a_240_47# _1037_/a_1059_315# 0
C46074 _0313_ _0219_ 0.02493f
C46075 _0276_ _0296_ 0
C46076 net160 comp0.B\[2\] 0
C46077 _0640_/a_215_297# _0431_ 0.00107f
C46078 clknet_1_1__leaf__0460_ _0368_ 0.02802f
C46079 _0326_ _0318_ 0.00148f
C46080 _1003_/a_891_413# _0760_/a_285_47# 0
C46081 _1000_/a_193_47# _0242_ 0
C46082 _0997_/a_193_47# _0405_ 0
C46083 hold20/a_391_47# net159 0
C46084 hold46/a_285_47# _0174_ 0.00354f
C46085 _0339_ _0568_/a_109_297# 0
C46086 _0459_ _0581_/a_109_297# 0.0049f
C46087 _0346_ net66 0.00211f
C46088 control0.count\[0\] _0484_ 0
C46089 clknet_1_0__leaf_clk _0162_ 0.08073f
C46090 net157 _1048_/a_891_413# 0
C46091 _0343_ hold74/a_285_47# 0.01182f
C46092 _1042_/a_27_47# hold51/a_49_47# 0
C46093 _0496_/a_27_47# _0563_/a_51_297# 0
C46094 _0212_ _0208_ 0.05372f
C46095 net240 clknet_1_0__leaf__0461_ 0
C46096 net93 net51 0
C46097 _0460_ _0759_/a_113_47# 0
C46098 _0353_ _0334_ 0.05119f
C46099 _0399_ _1014_/a_27_47# 0
C46100 _0546_/a_149_47# _1040_/a_27_47# 0
C46101 _0340_ _0345_ 0.00436f
C46102 net188 _0155_ 0.02909f
C46103 clknet_1_0__leaf__0461_ _0099_ 0
C46104 _1004_/a_27_47# _0379_ 0.00579f
C46105 net190 _0319_ 0
C46106 _0645_/a_47_47# acc0.A\[13\] 0.04746f
C46107 net55 _0730_/a_297_297# 0
C46108 acc0.A\[8\] _0989_/a_634_159# 0.03983f
C46109 acc0.A\[8\] hold1/a_391_47# 0
C46110 _0465_ _0431_ 0.00888f
C46111 pp[17] hold15/a_49_47# 0.02284f
C46112 net44 hold15/a_391_47# 0
C46113 output44/a_27_47# acc0.A\[31\] 0
C46114 _0346_ _0991_/a_27_47# 0.03305f
C46115 clknet_1_0__leaf__0458_ _0345_ 0.05972f
C46116 clkload3/a_268_47# _0181_ 0
C46117 pp[6] _0252_ 0.00213f
C46118 net201 acc0.A\[15\] 0.00174f
C46119 _0996_/a_634_159# net6 0
C46120 _0974_/a_79_199# _0487_ 0.02604f
C46121 _0291_ _0992_/a_193_47# 0
C46122 net168 _0191_ 0.1962f
C46123 _0712_/a_381_47# _0340_ 0.00188f
C46124 clknet_1_0__leaf__0464_ _0987_/a_27_47# 0
C46125 _0217_ net199 0.36863f
C46126 net69 _0852_/a_285_297# 0
C46127 _0387_ _0394_ 0.00509f
C46128 _0544_/a_245_297# _0544_/a_240_47# 0
C46129 _0345_ _0737_/a_35_297# 0.06069f
C46130 net133 _0177_ 0
C46131 _0730_/a_79_21# _0347_ 0.10701f
C46132 _0305_ clkbuf_1_1__f__0461_/a_110_47# 0.00815f
C46133 _0747_/a_215_47# _0460_ 0.00212f
C46134 VPWR _0524_/a_109_47# 0
C46135 _1034_/a_193_47# _1034_/a_381_47# 0.10164f
C46136 _1034_/a_634_159# _1034_/a_891_413# 0.03684f
C46137 _1034_/a_27_47# _1034_/a_561_413# 0.00163f
C46138 hold6/a_49_47# _0544_/a_51_297# 0
C46139 _0796_/a_79_21# _0410_ 0.10751f
C46140 _0796_/a_297_297# net238 0.00222f
C46141 _1021_/a_1059_315# acc0.A\[21\] 0.08405f
C46142 net168 _1053_/a_381_47# 0
C46143 _0960_/a_27_47# _0478_ 0.08831f
C46144 _0305_ _0426_ 0
C46145 VPWR _0972_/a_250_297# 0.30562f
C46146 clknet_1_0__leaf__0458_ hold2/a_49_47# 0.00345f
C46147 _0427_ _0291_ 0.05f
C46148 _0428_ acc0.A\[8\] 0
C46149 hold25/a_49_47# net180 0
C46150 _0982_/a_975_413# clknet_1_0__leaf__0461_ 0
C46151 hold88/a_285_47# _0259_ 0
C46152 _0499_/a_59_75# _0499_/a_145_75# 0.00658f
C46153 _1013_/a_634_159# _0219_ 0
C46154 control0.state\[0\] _1066_/a_466_413# 0
C46155 _0343_ _0583_/a_109_297# 0.0066f
C46156 clknet_0__0464_ _1045_/a_27_47# 0.00465f
C46157 clkbuf_0__0464_/a_110_47# _1045_/a_891_413# 0
C46158 clkbuf_0__0463_/a_110_47# _0214_ 0
C46159 _0086_ _0988_/a_634_159# 0
C46160 _0224_ _0378_ 0.00425f
C46161 _0225_ _0756_/a_285_47# 0.04129f
C46162 VPWR _0448_ 0.14139f
C46163 _0346_ _0350_ 0.75787f
C46164 control0.count\[3\] _0480_ 0
C46165 _0965_/a_285_47# _0169_ 0
C46166 control0.state\[0\] _1068_/a_466_413# 0
C46167 clkbuf_1_0__f__0458_/a_110_47# _0266_ 0
C46168 VPWR _1026_/a_1059_315# 0.40971f
C46169 _0483_ _1072_/a_466_413# 0
C46170 pp[28] acc0.A\[29\] 0.2309f
C46171 control0.count\[3\] _1072_/a_891_413# 0.04267f
C46172 net39 VPWR 1.61614f
C46173 _0225_ _0749_/a_299_297# 0
C46174 hold96/a_49_47# net50 0.30038f
C46175 net35 net49 0.00148f
C46176 net78 _0992_/a_891_413# 0
C46177 _0305_ _0185_ 0.01802f
C46178 VPWR _1024_/a_975_413# 0.00483f
C46179 hold32/a_285_47# hold32/a_391_47# 0.41909f
C46180 _0218_ _0848_/a_27_47# 0.0013f
C46181 output42/a_27_47# _1013_/a_466_413# 0
C46182 _0585_/a_27_297# _0112_ 0.17634f
C46183 _0172_ _0498_/a_240_47# 0.02801f
C46184 VPWR _1048_/a_1017_47# 0
C46185 net34 _0478_ 0
C46186 clknet_1_0__leaf__0460_ _1005_/a_466_413# 0.00427f
C46187 hold52/a_49_47# acc0.A\[25\] 0.07464f
C46188 _0259_ _0086_ 0
C46189 _1017_/a_634_159# _1017_/a_466_413# 0.23992f
C46190 _1017_/a_193_47# _1017_/a_1059_315# 0.03405f
C46191 _1017_/a_27_47# _1017_/a_891_413# 0.03089f
C46192 _0343_ _0610_/a_59_75# 0
C46193 _0487_ _1062_/a_193_47# 0.10429f
C46194 output56/a_27_47# net56 0.17436f
C46195 net86 _0307_ 0.00186f
C46196 _0273_ _0253_ 0.01609f
C46197 hold47/a_285_47# net194 0.00851f
C46198 _0984_/a_27_47# _0219_ 0.00599f
C46199 _0195_ _0127_ 0.00265f
C46200 _0179_ _0531_/a_109_297# 0
C46201 acc0.A\[28\] _0318_ 0
C46202 net117 net163 0.00395f
C46203 _1000_/a_1059_315# _1000_/a_1017_47# 0
C46204 _1000_/a_193_47# net86 0.01548f
C46205 _1000_/a_27_47# _0098_ 0.10109f
C46206 _0507_/a_27_297# _0507_/a_373_47# 0.01338f
C46207 _1006_/a_27_47# net52 0.00795f
C46208 _0629_/a_59_75# _0350_ 0
C46209 _0715_/a_27_47# acc0.A\[8\] 0
C46210 _1056_/a_27_47# hold34/a_49_47# 0
C46211 _0621_/a_35_297# net65 0
C46212 _0430_ _0989_/a_27_47# 0
C46213 _1051_/a_592_47# net154 0
C46214 _0129_ _1013_/a_193_47# 0
C46215 _0195_ _0399_ 0.96965f
C46216 _0168_ net164 0
C46217 _0192_ _0186_ 0
C46218 _0151_ net14 0.02494f
C46219 _0174_ net127 0
C46220 _1072_/a_975_413# VPWR 0.00473f
C46221 VPWR _0444_ 0.16285f
C46222 _0804_/a_79_21# _0804_/a_297_297# 0.01735f
C46223 _0463_ _0935_/a_27_47# 0
C46224 hold57/a_285_47# net29 0
C46225 acc0.A\[20\] _0236_ 0.00323f
C46226 _0174_ _0543_/a_150_297# 0.00146f
C46227 clknet_0__0463_ _0493_/a_27_47# 0.00563f
C46228 _0536_/a_51_297# _1046_/a_634_159# 0
C46229 _0233_ _0368_ 0
C46230 _0320_ _0365_ 0
C46231 _0520_/a_109_297# clknet_1_0__leaf__0465_ 0.00141f
C46232 control0.add clknet_1_1__leaf_clk 0
C46233 acc0.A\[5\] hold1/a_49_47# 0.32626f
C46234 acc0.A\[5\] _0989_/a_27_47# 0
C46235 _0292_ _0817_/a_585_47# 0
C46236 net240 _1063_/a_891_413# 0
C46237 _0216_ _0699_/a_150_297# 0
C46238 hold82/a_49_47# hold82/a_285_47# 0.22264f
C46239 _0582_/a_109_47# _0347_ 0
C46240 clknet_1_1__leaf__0459_ acc0.A\[10\] 0.07633f
C46241 _0401_ _0992_/a_27_47# 0
C46242 _0347_ _1007_/a_634_159# 0
C46243 net27 _0132_ 0
C46244 clknet_1_0__leaf__0460_ _1006_/a_193_47# 0.00218f
C46245 _0195_ _1031_/a_27_47# 0.0441f
C46246 _0457_ _1033_/a_592_47# 0
C46247 _0963_/a_117_297# _0481_ 0
C46248 _0375_ _0755_/a_109_297# 0
C46249 _0751_/a_111_297# clknet_1_0__leaf__0460_ 0
C46250 clknet_0__0457_ _0579_/a_27_297# 0.06561f
C46251 hold55/a_391_47# _0457_ 0.01464f
C46252 _1072_/a_193_47# clknet_0_clk 0.0467f
C46253 _1050_/a_193_47# _1050_/a_381_47# 0.09799f
C46254 _1050_/a_634_159# _1050_/a_891_413# 0.03684f
C46255 _1050_/a_27_47# _1050_/a_561_413# 0.0027f
C46256 output64/a_27_47# clknet_1_1__leaf__0458_ 0
C46257 _0643_/a_337_297# VPWR 0
C46258 VPWR _0367_ 1.09434f
C46259 _0330_ _0333_ 0.06052f
C46260 _1019_/a_891_413# clknet_1_0__leaf__0457_ 0.00444f
C46261 _0557_/a_240_47# comp0.B\[5\] 0
C46262 net36 _0854_/a_79_21# 0.01584f
C46263 _0398_ _0369_ 0
C46264 net90 net50 0
C46265 hold85/a_49_47# _0946_/a_30_53# 0
C46266 clkload1/Y _0432_ 0
C46267 _0221_ _1011_/a_381_47# 0.01678f
C46268 _0958_/a_27_47# _0958_/a_303_47# 0.00119f
C46269 _0869_/a_27_47# _0352_ 0
C46270 _0179_ _1049_/a_1017_47# 0
C46271 _0427_ _0290_ 0.01193f
C46272 _0337_ net44 0
C46273 _1036_/a_27_47# net28 0
C46274 _0565_/a_51_297# _0565_/a_512_297# 0.0116f
C46275 clknet_1_0__leaf__0462_ hold90/a_391_47# 0
C46276 net46 control0.add 0.26701f
C46277 _0178_ _0173_ 0
C46278 _0680_/a_80_21# VPWR 0.27478f
C46279 net203 net24 0.10177f
C46280 _0718_/a_285_47# VPWR 0.00234f
C46281 _0461_ _0769_/a_81_21# 0.00259f
C46282 _0222_ _0377_ 0.11693f
C46283 clknet_0__0464_ net132 0.36921f
C46284 _0997_/a_975_413# pp[14] 0
C46285 _0998_/a_466_413# net43 0
C46286 _1071_/a_1017_47# clknet_0_clk 0
C46287 _0640_/a_215_297# _0269_ 0
C46288 _0852_/a_35_297# _0399_ 0
C46289 _1054_/a_27_47# _1052_/a_1059_315# 0
C46290 net206 clknet_1_0__leaf__0457_ 0
C46291 hold88/a_49_47# _0186_ 0.04202f
C46292 _0470_ _0132_ 0
C46293 net224 _1009_/a_891_413# 0.00187f
C46294 _0403_ net38 0
C46295 _0176_ _1040_/a_27_47# 0.05166f
C46296 _0982_/a_634_159# net149 0
C46297 net1 _0181_ 0.28572f
C46298 _1039_/a_193_47# _0463_ 0.03247f
C46299 output61/a_27_47# pp[3] 0.33815f
C46300 clkbuf_1_1__f__0457_/a_110_47# _0526_/a_27_47# 0.00236f
C46301 _0538_/a_240_47# _1044_/a_466_413# 0
C46302 acc0.A\[27\] _0331_ 0
C46303 _0217_ VPWR 5.94174f
C46304 _1004_/a_27_47# net53 0
C46305 comp0.B\[11\] net129 0
C46306 _1056_/a_634_159# _0179_ 0.04423f
C46307 _0533_/a_27_297# control0.reset 0.02847f
C46308 hold46/a_285_47# comp0.B\[13\] 0.02036f
C46309 clknet_1_1__leaf__0461_ _0507_/a_27_297# 0
C46310 _0486_ _1068_/a_561_413# 0.00275f
C46311 _0143_ _1045_/a_381_47# 0
C46312 _0353_ _0724_/a_113_297# 0.00758f
C46313 _0555_/a_51_297# _0173_ 0.07918f
C46314 hold46/a_391_47# _1046_/a_27_47# 0
C46315 hold46/a_285_47# _1046_/a_193_47# 0
C46316 hold57/a_49_47# _0494_/a_27_47# 0
C46317 _0258_ acc0.A\[8\] 0
C46318 clkload4/Y _1016_/a_1059_315# 0.00161f
C46319 hold10/a_49_47# _0180_ 0.02082f
C46320 _0343_ _1000_/a_381_47# 0.00149f
C46321 _0574_/a_27_297# _1007_/a_27_47# 0
C46322 _0273_ net74 0
C46323 _0817_/a_81_21# clknet_1_1__leaf__0465_ 0.00378f
C46324 _1033_/a_466_413# _0208_ 0
C46325 _0183_ _1015_/a_193_47# 0.00249f
C46326 _0269_ _0465_ 0.07569f
C46327 _0081_ _0399_ 0.18399f
C46328 _0999_/a_1059_315# net85 0
C46329 _0426_ _0181_ 0
C46330 _1001_/a_891_413# _1019_/a_1059_315# 0
C46331 _1050_/a_27_47# clkbuf_1_0__f__0464_/a_110_47# 0
C46332 _0772_/a_215_47# net223 0.06325f
C46333 _0179_ _0433_ 0
C46334 clkbuf_1_1__f__0458_/a_110_47# _0988_/a_27_47# 0.00103f
C46335 hold76/a_391_47# clkbuf_1_0__f__0461_/a_110_47# 0.01112f
C46336 _0772_/a_297_297# _0391_ 0.00133f
C46337 net231 clknet_1_1__leaf_clk 0.14718f
C46338 _0310_ _0777_/a_47_47# 0
C46339 VPWR _0993_/a_975_413# 0.00464f
C46340 _1016_/a_193_47# net221 0.04977f
C46341 net168 input11/a_75_212# 0.03682f
C46342 _0752_/a_27_413# _0234_ 0.21503f
C46343 acc0.A\[2\] _0269_ 0
C46344 clknet_1_0__leaf__0462_ _1007_/a_975_413# 0
C46345 output56/a_27_47# _0345_ 0.01421f
C46346 _0732_/a_80_21# _0732_/a_209_297# 0.06257f
C46347 _0715_/a_27_47# _0423_ 0
C46348 _0271_ _0186_ 0.00145f
C46349 hold91/a_285_47# _0345_ 0.01934f
C46350 _0971_/a_81_21# clkbuf_1_1__f_clk/a_110_47# 0.00788f
C46351 hold31/a_49_47# acc0.A\[6\] 0.00911f
C46352 clknet_1_1__leaf__0459_ net43 0.0255f
C46353 _0983_/a_1059_315# _0183_ 0
C46354 VPWR _0542_/a_51_297# 0.46977f
C46355 net194 comp0.B\[14\] 0
C46356 net106 control0.reset 0
C46357 net47 _0347_ 0.07707f
C46358 _0312_ _0360_ 0.00138f
C46359 _0305_ _0289_ 0.03403f
C46360 _0186_ _0987_/a_891_413# 0
C46361 _0996_/a_1059_315# _0790_/a_35_297# 0
C46362 _0172_ _0954_/a_32_297# 0.00312f
C46363 _0232_ _0219_ 0.03341f
C46364 hold20/a_49_47# hold20/a_391_47# 0.00188f
C46365 _1043_/a_27_47# _0203_ 0
C46366 input32/a_75_212# _0140_ 0
C46367 B[9] net18 0
C46368 clknet_1_0__leaf__0465_ net147 0.11029f
C46369 _0273_ output61/a_27_47# 0
C46370 net81 _0297_ 0
C46371 hold38/a_49_47# _0564_/a_150_297# 0
C46372 _0818_/a_193_47# _0291_ 0
C46373 _0723_/a_27_413# _0705_/a_59_75# 0
C46374 _0181_ _0185_ 0.15746f
C46375 _0328_ _0745_/a_193_47# 0
C46376 _1001_/a_1059_315# net206 0
C46377 net185 B[2] 0
C46378 hold32/a_285_47# _0153_ 0.01023f
C46379 _0479_ _0975_/a_59_75# 0.00119f
C46380 _0274_ _0435_ 0
C46381 _1016_/a_466_413# _0459_ 0
C46382 hold88/a_285_47# _0253_ 0
C46383 _0648_/a_277_297# _0278_ 0
C46384 _0648_/a_109_297# _0280_ 0
C46385 _0285_ net228 0
C46386 _0217_ net48 0.02056f
C46387 VPWR _0142_ 1.56213f
C46388 _1030_/a_27_47# _0333_ 0
C46389 hold17/a_49_47# _0169_ 0.00106f
C46390 clknet_1_1__leaf__0459_ _0999_/a_27_47# 0.0077f
C46391 hold38/a_285_47# clknet_1_1__leaf_clk 0.01877f
C46392 net129 _0202_ 0.00406f
C46393 clknet_0__0458_ _0840_/a_68_297# 0.00509f
C46394 _0964_/a_109_297# clk 0
C46395 _1006_/a_561_413# _0219_ 0
C46396 _0288_ _0345_ 0.06013f
C46397 _0136_ comp0.B\[8\] 0
C46398 _0412_ net81 0
C46399 _0947_/a_109_297# _0166_ 0
C46400 _0467_ _1068_/a_592_47# 0
C46401 _0614_/a_111_297# _0245_ 0
C46402 hold100/a_285_47# hold100/a_391_47# 0.41909f
C46403 _0712_/a_79_21# _0195_ 0.00108f
C46404 _0985_/a_634_159# _0985_/a_975_413# 0
C46405 _0985_/a_466_413# _0985_/a_561_413# 0.00772f
C46406 hold39/a_49_47# comp0.B\[6\] 0.02567f
C46407 _0183_ hold29/a_391_47# 0
C46408 _0951_/a_109_93# _0175_ 0
C46409 hold19/a_391_47# net103 0.0017f
C46410 _0326_ _1007_/a_27_47# 0
C46411 _1018_/a_634_159# _1018_/a_381_47# 0
C46412 hold85/a_49_47# _0967_/a_109_93# 0.00193f
C46413 _0956_/a_32_297# clknet_1_0__leaf__0461_ 0
C46414 hold63/a_49_47# hold8/a_285_47# 0
C46415 _0086_ _0253_ 0.0167f
C46416 hold19/a_49_47# _1016_/a_27_47# 0
C46417 _0290_ net142 0.00296f
C46418 _0390_ _0217_ 0
C46419 comp0.B\[14\] _1046_/a_634_159# 0
C46420 _0596_/a_59_75# _0228_ 0.11157f
C46421 _0982_/a_27_47# _0982_/a_891_413# 0.03224f
C46422 _0982_/a_193_47# _0982_/a_1059_315# 0.03202f
C46423 _0982_/a_634_159# _0982_/a_466_413# 0.23992f
C46424 _0222_ net109 0.2705f
C46425 VPWR _0742_/a_299_297# 0.2152f
C46426 _0725_/a_303_47# _0335_ 0
C46427 _1049_/a_27_47# _1049_/a_1059_315# 0.04875f
C46428 _1049_/a_193_47# _1049_/a_466_413# 0.07402f
C46429 _0983_/a_1059_315# acc0.A\[15\] 0.00409f
C46430 clknet_1_1__leaf__0460_ _0732_/a_303_47# 0.00224f
C46431 control0.sh _0951_/a_209_311# 0
C46432 _0430_ _0257_ 0
C46433 net64 _0258_ 0.00503f
C46434 net148 _0522_/a_27_297# 0
C46435 _0524_/a_27_297# acc0.A\[6\] 0
C46436 _1019_/a_592_47# _0459_ 0
C46437 net207 _0869_/a_27_47# 0
C46438 _0324_ net93 0
C46439 _0359_ _0105_ 0.19199f
C46440 _0753_/a_465_47# _0233_ 0.01251f
C46441 _0753_/a_381_47# _0231_ 0
C46442 net180 _0540_/a_149_47# 0
C46443 net125 clknet_1_0__leaf__0465_ 0.00464f
C46444 clkbuf_0__0462_/a_110_47# _0366_ 0
C46445 _0461_ clknet_0__0461_ 0.09805f
C46446 clkload3/a_268_47# clknet_1_1__leaf__0461_ 0.0018f
C46447 clkbuf_1_0__f__0457_/a_110_47# _0345_ 0.01529f
C46448 _0172_ net173 0.20217f
C46449 _1054_/a_634_159# A[8] 0
C46450 hold98/a_49_47# net40 0.29291f
C46451 hold79/a_49_47# net226 0
C46452 hold11/a_391_47# _0172_ 0.00623f
C46453 _0218_ _0099_ 0.02992f
C46454 _0257_ acc0.A\[5\] 0
C46455 _1066_/a_27_47# _1066_/a_1059_315# 0.04755f
C46456 _1066_/a_193_47# _1066_/a_466_413# 0.0802f
C46457 _0473_ _1045_/a_1059_315# 0
C46458 net101 _0216_ 0.02743f
C46459 _0254_ _0431_ 0
C46460 _0782_/a_27_47# clkbuf_0__0457_/a_110_47# 0.00949f
C46461 VPWR _0248_ 0.62727f
C46462 hold37/a_285_47# _1050_/a_27_47# 0
C46463 hold37/a_49_47# _1050_/a_193_47# 0
C46464 hold45/a_285_47# net37 0
C46465 net56 _1010_/a_466_413# 0
C46466 net61 _0625_/a_59_75# 0.0044f
C46467 clknet_0__0459_ _0305_ 0.00741f
C46468 net89 _0381_ 0
C46469 net45 _0999_/a_1059_315# 0.01123f
C46470 clknet_1_1__leaf__0460_ clknet_0__0460_ 0.0406f
C46471 VPWR _1052_/a_891_413# 0.18672f
C46472 _1031_/a_466_413# acc0.A\[30\] 0
C46473 _1023_/a_27_47# _1022_/a_891_413# 0.00437f
C46474 _1023_/a_193_47# _1022_/a_1059_315# 0
C46475 _0080_ _0850_/a_68_297# 0
C46476 _0967_/a_403_297# clk 0
C46477 _1068_/a_27_47# _1068_/a_1059_315# 0.04875f
C46478 _1068_/a_193_47# _1068_/a_466_413# 0.07855f
C46479 _0557_/a_51_297# comp0.B\[4\] 0.01244f
C46480 _0134_ _1036_/a_1059_315# 0
C46481 _0677_/a_285_47# acc0.A\[17\] 0.08048f
C46482 VPWR _0971_/a_81_21# 0.20849f
C46483 _0460_ _0352_ 0.07157f
C46484 clkbuf_1_1__f__0464_/a_110_47# _1045_/a_1059_315# 0
C46485 net54 net244 0
C46486 _0255_ _0825_/a_150_297# 0
C46487 _0502_/a_27_47# net247 0.04421f
C46488 _0797_/a_207_413# _0297_ 0.00414f
C46489 _1032_/a_466_413# net23 0
C46490 net44 _0307_ 0.05315f
C46491 _0992_/a_27_47# hold70/a_49_47# 0.00533f
C46492 clkbuf_0__0465_/a_110_47# net47 0.00113f
C46493 net53 net54 0.00682f
C46494 hold53/a_285_47# hold53/a_391_47# 0.41909f
C46495 _0204_ net198 0.00113f
C46496 _0217_ clknet_1_0__leaf__0459_ 0.02706f
C46497 net71 _1048_/a_27_47# 0
C46498 _0519_/a_384_47# net65 0
C46499 _0519_/a_299_297# acc0.A\[7\] 0.03109f
C46500 _0946_/a_30_53# net17 0
C46501 _0358_ _0352_ 0.17372f
C46502 clkbuf_0__0460_/a_110_47# _0219_ 0.03188f
C46503 _0268_ _0263_ 0.83544f
C46504 clkbuf_1_0__f__0458_/a_110_47# _0399_ 0.02061f
C46505 _1034_/a_193_47# comp0.B\[2\] 0.04815f
C46506 _1051_/a_634_159# _0186_ 0.00154f
C46507 _0557_/a_149_47# net26 0.00245f
C46508 hold6/a_285_47# net18 0.00476f
C46509 _0765_/a_79_21# _0346_ 0
C46510 output65/a_27_47# acc0.A\[7\] 0
C46511 output65/a_27_47# _0989_/a_1059_315# 0.00155f
C46512 _0343_ acc0.A\[13\] 0.00325f
C46513 _0457_ _0352_ 0.00493f
C46514 acc0.A\[27\] _1008_/a_27_47# 0.03311f
C46515 pp[6] pp[8] 0
C46516 _0710_/a_109_297# clknet_1_1__leaf__0462_ 0
C46517 _0275_ _0785_/a_81_21# 0.03896f
C46518 net25 net27 0.48535f
C46519 VPWR _0164_ 0.24437f
C46520 _0413_ _0797_/a_27_413# 0
C46521 _0979_/a_109_297# _0466_ 0.01277f
C46522 _0979_/a_109_47# _0488_ 0.00487f
C46523 _0983_/a_27_47# _0181_ 0
C46524 net48 _0248_ 0
C46525 _0225_ _0618_/a_297_297# 0
C46526 _0958_/a_27_47# _0485_ 0
C46527 _0787_/a_209_47# net246 0
C46528 _0999_/a_1059_315# _0587_/a_27_47# 0.00242f
C46529 control0.state\[1\] clknet_1_1__leaf_clk 0.46579f
C46530 _0086_ net74 0.03018f
C46531 _0346_ _1006_/a_634_159# 0.04098f
C46532 hold57/a_285_47# comp0.B\[6\] 0.04107f
C46533 control0.state\[0\] _0166_ 0
C46534 _0450_ _0451_ 0.12881f
C46535 _0289_ _0181_ 0.00136f
C46536 clknet_1_0__leaf__0465_ _0473_ 0.00263f
C46537 VPWR _0424_ 0.13318f
C46538 net171 _0176_ 0.18794f
C46539 _0407_ net42 0.33439f
C46540 pp[30] _1031_/a_891_413# 0.00279f
C46541 _1058_/a_1059_315# net2 0
C46542 acc0.A\[17\] _0114_ 0
C46543 _1032_/a_193_47# clknet_1_0__leaf__0461_ 0.04058f
C46544 hold89/a_285_47# _0974_/a_448_47# 0
C46545 _0257_ _0443_ 0.24625f
C46546 _0973_/a_27_297# _0487_ 0.14337f
C46547 hold41/a_49_47# clknet_1_1__leaf__0465_ 0
C46548 _1071_/a_975_413# _0466_ 0
C46549 _1071_/a_592_47# _0488_ 0
C46550 VPWR clknet_0__0463_ 2.26248f
C46551 net85 _0397_ 0
C46552 _0217_ _0453_ 0
C46553 _0183_ _0266_ 0
C46554 _1008_/a_27_47# _0364_ 0
C46555 _0243_ _0372_ 0
C46556 hold8/a_49_47# _0365_ 0
C46557 _0390_ _0248_ 0
C46558 _0993_/a_561_413# _0286_ 0
C46559 _0853_/a_68_297# _0264_ 0
C46560 hold38/a_391_47# VPWR 0.19682f
C46561 clknet_1_0__leaf__0460_ _0103_ 0.039f
C46562 _1013_/a_27_47# clknet_1_1__leaf__0462_ 0
C46563 _0456_ _0117_ 0.00141f
C46564 _0343_ net85 0
C46565 _1017_/a_466_413# net103 0.03199f
C46566 _0708_/a_150_297# net60 0
C46567 _0751_/a_29_53# hold94/a_391_47# 0.00115f
C46568 _1017_/a_193_47# _1016_/a_27_47# 0
C46569 _1017_/a_27_47# _1016_/a_193_47# 0
C46570 clknet_1_0__leaf__0465_ clkbuf_1_1__f__0464_/a_110_47# 0.02118f
C46571 _0233_ _0234_ 0.27337f
C46572 _0343_ _0375_ 0.07129f
C46573 _0430_ _0429_ 0.0069f
C46574 _1052_/a_1017_47# net9 0.00173f
C46575 _0554_/a_68_297# _1036_/a_1059_315# 0
C46576 acc0.A\[8\] _0988_/a_193_47# 0
C46577 net24 _0176_ 0.05374f
C46578 _0966_/a_109_297# _0480_ 0
C46579 net127 comp0.B\[9\] 0
C46580 net10 _1040_/a_1059_315# 0
C46581 clknet_0__0457_ net36 0.05016f
C46582 _0507_/a_373_47# _0185_ 0
C46583 _1000_/a_975_413# net45 0.00196f
C46584 acc0.A\[5\] net11 0
C46585 control0.state\[1\] _0479_ 0
C46586 _0645_/a_47_47# VPWR 0.35379f
C46587 _0804_/a_215_47# _0092_ 0.0014f
C46588 net224 clkbuf_1_1__f__0460_/a_110_47# 0
C46589 _0470_ _0477_ 0.1405f
C46590 _1067_/a_27_47# _1065_/a_27_47# 0
C46591 _0458_ _0267_ 0
C46592 hold82/a_391_47# _0185_ 0
C46593 net44 _0780_/a_285_297# 0
C46594 _0690_/a_68_297# _0324_ 0
C46595 _0476_ _0561_/a_240_47# 0.00523f
C46596 _0521_/a_299_297# net230 0.08168f
C46597 _0521_/a_384_47# _0192_ 0.00157f
C46598 _0855_/a_299_297# acc0.A\[19\] 0
C46599 _0721_/a_27_47# clknet_1_0__leaf__0461_ 0
C46600 _1033_/a_193_47# _1033_/a_592_47# 0.00135f
C46601 _1033_/a_466_413# _1033_/a_561_413# 0.00772f
C46602 _1033_/a_634_159# _1033_/a_975_413# 0
C46603 hold3/a_49_47# net51 0.00131f
C46604 _0329_ net57 0.00967f
C46605 clknet_1_0__leaf__0465_ _0186_ 0.08587f
C46606 _0259_ net66 0.19495f
C46607 clknet_0__0458_ _0255_ 0.02232f
C46608 net194 hold37/a_49_47# 0.00316f
C46609 _1012_/a_193_47# _1012_/a_592_47# 0.00135f
C46610 _1012_/a_466_413# _1012_/a_561_413# 0.00772f
C46611 _1012_/a_634_159# _1012_/a_975_413# 0
C46612 _1039_/a_466_413# _0176_ 0.02342f
C46613 _0995_/a_891_413# net6 0
C46614 hold23/a_391_47# _0186_ 0
C46615 _0195_ _0327_ 0.07184f
C46616 _0712_/a_465_47# acc0.A\[30\] 0
C46617 net36 hold25/a_391_47# 0
C46618 hold79/a_391_47# _0485_ 0
C46619 _0347_ net93 0.18562f
C46620 _0107_ _1009_/a_381_47# 0.12066f
C46621 _0476_ _0472_ 0.00581f
C46622 _0343_ net245 0.11509f
C46623 _1019_/a_1059_315# net149 0
C46624 _0749_/a_299_297# _0462_ 0
C46625 _1009_/a_27_47# _0219_ 0.01381f
C46626 _1015_/a_27_47# comp0.B\[0\] 0
C46627 _0259_ _0991_/a_27_47# 0
C46628 _1050_/a_193_47# acc0.A\[4\] 0.14336f
C46629 hold67/a_391_47# VPWR 0.18515f
C46630 _0266_ acc0.A\[15\] 0.00133f
C46631 _0343_ _1030_/a_1059_315# 0.00283f
C46632 _1055_/a_634_159# acc0.A\[9\] 0
C46633 hold47/a_285_47# net132 0.00207f
C46634 hold26/a_49_47# _0540_/a_240_47# 0
C46635 hold26/a_285_47# _0540_/a_149_47# 0
C46636 _1041_/a_891_413# _0546_/a_240_47# 0
C46637 _1041_/a_27_47# net152 0
C46638 hold100/a_391_47# _0858_/a_27_47# 0
C46639 clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ 1.75875f
C46640 _0967_/a_109_93# net17 0
C46641 _0958_/a_303_47# _0477_ 0
C46642 _0221_ net57 0.43943f
C46643 _0487_ net17 0.10922f
C46644 clknet_0__0459_ _0181_ 0.00136f
C46645 _0746_/a_81_21# clkbuf_0__0460_/a_110_47# 0
C46646 _0508_/a_81_21# _0508_/a_299_297# 0.08213f
C46647 net61 pp[3] 0.12087f
C46648 _0565_/a_240_47# net201 0.05147f
C46649 clkload3/Y acc0.A\[17\] 0.0129f
C46650 comp0.B\[14\] _1045_/a_27_47# 0
C46651 _0294_ _0347_ 0.07853f
C46652 _0544_/a_240_47# _1043_/a_193_47# 0
C46653 net163 _0704_/a_68_297# 0.00251f
C46654 hold16/a_285_47# acc0.A\[30\] 0.00661f
C46655 _0960_/a_27_47# VPWR 0.19425f
C46656 comp0.B\[13\] hold37/a_285_47# 0
C46657 _1004_/a_27_47# _0575_/a_27_297# 0
C46658 net140 _1052_/a_634_159# 0.00109f
C46659 _0254_ _0269_ 0
C46660 _0716_/a_27_47# clkbuf_1_1__f__0459_/a_110_47# 0.00272f
C46661 _0513_/a_299_297# clknet_1_1__leaf__0465_ 0.02271f
C46662 _0181_ control0.sh 0
C46663 _0457_ net207 0
C46664 _0409_ _0277_ 0.16095f
C46665 hold24/a_285_47# net36 0.08785f
C46666 VPWR _0755_/a_109_297# 0.00431f
C46667 hold6/a_49_47# _1043_/a_27_47# 0
C46668 net68 net149 0.22301f
C46669 _1053_/a_27_47# input12/a_75_212# 0
C46670 _0179_ _1054_/a_975_413# 0.00124f
C46671 _0259_ _0350_ 0.02697f
C46672 _0199_ control0.reset 0.03882f
C46673 net64 _0988_/a_193_47# 0.01834f
C46674 net126 _0547_/a_68_297# 0.06977f
C46675 net45 _1018_/a_891_413# 0.00534f
C46676 net45 _0397_ 0.00338f
C46677 _0108_ hold95/a_285_47# 0
C46678 _1031_/a_891_413# _0339_ 0.0079f
C46679 _1003_/a_27_47# _0762_/a_215_47# 0
C46680 _1020_/a_1059_315# clknet_0__0457_ 0.01009f
C46681 _0997_/a_1059_315# _1013_/a_466_413# 0
C46682 _0271_ net62 0.02448f
C46683 net193 _1046_/a_381_47# 0
C46684 input6/a_75_212# net5 0
C46685 _0343_ net45 0.34372f
C46686 _0131_ _0208_ 0.02977f
C46687 comp0.B\[1\] _0173_ 0
C46688 _0779_/a_215_47# _0395_ 0.05495f
C46689 _0443_ _0640_/a_392_297# 0.0012f
C46690 _1001_/a_634_159# _0350_ 0
C46691 VPWR _0235_ 0.34593f
C46692 _0518_/a_109_297# acc0.A\[4\] 0
C46693 _1046_/a_1059_315# _1046_/a_891_413# 0.31086f
C46694 _1046_/a_193_47# _1046_/a_975_413# 0
C46695 _1046_/a_466_413# _1046_/a_381_47# 0.03733f
C46696 _0991_/a_466_413# _0263_ 0
C46697 net233 hold100/a_391_47# 0
C46698 _0183_ _0713_/a_27_47# 0.01103f
C46699 _0481_ _0485_ 0
C46700 _0227_ _0373_ 0
C46701 pp[26] _0570_/a_109_47# 0
C46702 net61 _0273_ 0.01698f
C46703 _1032_/a_561_413# clknet_1_0__leaf__0457_ 0
C46704 net169 net12 0
C46705 control0.state\[0\] _0168_ 0.0024f
C46706 net34 VPWR 2.253f
C46707 _0375_ _0376_ 0.05337f
C46708 hold68/a_391_47# _0122_ 0.0027f
C46709 _0753_/a_381_47# _0225_ 0
C46710 _0180_ hold7/a_285_47# 0
C46711 _1051_/a_1059_315# _1050_/a_27_47# 0.00493f
C46712 _1051_/a_466_413# _1050_/a_193_47# 0
C46713 _1051_/a_193_47# _1050_/a_466_413# 0
C46714 _1051_/a_27_47# _1050_/a_1059_315# 0.00493f
C46715 _1039_/a_193_47# clkbuf_1_0__f__0463_/a_110_47# 0.00594f
C46716 _0684_/a_59_75# _0684_/a_145_75# 0.00658f
C46717 VPWR _0583_/a_373_47# 0.00158f
C46718 _0179_ _0266_ 0
C46719 clknet_1_0__leaf__0462_ hold53/a_285_47# 0.00134f
C46720 _0985_/a_466_413# net175 0
C46721 _0985_/a_27_47# net9 0
C46722 net44 _0333_ 0
C46723 _1050_/a_27_47# _1045_/a_381_47# 0
C46724 hold58/a_391_47# net26 0
C46725 hold9/a_285_47# _1028_/a_27_47# 0
C46726 clkbuf_0__0462_/a_110_47# acc0.A\[24\] 0
C46727 acc0.A\[21\] _0487_ 0
C46728 _0982_/a_27_47# clkbuf_0__0457_/a_110_47# 0
C46729 _0996_/a_975_413# acc0.A\[15\] 0
C46730 hold91/a_49_47# _0301_ 0
C46731 clknet_1_0__leaf__0463_ _1038_/a_381_47# 0.00741f
C46732 _0785_/a_384_47# _0181_ 0
C46733 net196 _0542_/a_240_47# 0.00133f
C46734 net175 _1049_/a_27_47# 0
C46735 _0531_/a_109_297# _1049_/a_891_413# 0
C46736 _0430_ clknet_1_1__leaf__0458_ 0.30194f
C46737 _0183_ _0612_/a_59_75# 0.00619f
C46738 acc0.A\[12\] _1057_/a_975_413# 0
C46739 _0195_ _0306_ 0
C46740 _0292_ _0816_/a_68_297# 0
C46741 _0775_/a_297_297# _0347_ 0.00412f
C46742 _0467_ _0215_ 0
C46743 net166 _0459_ 0
C46744 _0457_ _1032_/a_891_413# 0.01622f
C46745 _0710_/a_109_297# hold92/a_49_47# 0
C46746 net44 _0999_/a_975_413# 0
C46747 _0246_ _0393_ 0
C46748 net59 _0129_ 0.00212f
C46749 acc0.A\[5\] clknet_1_1__leaf__0458_ 0.07918f
C46750 _0181_ net157 0.35714f
C46751 _1016_/a_1059_315# _0218_ 0
C46752 net117 net116 0
C46753 _0179_ hold35/a_49_47# 0
C46754 VPWR _0999_/a_1059_315# 0.41752f
C46755 _1024_/a_27_47# output52/a_27_47# 0
C46756 hold27/a_285_47# _0536_/a_149_47# 0
C46757 hold27/a_49_47# _0536_/a_240_47# 0
C46758 _1052_/a_466_413# acc0.A\[6\] 0.02484f
C46759 _1052_/a_27_47# net13 0
C46760 _0614_/a_29_53# _0352_ 0.013f
C46761 net89 _0468_ 0
C46762 _0226_ acc0.A\[21\] 0.13213f
C46763 _0316_ _0690_/a_68_297# 0.0263f
C46764 hold22/a_391_47# input15/a_75_212# 0.00301f
C46765 _0179_ _0522_/a_109_47# 0
C46766 net48 _0235_ 0.00901f
C46767 _0217_ pp[22] 0
C46768 _0183_ net50 0
C46769 _0984_/a_27_47# net58 0
C46770 comp0.B\[0\] _0215_ 0.7938f
C46771 _0240_ _0308_ 0.00623f
C46772 _0501_/a_27_47# _1061_/a_1059_315# 0
C46773 _0902_/a_27_47# control0.add 0.0265f
C46774 _1018_/a_381_47# net104 0
C46775 _0734_/a_47_47# _0350_ 0.0027f
C46776 net54 clkbuf_1_1__f__0462_/a_110_47# 0
C46777 clkbuf_0__0463_/a_110_47# _0472_ 0.03876f
C46778 _0369_ _0308_ 0
C46779 _0985_/a_193_47# acc0.A\[3\] 0.01649f
C46780 _0690_/a_68_297# _0347_ 0
C46781 comp0.B\[14\] net132 0.01725f
C46782 _0640_/a_215_297# clkbuf_0__0458_/a_110_47# 0
C46783 _0948_/a_109_297# _0468_ 0.01298f
C46784 _0346_ _1014_/a_27_47# 0.0035f
C46785 _0970_/a_27_297# _0162_ 0.16445f
C46786 _0298_ _0409_ 0.21591f
C46787 net194 acc0.A\[4\] 0
C46788 _1053_/a_1059_315# net15 0.00526f
C46789 _1053_/a_634_159# _0191_ 0
C46790 hold101/a_285_47# _0346_ 0.078f
C46791 _0982_/a_634_159# _0080_ 0.00364f
C46792 _0982_/a_466_413# net68 0
C46793 control0.reset _0560_/a_150_297# 0
C46794 net76 _0186_ 0
C46795 _0174_ B[7] 0
C46796 _1049_/a_891_413# _1049_/a_1017_47# 0.00617f
C46797 _1049_/a_193_47# _0147_ 0.28534f
C46798 _1049_/a_634_159# net135 0
C46799 _0653_/a_113_47# acc0.A\[11\] 0
C46800 _0642_/a_215_297# clkbuf_1_1__f__0458_/a_110_47# 0
C46801 net148 _0193_ 0.10034f
C46802 _0194_ acc0.A\[6\] 0
C46803 net40 clknet_1_1__leaf__0459_ 0
C46804 _0598_/a_79_21# hold3/a_49_47# 0.0013f
C46805 _0747_/a_79_21# net216 0.12851f
C46806 _0985_/a_634_159# _0504_/a_27_47# 0
C46807 _0606_/a_215_297# _0606_/a_297_297# 0.00659f
C46808 _0949_/a_59_75# _1062_/a_193_47# 0
C46809 VPWR _0530_/a_81_21# 0.2038f
C46810 _1070_/a_27_47# _1070_/a_1059_315# 0.04875f
C46811 _1070_/a_193_47# _1070_/a_466_413# 0.08301f
C46812 _1052_/a_1059_315# _0523_/a_299_297# 0
C46813 _1052_/a_891_413# _0523_/a_81_21# 0
C46814 _1053_/a_634_159# _1053_/a_381_47# 0
C46815 _0237_ _0460_ 0.00286f
C46816 _0647_/a_47_47# _0647_/a_377_297# 0.00899f
C46817 _1057_/a_634_159# acc0.A\[10\] 0.00115f
C46818 clknet_1_0__leaf__0465_ _1050_/a_634_159# 0.00232f
C46819 hold54/a_391_47# clknet_1_0__leaf__0461_ 0.0047f
C46820 _0329_ _1010_/a_1059_315# 0
C46821 _0465_ clkbuf_0__0458_/a_110_47# 0.0291f
C46822 net45 _0998_/a_193_47# 0.00826f
C46823 net186 _1065_/a_27_47# 0
C46824 net163 _0216_ 0.06673f
C46825 _1066_/a_634_159# clknet_1_1__leaf_clk 0
C46826 _1066_/a_891_413# _1066_/a_1017_47# 0.00617f
C46827 _0314_ _1007_/a_634_159# 0.00167f
C46828 _0313_ _1007_/a_193_47# 0
C46829 _0457_ net106 0.05886f
C46830 _0327_ _1010_/a_891_413# 0
C46831 net222 _0263_ 0
C46832 hold64/a_49_47# net36 0
C46833 _1034_/a_1059_315# _0175_ 0
C46834 _0309_ _0777_/a_47_47# 0.07292f
C46835 hold32/a_49_47# clknet_1_1__leaf__0465_ 0
C46836 net109 _1022_/a_466_413# 0.021f
C46837 _0305_ _0462_ 0.05537f
C46838 _1068_/a_891_413# _1068_/a_1017_47# 0.00617f
C46839 _1068_/a_193_47# _0166_ 0.26947f
C46840 _0290_ _0420_ 0
C46841 _1030_/a_466_413# _1030_/a_561_413# 0.00772f
C46842 _1030_/a_634_159# _1030_/a_975_413# 0
C46843 clkbuf_1_1__f__0464_/a_110_47# _1044_/a_466_413# 0.0068f
C46844 _0696_/a_109_297# acc0.A\[25\] 0
C46845 clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ 1.6264f
C46846 _1038_/a_27_47# _0552_/a_68_297# 0
C46847 clkbuf_1_1__f__0464_/a_110_47# net137 0
C46848 _0627_/a_109_93# _0255_ 0.1059f
C46849 clknet_1_1__leaf__0463_ _0957_/a_32_297# 0
C46850 _0995_/a_193_47# net42 0
C46851 _0270_ _0256_ 0.07401f
C46852 _0443_ clknet_1_1__leaf__0458_ 0.02387f
C46853 hold27/a_49_47# _1046_/a_27_47# 0
C46854 VPWR _0570_/a_373_47# 0
C46855 net202 net23 0.02485f
C46856 _1035_/a_1017_47# clknet_1_1__leaf__0463_ 0
C46857 _0601_/a_150_297# _0366_ 0
C46858 _0992_/a_381_47# net37 0
C46859 _0478_ _0166_ 0
C46860 _0786_/a_300_47# _0401_ 0.00349f
C46861 hold18/a_391_47# _0346_ 0
C46862 clknet_1_1__leaf__0463_ net23 0.0118f
C46863 _0598_/a_297_47# _0226_ 0.05267f
C46864 clkbuf_1_0__f__0459_/a_110_47# acc0.A\[13\] 0.00264f
C46865 _1015_/a_975_413# _0181_ 0.00106f
C46866 _0987_/a_27_47# _0987_/a_561_413# 0.0027f
C46867 _0987_/a_634_159# _0987_/a_891_413# 0.03684f
C46868 _0987_/a_193_47# _0987_/a_381_47# 0.09799f
C46869 _0180_ _0261_ 0.00222f
C46870 _0182_ _0263_ 0
C46871 _0667_/a_113_47# _0299_ 0.00981f
C46872 _0579_/a_109_297# _0183_ 0.07569f
C46873 net194 _1051_/a_466_413# 0
C46874 _0579_/a_373_47# _0217_ 0
C46875 _0261_ net218 0
C46876 _1021_/a_466_413# net106 0
C46877 net137 _0186_ 0.01634f
C46878 acc0.A\[1\] _1047_/a_193_47# 0
C46879 _0182_ _1047_/a_27_47# 0.0273f
C46880 _0713_/a_27_47# hold40/a_285_47# 0
C46881 _0313_ _0328_ 0.15686f
C46882 clknet_1_1__leaf__0457_ _0913_/a_27_47# 0.19403f
C46883 acc0.A\[20\] _0765_/a_297_297# 0.002f
C46884 _0992_/a_975_413# net67 0
C46885 _1000_/a_975_413# VPWR 0.00434f
C46886 _1004_/a_193_47# _1004_/a_466_413# 0.07482f
C46887 _1004_/a_27_47# _1004_/a_1059_315# 0.04819f
C46888 net126 net127 0
C46889 net162 _0128_ 0
C46890 _0557_/a_51_297# _1035_/a_193_47# 0
C46891 net238 net41 0.32678f
C46892 _1072_/a_1017_47# _0466_ 0
C46893 _0151_ _1053_/a_891_413# 0
C46894 _0183_ _0399_ 0.23965f
C46895 net43 _0095_ 0.39326f
C46896 clkload4/a_110_47# acc0.A\[16\] 0
C46897 control0.state\[2\] clknet_0_clk 0.02297f
C46898 _0476_ _0958_/a_197_47# 0.00123f
C46899 _0718_/a_285_47# net56 0
C46900 _0477_ _0485_ 0
C46901 _0195_ _0346_ 0.02262f
C46902 net120 clknet_0_clk 0
C46903 _0534_/a_299_297# _0145_ 0
C46904 input12/a_75_212# A[5] 0.22984f
C46905 _0346_ net92 0.07291f
C46906 _1029_/a_193_47# _1029_/a_381_47# 0.10164f
C46907 _1029_/a_634_159# _1029_/a_891_413# 0.03684f
C46908 _1029_/a_27_47# _1029_/a_561_413# 0.0027f
C46909 _0669_/a_29_53# net6 0
C46910 _0462_ hold73/a_49_47# 0.02669f
C46911 hold37/a_49_47# _1045_/a_27_47# 0
C46912 net211 _0580_/a_109_297# 0
C46913 hold67/a_391_47# hold35/a_391_47# 0
C46914 VPWR _0565_/a_512_297# 0.00729f
C46915 acc0.A\[1\] _0459_ 0
C46916 comp0.B\[15\] _0499_/a_59_75# 0.00579f
C46917 _0448_ _0345_ 0.06699f
C46918 net9 _0197_ 0
C46919 _0165_ _0487_ 0.02885f
C46920 clkbuf_1_1__f__0465_/a_110_47# acc0.A\[10\] 0
C46921 net39 _0345_ 0
C46922 _0268_ _0848_/a_27_47# 0
C46923 _0343_ _0998_/a_1017_47# 0
C46924 _0119_ _0352_ 0
C46925 net94 _0321_ 0
C46926 _0425_ net47 0
C46927 clkload0/a_27_47# _1072_/a_1059_315# 0.01217f
C46928 _0621_/a_35_297# _0253_ 0.17177f
C46929 comp0.B\[13\] _1045_/a_381_47# 0
C46930 acc0.A\[4\] _0987_/a_193_47# 0.0355f
C46931 _0218_ _0268_ 0
C46932 net99 _0219_ 0.03066f
C46933 acc0.A\[12\] _0304_ 0.18349f
C46934 clknet_1_0__leaf__0465_ _0200_ 0.00133f
C46935 acc0.A\[29\] _0701_/a_80_21# 0.00219f
C46936 _1041_/a_1059_315# clkbuf_1_0__f__0463_/a_110_47# 0
C46937 _0661_/a_109_297# _0289_ 0.00576f
C46938 _0661_/a_27_297# _0287_ 0.19391f
C46939 _0581_/a_109_297# _0347_ 0
C46940 clkbuf_0__0462_/a_110_47# _0691_/a_68_297# 0.00989f
C46941 A[10] _0514_/a_109_47# 0
C46942 clknet_1_0__leaf__0465_ net62 0
C46943 control0.count\[3\] _1068_/a_27_47# 0
C46944 _1037_/a_561_413# clknet_1_1__leaf__0463_ 0
C46945 _0378_ _1023_/a_634_159# 0
C46946 clknet_1_0__leaf__0465_ comp0.B\[8\] 0
C46947 _1033_/a_891_413# _0956_/a_32_297# 0
C46948 _0960_/a_181_47# _0976_/a_505_21# 0
C46949 _0555_/a_51_297# net204 0.07935f
C46950 _1028_/a_634_159# _1028_/a_1059_315# 0
C46951 _1028_/a_27_47# _1028_/a_381_47# 0.05761f
C46952 _1028_/a_193_47# _1028_/a_891_413# 0.19226f
C46953 hold41/a_391_47# hold42/a_285_47# 0
C46954 hold41/a_285_47# hold42/a_391_47# 0
C46955 net201 _0171_ 0.08198f
C46956 _0182_ clknet_1_0__leaf__0461_ 0.00124f
C46957 _0371_ _0324_ 0
C46958 clknet_0__0459_ clknet_1_1__leaf__0461_ 0.02112f
C46959 _0369_ _0989_/a_634_159# 0
C46960 _0399_ acc0.A\[15\] 0.09915f
C46961 _0452_ net165 0
C46962 _0441_ _0835_/a_78_199# 0.10637f
C46963 _0837_/a_266_297# _0255_ 0
C46964 _0440_ _0835_/a_292_297# 0
C46965 _0216_ hold60/a_285_47# 0
C46966 net58 _0986_/a_561_413# 0
C46967 _1033_/a_1059_315# comp0.B\[1\] 0.08468f
C46968 _1033_/a_561_413# _0131_ 0
C46969 _0369_ _0992_/a_634_159# 0
C46970 _0852_/a_35_297# _0346_ 0.03234f
C46971 _0985_/a_381_47# VPWR 0.07715f
C46972 net63 _0987_/a_975_413# 0
C46973 _0553_/a_51_297# _0176_ 0.00277f
C46974 _0554_/a_150_297# net26 0
C46975 _0444_ _0345_ 0.05312f
C46976 VPWR _0397_ 0.2035f
C46977 VPWR _1018_/a_891_413# 0.17994f
C46978 acc0.A\[11\] _0651_/a_113_47# 0
C46979 _0722_/a_79_21# net239 0.00117f
C46980 clknet_1_1__leaf__0460_ _0355_ 0
C46981 _0343_ _0439_ 0
C46982 VPWR _1049_/a_466_413# 0.25026f
C46983 _0244_ net221 0
C46984 _0802_/a_59_75# _0647_/a_47_47# 0
C46985 _0647_/a_285_47# clknet_1_1__leaf__0459_ 0.04376f
C46986 hold55/a_391_47# _0130_ 0
C46987 _0179_ _0516_/a_27_297# 0
C46988 _0343_ VPWR 8.4788f
C46989 _0743_/a_240_47# _0315_ 0
C46990 _0743_/a_149_47# _0367_ 0.018f
C46991 acc0.A\[1\] _0265_ 0.12334f
C46992 _0100_ hold93/a_285_47# 0.00147f
C46993 _1041_/a_193_47# net31 0.13201f
C46994 net88 hold93/a_391_47# 0.02624f
C46995 _0662_/a_81_21# net67 0
C46996 net61 acc0.A\[4\] 0
C46997 hold97/a_285_47# _1008_/a_27_47# 0.00403f
C46998 VPWR _1066_/a_466_413# 0.28054f
C46999 _0285_ _0401_ 0
C47000 _0172_ clknet_1_1__leaf__0457_ 0.08158f
C47001 VPWR net95 0.40376f
C47002 _0118_ _0216_ 0
C47003 VPWR _1068_/a_466_413# 0.24331f
C47004 net141 acc0.A\[9\] 0
C47005 _0428_ _0369_ 0.14699f
C47006 _0454_ _0853_/a_68_297# 0.05587f
C47007 _0081_ _0346_ 0
C47008 hold13/a_49_47# _0463_ 0.00243f
C47009 _0367_ _0345_ 0.18128f
C47010 _0258_ hold101/a_391_47# 0
C47011 _0300_ _0406_ 0
C47012 _1051_/a_1059_315# _0987_/a_27_47# 0
C47013 _0388_ _0459_ 0
C47014 _0462_ _0181_ 0.02729f
C47015 _0993_/a_193_47# _0419_ 0
C47016 _0993_/a_466_413# _0417_ 0
C47017 VPWR net198 0.33058f
C47018 clknet_0__0457_ hold60/a_391_47# 0
C47019 _0518_/a_27_297# acc0.A\[8\] 0.06074f
C47020 clknet_0__0458_ _0843_/a_68_297# 0
C47021 _0828_/a_113_297# _0435_ 0.05193f
C47022 A[7] input15/a_75_212# 0
C47023 net1 _1015_/a_27_47# 0.03878f
C47024 clknet_1_0__leaf__0460_ _1067_/a_975_413# 0
C47025 net18 _1043_/a_381_47# 0
C47026 net198 _1043_/a_561_413# 0
C47027 _0478_ _0168_ 0
C47028 clknet_1_0__leaf__0465_ _1046_/a_466_413# 0.0022f
C47029 clknet_1_1__leaf__0460_ _0693_/a_150_297# 0
C47030 _0642_/a_298_297# acc0.A\[8\] 0
C47031 _0343_ _0983_/a_381_47# 0
C47032 _0531_/a_109_47# net175 0
C47033 _0170_ _1071_/a_634_159# 0
C47034 _1016_/a_27_47# net219 0
C47035 _0996_/a_193_47# acc0.A\[13\] 0
C47036 _0699_/a_150_297# _0319_ 0
C47037 _0718_/a_285_47# _0345_ 0
C47038 acc0.A\[21\] _0760_/a_47_47# 0.01253f
C47039 _0343_ output62/a_27_47# 0
C47040 net45 _0793_/a_51_297# 0.00301f
C47041 _1019_/a_634_159# clkbuf_0__0457_/a_110_47# 0.0075f
C47042 _0998_/a_634_159# _0998_/a_592_47# 0
C47043 _0093_ net42 0
C47044 _0579_/a_27_297# hold40/a_391_47# 0.00604f
C47045 _0579_/a_109_297# hold40/a_285_47# 0
C47046 _1009_/a_193_47# _0318_ 0
C47047 clknet_1_1__leaf__0459_ _0806_/a_113_297# 0.00315f
C47048 _0621_/a_35_297# net74 0.04005f
C47049 _0179_ _0399_ 0.12057f
C47050 _0529_/a_373_47# _0186_ 0.00128f
C47051 _0498_/a_512_297# _0465_ 0
C47052 hold10/a_391_47# net247 0
C47053 _0410_ _0400_ 0.67728f
C47054 _0217_ _0345_ 0.06635f
C47055 _0122_ _1023_/a_891_413# 0
C47056 _1024_/a_634_159# acc0.A\[23\] 0
C47057 _0404_ _0788_/a_68_297# 0.11246f
C47058 _0343_ net48 0
C47059 clkbuf_1_1__f__0463_/a_110_47# comp0.B\[6\] 0.0269f
C47060 clknet_0__0463_ comp0.B\[3\] 0
C47061 hold38/a_391_47# comp0.B\[3\] 0.0674f
C47062 hold38/a_49_47# comp0.B\[5\] 0
C47063 _1059_/a_27_47# _0294_ 0
C47064 _0496_/a_27_47# _0173_ 0.00741f
C47065 _0174_ _1044_/a_891_413# 0
C47066 _1019_/a_1059_315# _1019_/a_891_413# 0.31086f
C47067 _1019_/a_193_47# _1019_/a_975_413# 0
C47068 _1019_/a_466_413# _1019_/a_381_47# 0.03733f
C47069 _0089_ _0263_ 0
C47070 _1058_/a_27_47# net37 0.03242f
C47071 comp0.B\[2\] _0171_ 0
C47072 clknet_1_0__leaf__0464_ net8 0
C47073 net133 _0182_ 0.00771f
C47074 net72 _0986_/a_466_413# 0
C47075 VPWR _1012_/a_381_47# 0.07964f
C47076 _0482_ _0484_ 0.09855f
C47077 hold54/a_49_47# _0208_ 0.00603f
C47078 _0469_ _1063_/a_193_47# 0
C47079 clkbuf_0_clk/a_110_47# _0468_ 0.15275f
C47080 _0083_ net175 0
C47081 _1050_/a_466_413# net184 0
C47082 acc0.A\[4\] _1045_/a_27_47# 0
C47083 _1050_/a_1059_315# net131 0
C47084 _0726_/a_51_297# _0726_/a_512_297# 0.0116f
C47085 _0217_ hold2/a_49_47# 0
C47086 net117 _0220_ 0.04962f
C47087 _1058_/a_634_159# net67 0.01912f
C47088 net9 _1049_/a_975_413# 0.00103f
C47089 input2/a_75_212# net66 0.00223f
C47090 net44 _0998_/a_891_413# 0
C47091 hold58/a_49_47# _1035_/a_27_47# 0.00146f
C47092 _0982_/a_27_47# _0350_ 0
C47093 acc0.A\[1\] _0585_/a_109_297# 0.00117f
C47094 _0533_/a_109_297# net149 0
C47095 _0182_ _0585_/a_27_297# 0
C47096 net162 _1031_/a_1059_315# 0
C47097 VPWR _0998_/a_193_47# 0.2965f
C47098 hold3/a_49_47# hold3/a_391_47# 0.00188f
C47099 _0338_ hold61/a_49_47# 0.04808f
C47100 _0335_ hold61/a_285_47# 0
C47101 clknet_1_0__leaf__0465_ _0987_/a_634_159# 0.005f
C47102 _0373_ _0352_ 0.00128f
C47103 _0991_/a_27_47# _0446_ 0
C47104 _1021_/a_891_413# _0578_/a_109_297# 0
C47105 _0758_/a_297_297# _0352_ 0.0059f
C47106 _0758_/a_79_21# _0102_ 0.05113f
C47107 net36 _0210_ 0
C47108 _0221_ _0700_/a_113_47# 0
C47109 _0589_/a_113_47# _0332_ 0
C47110 _0950_/a_75_212# _1063_/a_381_47# 0
C47111 _1024_/a_975_413# net52 0
C47112 _0786_/a_80_21# net67 0
C47113 clkload3/Y net84 0.00961f
C47114 _0216_ _0320_ 0
C47115 _0294_ _0991_/a_1059_315# 0.01715f
C47116 _0991_/a_466_413# _0218_ 0
C47117 _0376_ VPWR 0.42902f
C47118 _0990_/a_466_413# _0990_/a_561_413# 0.00772f
C47119 _0990_/a_634_159# _0990_/a_975_413# 0
C47120 net63 clkbuf_1_1__f__0458_/a_110_47# 0
C47121 _0404_ _0406_ 0
C47122 clknet_0__0461_ _0115_ 0
C47123 _0461_ _0771_/a_215_297# 0.00288f
C47124 _0769_/a_299_297# _0614_/a_29_53# 0
C47125 clknet_1_0__leaf__0465_ input12/a_75_212# 0.01818f
C47126 net76 net62 0.20644f
C47127 _1002_/a_1059_315# clknet_1_0__leaf__0457_ 0.00241f
C47128 _1002_/a_634_159# _0460_ 0.00968f
C47129 _0361_ clkbuf_0__0462_/a_110_47# 0.02295f
C47130 _0329_ clkbuf_1_1__f__0460_/a_110_47# 0
C47131 _0571_/a_109_297# hold8/a_391_47# 0
C47132 _0304_ net42 0.07266f
C47133 _0288_ _0809_/a_299_297# 0
C47134 _0172_ net19 0.08852f
C47135 _0357_ _0722_/a_79_21# 0
C47136 clknet_1_0__leaf__0458_ _0635_/a_27_47# 0.00523f
C47137 hold86/a_391_47# _0268_ 0
C47138 hold49/a_285_47# _0176_ 0
C47139 _0254_ clkbuf_0__0458_/a_110_47# 0
C47140 _0393_ _0774_/a_68_297# 0.10705f
C47141 pp[18] net60 0.00452f
C47142 output44/a_27_47# pp[17] 0.16974f
C47143 hold24/a_285_47# _1039_/a_27_47# 0
C47144 _0805_/a_27_47# _0992_/a_1059_315# 0
C47145 net68 _0080_ 0.00809f
C47146 hold53/a_285_47# _1025_/a_891_413# 0
C47147 _0123_ _1025_/a_193_47# 0
C47148 hold66/a_49_47# clknet_1_0__leaf__0460_ 0
C47149 net155 net113 0
C47150 _1034_/a_891_413# _0955_/a_32_297# 0
C47151 _1051_/a_27_47# _1051_/a_193_47# 0.9705f
C47152 _0446_ _0350_ 0.97977f
C47153 clknet_1_1__leaf_clk _0564_/a_68_297# 0
C47154 clknet_1_0__leaf__0459_ _1018_/a_891_413# 0
C47155 VPWR net38 1.42176f
C47156 _0371_ _0104_ 0
C47157 _0280_ _0405_ 0
C47158 _0218_ clkbuf_1_0__f__0461_/a_110_47# 0.18382f
C47159 VPWR A[14] 0.26501f
C47160 _0258_ _0369_ 0
C47161 _0606_/a_109_53# _0238_ 0
C47162 _0606_/a_392_297# _0236_ 0.00267f
C47163 _0850_/a_150_297# _0264_ 0.00154f
C47164 _1070_/a_891_413# _1070_/a_1017_47# 0.00617f
C47165 _1070_/a_466_413# VPWR 0.29326f
C47166 _1070_/a_193_47# _0168_ 0.21118f
C47167 net106 _1033_/a_193_47# 0
C47168 _1045_/a_634_159# _1045_/a_466_413# 0.23992f
C47169 _1045_/a_193_47# _1045_/a_1059_315# 0.03405f
C47170 _1045_/a_27_47# _1045_/a_891_413# 0.03224f
C47171 _1052_/a_975_413# _0150_ 0
C47172 _0348_ _0219_ 0
C47173 _1053_/a_381_47# net139 0
C47174 _0170_ _0978_/a_27_297# 0
C47175 _0231_ _0693_/a_68_297# 0
C47176 _0343_ clknet_1_0__leaf__0459_ 0.22247f
C47177 net44 _1030_/a_1017_47# 0.00125f
C47178 clknet_1_0__leaf__0465_ net136 0.0011f
C47179 clkbuf_1_0__f__0458_/a_110_47# _0346_ 0
C47180 clknet_1_0__leaf__0462_ hold30/a_285_47# 0.02497f
C47181 _0426_ clknet_1_1__leaf__0465_ 0.03112f
C47182 _1066_/a_592_47# control0.sh 0
C47183 comp0.B\[12\] _0541_/a_68_297# 0
C47184 _1014_/a_381_47# _0465_ 0
C47185 _0552_/a_68_297# B[6] 0
C47186 VPWR _1030_/a_381_47# 0.07542f
C47187 clknet_1_0__leaf__0464_ net10 0.35545f
C47188 clknet_1_1__leaf__0463_ _0213_ 0.0568f
C47189 _0314_ net93 0
C47190 _0378_ _0377_ 0.06597f
C47191 _0783_/a_79_21# _0397_ 0.06429f
C47192 _0135_ _0176_ 0.01234f
C47193 _1043_/a_634_159# _1043_/a_466_413# 0.23992f
C47194 _1043_/a_193_47# _1043_/a_1059_315# 0.03405f
C47195 _1043_/a_27_47# _1043_/a_891_413# 0.03224f
C47196 _0531_/a_27_297# net157 0
C47197 _0376_ net48 0.00174f
C47198 A[3] B[10] 0.17476f
C47199 net109 net151 0.10546f
C47200 _0248_ _0345_ 0.04752f
C47201 pp[27] net116 0
C47202 _1038_/a_1059_315# _0209_ 0.08707f
C47203 _0367_ net52 0.00338f
C47204 hold63/a_391_47# net200 0
C47205 net216 _0745_/a_193_47# 0
C47206 _0747_/a_79_21# _0370_ 0.02886f
C47207 pp[28] net242 0
C47208 hold52/a_285_47# _0217_ 0.01334f
C47209 _0763_/a_193_47# _0460_ 0
C47210 _1021_/a_634_159# _1002_/a_466_413# 0
C47211 _1021_/a_466_413# _1002_/a_634_159# 0.00564f
C47212 _1004_/a_466_413# VPWR 0.25976f
C47213 _1021_/a_891_413# _1002_/a_27_47# 0
C47214 _1021_/a_1059_315# _1002_/a_193_47# 0
C47215 _1021_/a_27_47# _1002_/a_891_413# 0
C47216 hold89/a_285_47# _0484_ 0
C47217 _0153_ input16/a_75_212# 0.02696f
C47218 _0216_ _0720_/a_68_297# 0.00118f
C47219 clknet_1_1__leaf__0465_ _0185_ 0.03435f
C47220 comp0.B\[7\] _1040_/a_1059_315# 0
C47221 clknet_1_0__leaf__0462_ _0102_ 0.00628f
C47222 clknet_1_0__leaf__0458_ _1047_/a_891_413# 0
C47223 _0174_ _1042_/a_27_47# 0.00176f
C47224 _0645_/a_285_47# _0277_ 0.04387f
C47225 hold65/a_285_47# acc0.A\[6\] 0.03101f
C47226 _0180_ _0173_ 0
C47227 _1056_/a_466_413# _1056_/a_561_413# 0.00772f
C47228 _1032_/a_592_47# net17 0
C47229 hold28/a_285_47# _0180_ 0.00232f
C47230 _0407_ net5 0
C47231 comp0.B\[10\] _1042_/a_634_159# 0
C47232 acc0.A\[5\] _0218_ 0.1049f
C47233 _0294_ _0425_ 0.02738f
C47234 _0401_ _0218_ 0
C47235 _0179_ _0295_ 0
C47236 output55/a_27_47# _0357_ 0.00108f
C47237 hold28/a_285_47# net218 0
C47238 net194 _1044_/a_1059_315# 0
C47239 _0680_/a_80_21# net52 0
C47240 _0332_ _0219_ 0.01271f
C47241 _0987_/a_1059_315# _0085_ 0.06492f
C47242 _0987_/a_891_413# net73 0
C47243 _0704_/a_150_297# hold92/a_49_47# 0
C47244 _0651_/a_113_47# _0281_ 0
C47245 net194 _0149_ 0
C47246 _0130_ _0352_ 0
C47247 clkload2/Y clknet_1_0__leaf__0464_ 0.33832f
C47248 _0664_/a_79_21# net37 0
C47249 clknet_1_0__leaf__0458_ _0850_/a_68_297# 0
C47250 _0212_ clknet_1_1__leaf__0463_ 0.04302f
C47251 _0849_/a_79_21# _0451_ 0.071f
C47252 pp[15] pp[31] 0
C47253 _0199_ _1047_/a_561_413# 0
C47254 acc0.A\[31\] _0219_ 0
C47255 _0219_ _0685_/a_68_297# 0
C47256 _0217_ net52 0.03579f
C47257 _0728_/a_59_75# _0332_ 0.01845f
C47258 VPWR hold81/a_285_47# 0.29109f
C47259 _1004_/a_891_413# _1004_/a_1017_47# 0.00617f
C47260 net171 net28 0
C47261 _0949_/a_59_75# net17 0
C47262 _0218_ net222 0.00181f
C47263 _1027_/a_1059_315# _1008_/a_381_47# 0
C47264 clknet_0__0462_ acc0.A\[25\] 0.0031f
C47265 output57/a_27_47# hold80/a_285_47# 0
C47266 hold47/a_49_47# _0196_ 0
C47267 net162 _0712_/a_561_47# 0
C47268 _1059_/a_193_47# _0158_ 0
C47269 _0157_ _1060_/a_193_47# 0
C47270 _1067_/a_891_413# hold93/a_391_47# 0
C47271 _0983_/a_193_47# _0983_/a_634_159# 0.12497f
C47272 _0983_/a_27_47# _0983_/a_466_413# 0.26005f
C47273 _0148_ _0186_ 0.22853f
C47274 _0222_ _0460_ 0
C47275 _0305_ _0312_ 0.04614f
C47276 hold34/a_49_47# net16 0.00117f
C47277 net45 clkbuf_0__0461_/a_110_47# 0.0038f
C47278 _0224_ VPWR 0.43744f
C47279 clknet_1_0__leaf__0465_ _1045_/a_193_47# 0.00546f
C47280 _0343_ hold35/a_391_47# 0
C47281 hold69/a_391_47# clknet_0__0460_ 0
C47282 _1029_/a_1059_315# net191 0
C47283 hold98/a_49_47# _0995_/a_27_47# 0.01168f
C47284 net138 _0150_ 0
C47285 _0245_ _0350_ 0
C47286 net24 net28 0.51006f
C47287 _0334_ hold80/a_391_47# 0.00451f
C47288 acc0.A\[22\] clknet_1_0__leaf__0460_ 0.00177f
C47289 _0244_ _0772_/a_215_47# 0
C47290 _0769_/a_81_21# net223 0
C47291 _0330_ acc0.A\[29\] 0.00291f
C47292 comp0.B\[13\] _1044_/a_891_413# 0
C47293 _0328_ _0321_ 0.0495f
C47294 _0424_ _0345_ 0.01544f
C47295 clknet_0__0459_ clkbuf_1_1__f__0459_/a_110_47# 0.31414f
C47296 _0424_ _0814_/a_27_47# 0.08818f
C47297 clknet_1_0__leaf__0462_ _0574_/a_109_47# 0
C47298 _0830_/a_79_21# pp[5] 0
C47299 _0328_ clkbuf_0__0460_/a_110_47# 0.00206f
C47300 clkbuf_1_1__f__0463_/a_110_47# net26 0.00203f
C47301 net213 net241 0
C47302 clknet_1_0__leaf__0459_ _0998_/a_193_47# 0.00377f
C47303 _1020_/a_891_413# _0183_ 0
C47304 _0278_ net80 0
C47305 _1003_/a_27_47# net150 0
C47306 _0806_/a_199_47# _0281_ 0.01114f
C47307 _0287_ _0293_ 0.00162f
C47308 net162 hold16/a_391_47# 0.002f
C47309 _1013_/a_27_47# _0218_ 0.02453f
C47310 _0854_/a_215_47# clknet_1_0__leaf__0461_ 0
C47311 _1016_/a_634_159# _1016_/a_381_47# 0
C47312 hold13/a_391_47# _0176_ 0
C47313 _0548_/a_51_297# net147 0
C47314 _0138_ _1061_/a_27_47# 0
C47315 _0699_/a_68_297# _0330_ 0.0272f
C47316 VPWR _0726_/a_512_297# 0.00729f
C47317 hold11/a_49_47# _0465_ 0
C47318 _0179_ _0619_/a_68_297# 0
C47319 _0607_/a_27_297# _0218_ 0
C47320 acc0.A\[20\] _0369_ 0.30405f
C47321 _0378_ net109 0
C47322 clknet_0__0457_ acc0.A\[20\] 0.07502f
C47323 hold25/a_391_47# _1041_/a_466_413# 0
C47324 _1028_/a_27_47# acc0.A\[28\] 0.00674f
C47325 hold31/a_285_47# _0252_ 0.06225f
C47326 _0343_ _0996_/a_1017_47# 0
C47327 _0723_/a_207_413# _0723_/a_297_47# 0.00476f
C47328 hold87/a_285_47# _0982_/a_1059_315# 0.00274f
C47329 hold42/a_49_47# _0187_ 0
C47330 _0443_ _0218_ 0.12464f
C47331 _1067_/a_891_413# control0.reset 0
C47332 _1057_/a_466_413# _0187_ 0.02324f
C47333 _1057_/a_891_413# net4 0
C47334 _0224_ net48 0.00234f
C47335 net220 _0460_ 0.01898f
C47336 _0812_/a_215_47# net217 0.08901f
C47337 _0812_/a_297_297# _0422_ 0.00282f
C47338 VPWR _0990_/a_381_47# 0.07359f
C47339 _0999_/a_891_413# _0096_ 0
C47340 _0999_/a_381_47# _0399_ 0
C47341 net85 _0783_/a_215_47# 0
C47342 VPWR _0793_/a_51_297# 0.50801f
C47343 hold28/a_49_47# net10 0
C47344 clknet_0__0462_ _0737_/a_117_297# 0.0017f
C47345 clkbuf_1_0__f__0459_/a_110_47# VPWR 1.23973f
C47346 VPWR _0564_/a_150_297# 0.00228f
C47347 net39 _0994_/a_27_47# 0.04414f
C47348 _0343_ net182 0
C47349 _0655_/a_109_93# clkbuf_1_1__f__0459_/a_110_47# 0
C47350 acc0.A\[16\] hold19/a_285_47# 0.0515f
C47351 _0557_/a_240_47# _1037_/a_891_413# 0
C47352 VPWR _0147_ 0.22786f
C47353 _1059_/a_193_47# acc0.A\[14\] 0.29026f
C47354 VPWR _0282_ 0.34967f
C47355 _0216_ net116 0.11135f
C47356 _0179_ _0190_ 0.00968f
C47357 net206 _0774_/a_68_297# 0
C47358 _0201_ _0540_/a_51_297# 0.00195f
C47359 _1041_/a_193_47# net7 0.05702f
C47360 hold59/a_391_47# _0181_ 0
C47361 hold97/a_49_47# _0318_ 0
C47362 hold4/a_391_47# _1022_/a_27_47# 0
C47363 hold4/a_285_47# _1022_/a_193_47# 0
C47364 hold4/a_49_47# _1022_/a_634_159# 0
C47365 _0636_/a_59_75# acc0.A\[3\] 0.08273f
C47366 _0090_ net228 0
C47367 _1017_/a_891_413# clknet_0__0461_ 0.01084f
C47368 _0460_ _1006_/a_592_47# 0
C47369 hold54/a_49_47# hold55/a_49_47# 0
C47370 _0742_/a_299_297# net52 0.01034f
C47371 _0532_/a_299_297# _1047_/a_891_413# 0
C47372 _0198_ _1047_/a_193_47# 0
C47373 _0764_/a_299_297# _0346_ 0.02782f
C47374 _1056_/a_27_47# input16/a_75_212# 0
C47375 _0170_ _1072_/a_1059_315# 0
C47376 _0753_/a_79_21# _0754_/a_149_47# 0
C47377 A[11] _0512_/a_109_297# 0.05359f
C47378 hold27/a_49_47# hold27/a_391_47# 0.00188f
C47379 VPWR _0166_ 0.39163f
C47380 net77 _0267_ 0.00192f
C47381 _0566_/a_27_47# _0526_/a_27_47# 0.0033f
C47382 clkload0/X _0183_ 0
C47383 hold23/a_49_47# hold23/a_285_47# 0.22264f
C47384 _1054_/a_193_47# VPWR 0.30029f
C47385 pp[27] hold80/a_285_47# 0
C47386 net149 _0264_ 0.14243f
C47387 net137 _0987_/a_634_159# 0
C47388 _1051_/a_193_47# _0085_ 0.00148f
C47389 clknet_1_0__leaf__0462_ _1025_/a_1059_315# 0
C47390 _1056_/a_381_47# VPWR 0.07542f
C47391 _0993_/a_1017_47# _0091_ 0
C47392 net122 net27 0
C47393 _0770_/a_382_297# _0389_ 0.01495f
C47394 _0770_/a_79_21# _0243_ 0.00139f
C47395 _0216_ hold92/a_285_47# 0.05641f
C47396 _0191_ acc0.A\[8\] 0
C47397 _1038_/a_27_47# VPWR 0.64771f
C47398 _0289_ clknet_1_1__leaf__0465_ 0.06051f
C47399 net61 _0350_ 0.00243f
C47400 _1041_/a_27_47# A[15] 0.00346f
C47401 _0248_ net52 0
C47402 _0742_/a_384_47# clknet_1_0__leaf__0460_ 0
C47403 _0767_/a_59_75# _0347_ 0
C47404 net36 clknet_1_0__leaf__0463_ 0.02284f
C47405 _1018_/a_634_159# acc0.A\[18\] 0.03558f
C47406 _0183_ _0576_/a_27_297# 0.19935f
C47407 _0217_ _0576_/a_109_47# 0.00171f
C47408 output58/a_27_47# acc0.A\[8\] 0
C47409 net189 _0181_ 0
C47410 _0247_ clknet_1_0__leaf__0457_ 0
C47411 _0387_ _0246_ 0
C47412 hold57/a_391_47# _1039_/a_891_413# 0
C47413 _0996_/a_592_47# net5 0.00178f
C47414 net114 _0347_ 0.09396f
C47415 clknet_0__0458_ _0257_ 0.00134f
C47416 clknet_0_clk _1068_/a_561_413# 0
C47417 net120 _1065_/a_27_47# 0
C47418 clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ 1.66521f
C47419 _0998_/a_592_47# net84 0.00107f
C47420 net105 clkbuf_0__0457_/a_110_47# 0.04316f
C47421 hold1/a_285_47# net148 0.00806f
C47422 pp[9] acc0.A\[9\] 0.00338f
C47423 clknet_1_0__leaf__0460_ _0379_ 0.00896f
C47424 _0159_ _0465_ 0
C47425 _0159_ _1061_/a_381_47# 0.11467f
C47426 hold30/a_285_47# hold30/a_391_47# 0.41909f
C47427 net110 acc0.A\[23\] 0.0915f
C47428 _0369_ _0988_/a_193_47# 0.00306f
C47429 acc0.A\[30\] net239 0
C47430 _0984_/a_1017_47# net47 0
C47431 _0372_ clknet_1_0__leaf__0460_ 0.23392f
C47432 _1001_/a_27_47# _0216_ 0
C47433 net190 acc0.A\[29\] 0.00959f
C47434 clknet_1_1__leaf__0463_ _0161_ 0
C47435 _1019_/a_381_47# net207 0.14614f
C47436 _0792_/a_303_47# net41 0
C47437 net35 _1071_/a_634_159# 0.0017f
C47438 _0965_/a_377_297# _0483_ 0.00282f
C47439 _0965_/a_285_47# control0.count\[3\] 0.03532f
C47440 _0539_/a_150_297# comp0.B\[12\] 0
C47441 net51 _1005_/a_381_47# 0
C47442 _0336_ _0334_ 0
C47443 _0694_/a_113_47# _0326_ 0.00937f
C47444 comp0.B\[13\] _1042_/a_27_47# 0.0016f
C47445 _0216_ hold8/a_49_47# 0
C47446 _0195_ hold8/a_391_47# 0.01267f
C47447 net155 hold8/a_285_47# 0.00977f
C47448 _0358_ acc0.A\[27\] 0
C47449 VPWR _0584_/a_373_47# 0
C47450 _0782_/a_27_47# _1014_/a_27_47# 0.00898f
C47451 _0760_/a_285_47# hold3/a_285_47# 0
C47452 _0082_ net146 0
C47453 _0312_ _0181_ 0
C47454 _0237_ _0373_ 0.17307f
C47455 _0233_ net50 0
C47456 _0343_ _0995_/a_634_159# 0.00362f
C47457 _1014_/a_466_413# clknet_1_0__leaf__0461_ 0.02309f
C47458 _0575_/a_109_297# net50 0
C47459 _0726_/a_51_297# _0109_ 0.10262f
C47460 _0726_/a_240_47# _0355_ 0.05299f
C47461 net144 net67 0
C47462 comp0.B\[1\] _1032_/a_27_47# 0.00131f
C47463 _0223_ net51 0.10238f
C47464 net242 _1010_/a_975_413# 0
C47465 _0287_ _0655_/a_369_297# 0
C47466 acc0.A\[1\] _0178_ 0.02371f
C47467 _0781_/a_68_297# _0459_ 0
C47468 _0753_/a_79_21# _0228_ 0
C47469 _0465_ _0447_ 0.01207f
C47470 _0800_/a_245_297# clknet_1_1__leaf__0459_ 0.00131f
C47471 net45 _0783_/a_215_47# 0.00415f
C47472 control0.state\[0\] _1064_/a_891_413# 0
C47473 net34 _1064_/a_466_413# 0.03264f
C47474 control0.state\[1\] _1064_/a_1059_315# 0
C47475 clkbuf_0__0465_/a_110_47# clkbuf_1_1__f__0458_/a_110_47# 0
C47476 _0996_/a_1059_315# clkbuf_1_1__f__0459_/a_110_47# 0
C47477 _0274_ _0826_/a_301_297# 0
C47478 _1033_/a_466_413# clknet_1_1__leaf__0463_ 0
C47479 input30/a_75_212# A[1] 0.00298f
C47480 B[7] input8/a_75_212# 0.00298f
C47481 _1015_/a_27_47# net157 0
C47482 hold86/a_391_47# net222 0
C47483 _0183_ _0891_/a_27_47# 0
C47484 _0381_ _0487_ 0
C47485 _0283_ hold81/a_285_47# 0.05217f
C47486 _0286_ hold81/a_49_47# 0.00253f
C47487 _1050_/a_634_159# _0148_ 0.00364f
C47488 hold46/a_285_47# net10 0.06832f
C47489 _1020_/a_193_47# _0181_ 0
C47490 _1001_/a_1059_315# _0247_ 0
C47491 net43 _0219_ 0.19376f
C47492 _0182_ _0112_ 0
C47493 _0179_ _0515_/a_299_297# 0.09747f
C47494 acc0.A\[2\] _0447_ 0
C47495 _0716_/a_27_47# _0296_ 0
C47496 clknet_0__0457_ _1001_/a_193_47# 0.00853f
C47497 net71 _0530_/a_299_297# 0.00246f
C47498 _1020_/a_1059_315# hold40/a_391_47# 0.01554f
C47499 _0467_ _1065_/a_193_47# 0.05293f
C47500 clknet_1_0__leaf__0465_ net73 0.02688f
C47501 _0347_ _0365_ 0.42664f
C47502 _0119_ _0578_/a_373_47# 0
C47503 _0216_ _1047_/a_193_47# 0
C47504 VPWR _0842_/a_59_75# 0.20809f
C47505 _0446_ _0847_/a_109_297# 0.00303f
C47506 _1014_/a_1059_315# net47 0
C47507 hold12/a_49_47# _0486_ 0
C47508 pp[28] hold80/a_49_47# 0.00329f
C47509 _0465_ _1048_/a_561_413# 0
C47510 _1048_/a_27_47# net147 0.00175f
C47511 _0089_ _0218_ 0.02058f
C47512 clknet_0__0459_ clknet_1_1__leaf__0465_ 0
C47513 _0176_ _0206_ 0.21016f
C47514 _0495_/a_150_297# _0173_ 0
C47515 _0514_/a_27_297# net66 0.0079f
C47516 _0244_ _0245_ 0.21148f
C47517 net152 net153 0
C47518 net32 net127 0
C47519 comp0.B\[5\] _1066_/a_193_47# 0
C47520 comp0.B\[3\] _1066_/a_466_413# 0
C47521 net88 _0460_ 0.0202f
C47522 _0999_/a_27_47# _0219_ 0.00238f
C47523 _0999_/a_1059_315# _0345_ 0.00247f
C47524 _0793_/a_245_297# _0407_ 0.00193f
C47525 _0322_ acc0.A\[26\] 0
C47526 hold83/a_285_47# _0150_ 0.00323f
C47527 acc0.A\[16\] _1017_/a_634_159# 0.00459f
C47528 _0234_ _0754_/a_51_297# 0.0802f
C47529 _0482_ hold89/a_391_47# 0
C47530 _1060_/a_27_47# _0505_/a_27_297# 0
C47531 net64 output58/a_27_47# 0.00755f
C47532 net31 comp0.B\[10\] 0.02212f
C47533 _0226_ _0381_ 0.12227f
C47534 _0211_ _1035_/a_466_413# 0
C47535 hold56/a_49_47# hold56/a_391_47# 0.00188f
C47536 _1050_/a_975_413# _0180_ 0.00107f
C47537 VPWR _0996_/a_193_47# 0.31417f
C47538 _0995_/a_193_47# net60 0
C47539 _0698_/a_113_297# _1008_/a_27_47# 0
C47540 _0647_/a_47_47# _0414_ 0
C47541 _1065_/a_193_47# comp0.B\[0\] 0.03286f
C47542 comp0.B\[7\] _1039_/a_561_413# 0
C47543 _0856_/a_79_21# _0850_/a_150_297# 0
C47544 _0216_ _0459_ 0.0396f
C47545 hold53/a_49_47# acc0.A\[25\] 0
C47546 net215 _0575_/a_27_297# 0.14453f
C47547 clknet_1_1__leaf__0460_ hold77/a_285_47# 0.02727f
C47548 _1037_/a_466_413# net28 0.00334f
C47549 _1034_/a_891_413# _0474_ 0.0036f
C47550 net237 _0319_ 0
C47551 clknet_1_0__leaf__0459_ _0793_/a_51_297# 0
C47552 _1051_/a_466_413# _1051_/a_592_47# 0.00553f
C47553 _1051_/a_634_159# _1051_/a_1017_47# 0
C47554 clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ 1.67652f
C47555 _1045_/a_466_413# _1044_/a_193_47# 0
C47556 _1045_/a_1059_315# _1044_/a_27_47# 0
C47557 _1045_/a_193_47# _1044_/a_466_413# 0
C47558 _1045_/a_634_159# _1044_/a_634_159# 0
C47559 net88 _0457_ 0
C47560 comp0.B\[14\] _1042_/a_891_413# 0
C47561 _0220_ _0704_/a_68_297# 0
C47562 _0227_ _1005_/a_466_413# 0
C47563 acc0.A\[21\] _1005_/a_1059_315# 0
C47564 _0368_ _0219_ 0.13639f
C47565 _0992_/a_1059_315# _0650_/a_68_297# 0.00151f
C47566 _1051_/a_193_47# net131 0
C47567 pp[27] _0220_ 0.01275f
C47568 net62 _0986_/a_193_47# 0.03661f
C47569 _1070_/a_592_47# control0.count\[1\] 0
C47570 VPWR _0168_ 0.50581f
C47571 _1045_/a_466_413# net131 0
C47572 _1045_/a_634_159# net184 0
C47573 _0467_ net33 0.17208f
C47574 hold56/a_391_47# _1032_/a_27_47# 0
C47575 hold56/a_285_47# _1032_/a_193_47# 0
C47576 net23 _1067_/a_466_413# 0.02902f
C47577 _1003_/a_634_159# net213 0
C47578 _0429_ clknet_0__0458_ 0
C47579 _1072_/a_193_47# clknet_1_0__leaf_clk 0.00433f
C47580 _0130_ net106 0.06804f
C47581 VPWR _1043_/a_592_47# 0
C47582 acc0.A\[8\] clkbuf_1_0__f__0465_/a_110_47# 0
C47583 acc0.A\[0\] _0465_ 0.00602f
C47584 _0618_/a_215_47# _0219_ 0.00409f
C47585 _0501_/a_27_47# net149 0
C47586 clknet_1_0__leaf__0458_ hold100/a_285_47# 0.00416f
C47587 _1038_/a_891_413# _0175_ 0
C47588 _0733_/a_222_93# _0322_ 0
C47589 VPWR clkbuf_0__0461_/a_110_47# 1.2643f
C47590 _1043_/a_634_159# net196 0.00122f
C47591 _1043_/a_466_413# net129 0
C47592 _0984_/a_27_47# _0158_ 0
C47593 hold32/a_285_47# net16 0.01654f
C47594 _1060_/a_27_47# _0506_/a_81_21# 0
C47595 VPWR _0568_/a_27_297# 0.29049f
C47596 VPWR _1015_/a_891_413# 0.18678f
C47597 clknet_1_0__leaf__0464_ _0146_ 0.00126f
C47598 _0195_ _0782_/a_27_47# 0.08223f
C47599 acc0.A\[21\] _0765_/a_79_21# 0.02066f
C47600 _0183_ _0346_ 0.24743f
C47601 net125 _1048_/a_27_47# 0
C47602 _0467_ hold12/a_391_47# 0.00299f
C47603 _0514_/a_27_297# _0350_ 0
C47604 clknet_1_0__leaf__0458_ _0982_/a_634_159# 0
C47605 _0579_/a_27_297# net1 0
C47606 acc0.A\[2\] acc0.A\[0\] 0
C47607 clkbuf_0__0464_/a_110_47# _0540_/a_240_47# 0
C47608 _1016_/a_27_47# hold72/a_285_47# 0
C47609 _1050_/a_1059_315# _0525_/a_81_21# 0
C47610 _0176_ _1046_/a_1059_315# 0
C47611 _0283_ _0282_ 0.15586f
C47612 control0.state\[0\] hold84/a_49_47# 0
C47613 VPWR _0654_/a_297_47# 0
C47614 _1030_/a_1059_315# _0128_ 0
C47615 clknet_1_1__leaf__0458_ _0825_/a_150_297# 0
C47616 _1021_/a_634_159# _0100_ 0
C47617 _1021_/a_466_413# net88 0.01755f
C47618 pp[25] output52/a_27_47# 0
C47619 _1032_/a_27_47# _1032_/a_634_159# 0.14145f
C47620 _0774_/a_68_297# _0774_/a_150_297# 0.00477f
C47621 _1054_/a_634_159# _1054_/a_592_47# 0
C47622 net9 _0522_/a_27_297# 0
C47623 net166 _0347_ 0
C47624 _1071_/a_381_47# control0.count\[0\] 0
C47625 net33 comp0.B\[0\] 0
C47626 _1015_/a_634_159# _1015_/a_381_47# 0
C47627 _0107_ clknet_1_1__leaf__0460_ 0.0401f
C47628 _0498_/a_51_297# _0173_ 0
C47629 _0983_/a_975_413# VPWR 0.0045f
C47630 _0358_ _1010_/a_193_47# 0.00267f
C47631 _0357_ _1010_/a_634_159# 0
C47632 _0096_ acc0.A\[17\] 0
C47633 _0557_/a_245_297# _0173_ 0.00103f
C47634 _0343_ net56 0
C47635 _0751_/a_111_297# _0227_ 0
C47636 comp0.B\[10\] net128 0
C47637 _0532_/a_81_21# net149 0.01159f
C47638 clknet_1_1__leaf__0462_ _1027_/a_381_47# 0.00315f
C47639 net113 _1027_/a_1059_315# 0
C47640 acc0.A\[12\] _0421_ 0
C47641 _0352_ _0773_/a_117_297# 0.00314f
C47642 net65 output63/a_27_47# 0.00589f
C47643 _0989_/a_466_413# output63/a_27_47# 0
C47644 _0792_/a_209_297# _0408_ 0.00295f
C47645 _0343_ _1031_/a_634_159# 0.00963f
C47646 _0216_ _0265_ 0
C47647 _0216_ clkbuf_1_0__f__0462_/a_110_47# 0
C47648 VPWR _0550_/a_245_297# 0.00524f
C47649 _0398_ clkbuf_1_1__f__0461_/a_110_47# 0.02109f
C47650 net247 _1047_/a_193_47# 0
C47651 net36 net165 0
C47652 _0319_ _0686_/a_27_53# 0
C47653 _1038_/a_1059_315# _1038_/a_891_413# 0.31086f
C47654 _1038_/a_193_47# _1038_/a_975_413# 0
C47655 _1038_/a_466_413# _1038_/a_381_47# 0.03733f
C47656 _1053_/a_466_413# _0180_ 0
C47657 _0211_ _1037_/a_27_47# 0
C47658 _0121_ _0757_/a_68_297# 0.00125f
C47659 _0829_/a_27_47# _0436_ 0.00471f
C47660 _0715_/a_27_47# _0084_ 0
C47661 _0319_ _1008_/a_891_413# 0
C47662 pp[20] VPWR 0.23729f
C47663 _1067_/a_193_47# clknet_1_0__leaf__0461_ 0.04228f
C47664 _0745_/a_193_47# _0370_ 0.01172f
C47665 net45 _0777_/a_377_297# 0
C47666 _0183_ _0629_/a_59_75# 0.001f
C47667 _0369_ net107 0
C47668 _0290_ _0812_/a_79_21# 0.0017f
C47669 net40 _0646_/a_47_47# 0.38836f
C47670 A[6] A[7] 0.18107f
C47671 pp[30] _0705_/a_145_75# 0
C47672 control0.state\[0\] _1065_/a_381_47# 0
C47673 clknet_1_0__leaf__0465_ _1044_/a_27_47# 0.00601f
C47674 clknet_1_1__leaf__0459_ _0995_/a_27_47# 0
C47675 _0983_/a_1059_315# _0983_/a_1017_47# 0
C47676 _0983_/a_193_47# net69 0.01434f
C47677 _0946_/a_30_53# _0468_ 0
C47678 clknet_1_0__leaf__0465_ _1051_/a_1017_47# 0
C47679 _0995_/a_891_413# input6/a_75_212# 0
C47680 net36 acc0.A\[19\] 0.00431f
C47681 _0401_ net228 0.23596f
C47682 _0346_ acc0.A\[15\] 0.0615f
C47683 net245 _0995_/a_1059_315# 0
C47684 net40 _0995_/a_381_47# 0
C47685 hold89/a_285_47# hold89/a_391_47# 0.41909f
C47686 _0659_/a_68_297# net66 0.12217f
C47687 net21 comp0.B\[12\] 0.1407f
C47688 net188 hold45/a_285_47# 0.0127f
C47689 _0984_/a_27_47# acc0.A\[14\] 0
C47690 hold69/a_49_47# VPWR 0.28234f
C47691 net71 _1049_/a_1059_315# 0
C47692 _0997_/a_27_47# net42 0.09308f
C47693 _0747_/a_79_21# _1006_/a_466_413# 0
C47694 acc0.A\[25\] _0687_/a_59_75# 0
C47695 _1056_/a_381_47# hold35/a_391_47# 0.00142f
C47696 _0466_ _1068_/a_891_413# 0.04625f
C47697 net90 _1007_/a_381_47# 0
C47698 _0318_ _0685_/a_150_297# 0
C47699 hold21/a_49_47# clknet_1_0__leaf__0465_ 0
C47700 _1048_/a_1059_315# _1047_/a_27_47# 0
C47701 _1048_/a_466_413# _1047_/a_193_47# 0
C47702 _1048_/a_634_159# _1047_/a_634_159# 0
C47703 _0851_/a_113_47# _0452_ 0
C47704 _0279_ _0276_ 0.00173f
C47705 _1003_/a_1017_47# _0217_ 0
C47706 _1004_/a_891_413# net50 0.02266f
C47707 _0935_/a_27_47# acc0.A\[15\] 0
C47708 clknet_1_0__leaf__0462_ _1005_/a_193_47# 0.00119f
C47709 _0553_/a_51_297# net28 0
C47710 _1061_/a_193_47# acc0.A\[15\] 0
C47711 net48 pp[20] 0.05148f
C47712 VPWR _0109_ 0.40843f
C47713 comp0.B\[2\] _0494_/a_27_47# 0.00205f
C47714 _0618_/a_79_21# acc0.A\[23\] 0
C47715 _0151_ _0180_ 0.00287f
C47716 _0629_/a_59_75# acc0.A\[15\] 0.01849f
C47717 _0998_/a_466_413# _0399_ 0.00346f
C47718 _0998_/a_634_159# _0096_ 0.02068f
C47719 _0216_ _0220_ 0.14804f
C47720 _0290_ _0347_ 0
C47721 hold17/a_285_47# _0168_ 0
C47722 hold87/a_391_47# _0080_ 0
C47723 _0476_ net203 0
C47724 _0780_/a_117_297# _0308_ 0.00795f
C47725 _0780_/a_35_297# _0306_ 0.00113f
C47726 net189 _0187_ 0.02544f
C47727 _0555_/a_240_47# _0176_ 0.0061f
C47728 _0350_ _0431_ 0
C47729 _0354_ _0568_/a_373_47# 0
C47730 clkbuf_0__0465_/a_110_47# _0291_ 0
C47731 clkbuf_1_0__f__0464_/a_110_47# net10 0.29425f
C47732 _0141_ hold51/a_285_47# 0
C47733 clknet_0__0458_ clknet_1_1__leaf__0458_ 0.3586f
C47734 _0559_/a_149_47# VPWR 0.00647f
C47735 _0179_ net192 0.22521f
C47736 _1008_/a_193_47# hold50/a_49_47# 0.00243f
C47737 _1008_/a_27_47# hold50/a_285_47# 0.00512f
C47738 _0216_ _0585_/a_109_297# 0.01376f
C47739 VPWR clkbuf_0__0462_/a_110_47# 1.20021f
C47740 _1052_/a_634_159# net154 0
C47741 _0961_/a_113_297# _0488_ 0.06461f
C47742 hold62/a_285_47# net209 0.01002f
C47743 _0982_/a_27_47# _1014_/a_27_47# 0
C47744 net247 _0265_ 0
C47745 _0985_/a_634_159# _0219_ 0
C47746 _0217_ _0634_/a_113_47# 0
C47747 hold54/a_285_47# comp0.B\[1\] 0.09364f
C47748 _0195_ _1017_/a_27_47# 0.42289f
C47749 net160 _1035_/a_1059_315# 0
C47750 clknet_1_1__leaf__0459_ _1057_/a_561_413# 0
C47751 hold64/a_285_47# _1001_/a_27_47# 0
C47752 _0179_ _0527_/a_109_297# 0.00869f
C47753 _0179_ _0346_ 0.05398f
C47754 _1016_/a_193_47# clknet_0__0461_ 0
C47755 _1057_/a_27_47# VPWR 0.66002f
C47756 net87 VPWR 0.38067f
C47757 comp0.B\[4\] _1034_/a_1059_315# 0.01431f
C47758 _1048_/a_27_47# _0186_ 0
C47759 _1052_/a_1059_315# _0252_ 0
C47760 hold33/a_285_47# net174 0.03146f
C47761 _0343_ _0345_ 0.11598f
C47762 VPWR B[6] 0.22365f
C47763 net44 acc0.A\[29\] 0.00334f
C47764 _1056_/a_381_47# net182 0.12224f
C47765 _0647_/a_47_47# _0404_ 0.0106f
C47766 acc0.A\[17\] _0395_ 0
C47767 _0179_ net65 0.00699f
C47768 _0179_ _0989_/a_466_413# 0
C47769 _0717_/a_209_297# _0705_/a_59_75# 0.00112f
C47770 _0734_/a_285_47# _1009_/a_466_413# 0
C47771 clknet_0_clk _0175_ 0
C47772 clknet_1_1__leaf__0465_ pp[4] 0
C47773 clknet_1_1__leaf__0459_ _0399_ 0.28792f
C47774 clknet_1_0__leaf__0459_ clkbuf_0__0461_/a_110_47# 0.0834f
C47775 net137 net73 0
C47776 clknet_1_0__leaf__0459_ _1015_/a_891_413# 0
C47777 _0174_ _0548_/a_512_297# 0
C47778 _0163_ _1065_/a_561_413# 0
C47779 _0513_/a_81_21# net192 0
C47780 _0188_ _0511_/a_299_297# 0
C47781 VPWR _0783_/a_215_47# 0.00122f
C47782 clknet_0__0458_ _0263_ 0.056f
C47783 _0256_ net170 0
C47784 _0953_/a_32_297# _0138_ 0
C47785 _0257_ _0837_/a_266_297# 0
C47786 _0500_/a_27_47# _0465_ 0.01935f
C47787 _0179_ _1061_/a_193_47# 0
C47788 net104 acc0.A\[18\] 0.08552f
C47789 _0989_/a_634_159# net75 0
C47790 net46 _0902_/a_27_47# 0
C47791 _0323_ clkbuf_1_0__f__0460_/a_110_47# 0
C47792 net35 _1072_/a_1059_315# 0.03212f
C47793 net114 _0106_ 0
C47794 _1067_/a_561_413# clknet_1_0__leaf__0457_ 0
C47795 _1067_/a_891_413# _0460_ 0.00104f
C47796 _0967_/a_109_93# _0468_ 0.00442f
C47797 hold10/a_49_47# _0181_ 0
C47798 _0690_/a_68_297# _0360_ 0
C47799 _0487_ _0468_ 0.42944f
C47800 hold21/a_391_47# A[4] 0.00389f
C47801 net22 _1061_/a_27_47# 0
C47802 _0783_/a_79_21# clkbuf_0__0461_/a_110_47# 0
C47803 _0172_ net135 0
C47804 _0473_ _0954_/a_220_297# 0
C47805 hold101/a_49_47# net62 0
C47806 net185 hold39/a_49_47# 0.0046f
C47807 _0323_ _0250_ 0.22166f
C47808 _0416_ _0276_ 0
C47809 _1059_/a_634_159# net41 0
C47810 _1020_/a_466_413# net118 0
C47811 _0760_/a_47_47# _0381_ 0.40994f
C47812 _0557_/a_240_47# net27 0.05798f
C47813 _0757_/a_150_297# _0350_ 0
C47814 _0757_/a_68_297# _0380_ 0.11118f
C47815 clknet_1_0__leaf__0458_ _0858_/a_27_47# 0
C47816 hold55/a_391_47# net187 0
C47817 _0286_ _0654_/a_207_413# 0.08527f
C47818 _1053_/a_193_47# _0152_ 0.00175f
C47819 _0326_ _0350_ 0
C47820 _0343_ hold16/a_49_47# 0
C47821 _1031_/a_1059_315# _1030_/a_1059_315# 0
C47822 _1031_/a_466_413# _1030_/a_891_413# 0
C47823 _0243_ _0617_/a_68_297# 0
C47824 _0457_ _1067_/a_891_413# 0
C47825 hold58/a_49_47# _0173_ 0.01284f
C47826 VPWR _0794_/a_326_47# 0.00137f
C47827 clknet_1_0__leaf__0463_ _1061_/a_27_47# 0.04463f
C47828 clknet_1_1__leaf__0460_ _0322_ 0.00821f
C47829 control0.state\[0\] _0471_ 0.16835f
C47830 _0962_/a_109_297# _0478_ 0.0031f
C47831 _1038_/a_27_47# net30 0
C47832 clknet_1_1__leaf__0460_ _0327_ 0.37142f
C47833 net160 _1037_/a_193_47# 0
C47834 _0712_/a_297_297# net60 0.01767f
C47835 _1025_/a_1059_315# _1025_/a_891_413# 0.31086f
C47836 _1025_/a_193_47# _1025_/a_975_413# 0
C47837 _1025_/a_466_413# _1025_/a_381_47# 0.03733f
C47838 _0458_ _0180_ 0.00433f
C47839 _0350_ hold95/a_391_47# 0
C47840 _0359_ _1006_/a_891_413# 0
C47841 _0324_ _1006_/a_1059_315# 0
C47842 _0292_ _0399_ 0.18025f
C47843 hold64/a_285_47# _0459_ 0.00846f
C47844 _0458_ net218 0
C47845 clkbuf_0__0465_/a_110_47# _0290_ 0
C47846 _0439_ acc0.A\[6\] 0
C47847 net58 _0627_/a_369_297# 0
C47848 hold5/a_285_47# _1042_/a_27_47# 0.00129f
C47849 rst clknet_1_0__leaf_clk 0
C47850 _0131_ clknet_1_1__leaf__0463_ 0.0417f
C47851 _0982_/a_27_47# _0195_ 0
C47852 _0113_ _0584_/a_373_47# 0
C47853 _1055_/a_891_413# _0181_ 0
C47854 _0410_ hold91/a_391_47# 0
C47855 VPWR acc0.A\[6\] 3.09582f
C47856 net136 _0148_ 0
C47857 control0.count\[1\] _0976_/a_76_199# 0.06242f
C47858 _1070_/a_381_47# _0488_ 0
C47859 _1070_/a_891_413# _0466_ 0
C47860 VPWR _0976_/a_439_47# 0
C47861 net178 clknet_1_1__leaf__0458_ 0.04396f
C47862 hold100/a_391_47# _0856_/a_79_21# 0
C47863 hold38/a_49_47# control0.reset 0
C47864 net248 _0625_/a_59_75# 0.0692f
C47865 _0369_ _0772_/a_297_297# 0.00457f
C47866 hold54/a_285_47# _1032_/a_634_159# 0
C47867 hold54/a_49_47# _1032_/a_466_413# 0
C47868 _0365_ _0106_ 0.06229f
C47869 _1046_/a_975_413# net10 0.00208f
C47870 clknet_1_1__leaf__0459_ _0808_/a_266_297# 0.0017f
C47871 _0955_/a_32_297# _0215_ 0
C47872 _0982_/a_466_413# _0856_/a_79_21# 0
C47873 _0982_/a_193_47# _0856_/a_215_47# 0.00119f
C47874 _0972_/a_93_21# _1063_/a_27_47# 0.00287f
C47875 net38 _0808_/a_266_47# 0
C47876 _0763_/a_193_47# _0373_ 0
C47877 _0403_ _0994_/a_634_159# 0
C47878 clknet_0__0463_ _1061_/a_466_413# 0
C47879 _0195_ _0145_ 0
C47880 _0533_/a_109_297# comp0.B\[15\] 0.00758f
C47881 net233 clknet_1_0__leaf__0458_ 0
C47882 net206 _0264_ 0.05726f
C47883 _1003_/a_381_47# control0.state\[2\] 0
C47884 hold18/a_391_47# _0446_ 0.03137f
C47885 hold18/a_285_47# _0450_ 0
C47886 hold58/a_285_47# _0212_ 0.02456f
C47887 hold58/a_391_47# net185 0
C47888 _0216_ net51 0.01306f
C47889 _0996_/a_634_159# _0996_/a_592_47# 0
C47890 _0539_/a_68_297# _0203_ 0
C47891 _1055_/a_466_413# _0517_/a_81_21# 0.00453f
C47892 hold59/a_49_47# net104 0.03504f
C47893 net203 clkbuf_0__0463_/a_110_47# 0
C47894 _0388_ _0347_ 0.00311f
C47895 net45 _1031_/a_1059_315# 0.00112f
C47896 _0189_ net66 0.46149f
C47897 clknet_0__0463_ net171 0
C47898 _1066_/a_27_47# hold84/a_285_47# 0.00178f
C47899 _1066_/a_193_47# hold84/a_49_47# 0.00209f
C47900 input15/a_75_212# net11 0
C47901 hold64/a_391_47# clknet_1_0__leaf__0461_ 0.01772f
C47902 _0080_ _0264_ 0
C47903 _0294_ _0679_/a_150_297# 0.00122f
C47904 clknet_1_0__leaf__0464_ _1048_/a_381_47# 0
C47905 hold53/a_49_47# net210 0
C47906 clknet_1_1__leaf__0457_ _1061_/a_1059_315# 0.01157f
C47907 _0518_/a_27_297# _0369_ 0
C47908 net7 comp0.B\[10\] 0.02009f
C47909 acc0.A\[16\] net103 0.17453f
C47910 _0976_/a_505_21# clkbuf_1_0__f_clk/a_110_47# 0.00164f
C47911 _0375_ _0377_ 0.01817f
C47912 _0234_ _0219_ 0.11474f
C47913 _0376_ _0345_ 0.12181f
C47914 _1060_/a_27_47# _0184_ 0
C47915 _1060_/a_634_159# net6 0
C47916 _0732_/a_303_47# _0219_ 0
C47917 _0559_/a_51_297# _0559_/a_240_47# 0.03076f
C47918 _0714_/a_51_297# _0341_ 0.09462f
C47919 _0211_ _0133_ 0
C47920 _0317_ _0686_/a_301_297# 0
C47921 hold42/a_49_47# clknet_1_1__leaf__0465_ 0.03193f
C47922 _0701_/a_80_21# clknet_1_1__leaf__0462_ 0.00766f
C47923 hold70/a_49_47# net228 0.14266f
C47924 clknet_1_0__leaf__0463_ _1039_/a_27_47# 0.00412f
C47925 _1057_/a_466_413# clknet_1_1__leaf__0465_ 0.01393f
C47926 VPWR _1036_/a_634_159# 0.18069f
C47927 _0344_ _0999_/a_891_413# 0
C47928 clknet_0__0457_ _0208_ 0
C47929 hold24/a_285_47# _0174_ 0.0192f
C47930 comp0.B\[7\] _0553_/a_240_47# 0
C47931 _1044_/a_27_47# _1044_/a_466_413# 0.27314f
C47932 _1044_/a_193_47# _1044_/a_634_159# 0.11072f
C47933 _0251_ _0274_ 0.04855f
C47934 _0274_ _0640_/a_109_53# 0.00643f
C47935 _0275_ _0640_/a_215_297# 0
C47936 VPWR _0725_/a_80_21# 0.15428f
C47937 VPWR _0523_/a_384_47# 0
C47938 clknet_0__0463_ net24 0.0117f
C47939 _0329_ clkbuf_1_1__f__0462_/a_110_47# 0.03588f
C47940 _1051_/a_27_47# net130 0
C47941 net137 _1044_/a_27_47# 0
C47942 _0135_ net28 0.28999f
C47943 _0815_/a_113_297# _0815_/a_199_47# 0
C47944 hold65/a_391_47# _0437_ 0.00138f
C47945 hold65/a_49_47# _0087_ 0
C47946 _1051_/a_381_47# acc0.A\[5\] 0
C47947 _0174_ input7/a_75_212# 0
C47948 net131 _1044_/a_634_159# 0
C47949 net184 _1044_/a_193_47# 0
C47950 _0222_ _0373_ 0
C47951 net237 _0250_ 0
C47952 _0227_ _0103_ 0.03262f
C47953 net247 _0267_ 0
C47954 _1021_/a_27_47# _0764_/a_81_21# 0
C47955 _0441_ _0346_ 0.00339f
C47956 clknet_0__0460_ _0219_ 0.05767f
C47957 VPWR _0777_/a_377_297# 0.00615f
C47958 output43/a_27_47# net42 0.00169f
C47959 net131 net184 0.17111f
C47960 _0269_ _0350_ 0.05143f
C47961 clknet_1_1__leaf__0459_ _0299_ 0.01972f
C47962 _0399_ _0990_/a_975_413# 0.00174f
C47963 _0319_ _0320_ 0.16496f
C47964 net46 _1023_/a_193_47# 0.00819f
C47965 output46/a_27_47# _1023_/a_1059_315# 0.00124f
C47966 control0.state\[0\] hold93/a_391_47# 0
C47967 control0.state\[1\] hold93/a_285_47# 0.00606f
C47968 hold49/a_49_47# _0540_/a_149_47# 0
C47969 clknet_1_0__leaf__0459_ net87 0.16569f
C47970 _0789_/a_544_297# VPWR 0.0083f
C47971 _0275_ _0465_ 0.01003f
C47972 acc0.A\[28\] _0350_ 0.02576f
C47973 net40 _0219_ 0
C47974 clknet_1_1__leaf__0459_ _0295_ 0.0019f
C47975 net129 net196 0.00532f
C47976 _1039_/a_466_413# clknet_0__0463_ 0.01118f
C47977 _0714_/a_240_47# _1013_/a_193_47# 0
C47978 clkbuf_1_1__f__0462_/a_110_47# _0221_ 0
C47979 VPWR _0128_ 0.20192f
C47980 _0343_ net52 0.23912f
C47981 clknet_1_1__leaf__0460_ _0306_ 0.00146f
C47982 _0189_ _0350_ 0
C47983 input29/a_75_212# net29 0.10849f
C47984 clknet_1_0__leaf__0458_ net68 0.12551f
C47985 pp[8] output47/a_27_47# 0.0119f
C47986 VPWR _0673_/a_253_297# 0.0015f
C47987 _0343_ _0819_/a_81_21# 0.03301f
C47988 _1030_/a_381_47# _0345_ 0.0022f
C47989 clknet_0__0464_ net20 0.056f
C47990 _0350_ net209 0
C47991 _1072_/a_466_413# net159 0
C47992 VPWR _0672_/a_297_297# 0.00952f
C47993 _0627_/a_109_93# clknet_1_1__leaf__0458_ 0.00253f
C47994 hold76/a_49_47# _1000_/a_1059_315# 0
C47995 _0972_/a_250_297# _1062_/a_466_413# 0
C47996 _0849_/a_79_21# _0849_/a_510_47# 0.00844f
C47997 _0849_/a_297_297# _0849_/a_215_47# 0
C47998 hold101/a_391_47# _0987_/a_27_47# 0
C47999 _0119_ net88 0.25867f
C48000 _1032_/a_891_413# _1032_/a_975_413# 0.00851f
C48001 _1032_/a_381_47# _1032_/a_561_413# 0.00123f
C48002 net9 _0193_ 0
C48003 pp[15] hold98/a_285_47# 0.0278f
C48004 _0568_/a_109_297# net208 0.01151f
C48005 _0251_ pp[5] 0
C48006 _0198_ _0178_ 0
C48007 _1015_/a_891_413# _0113_ 0.03672f
C48008 pp[12] output40/a_27_47# 0.01004f
C48009 net77 _0347_ 0.03158f
C48010 net175 net71 0.14756f
C48011 _0624_/a_59_75# VPWR 0.22451f
C48012 _1051_/a_891_413# _0180_ 0
C48013 _0575_/a_27_297# clknet_1_0__leaf__0460_ 0
C48014 _0852_/a_35_297# _0446_ 0.00841f
C48015 net100 _0585_/a_109_297# 0
C48016 _1014_/a_466_413# _0112_ 0
C48017 _0769_/a_384_47# _0773_/a_35_297# 0
C48018 _0783_/a_79_21# _0783_/a_215_47# 0.04584f
C48019 _1038_/a_381_47# net172 0.13436f
C48020 net33 _1066_/a_381_47# 0.0208f
C48021 hold21/a_285_47# hold21/a_391_47# 0.41909f
C48022 net220 _0373_ 0
C48023 _0456_ _0399_ 0
C48024 clknet_0__0459_ _0277_ 0
C48025 net242 _0701_/a_80_21# 0
C48026 net1 net33 0
C48027 _0476_ _0176_ 0.16609f
C48028 _0343_ _1055_/a_27_47# 0.03877f
C48029 _0366_ _0460_ 0
C48030 _0401_ _0090_ 0
C48031 hold25/a_49_47# comp0.B\[8\] 0
C48032 _0343_ _0791_/a_113_297# 0.03676f
C48033 _0750_/a_181_47# _0383_ 0
C48034 _0268_ net222 0
C48035 control0.count\[2\] _0976_/a_505_21# 0
C48036 _0536_/a_51_297# _0159_ 0
C48037 hold81/a_285_47# _0345_ 0.01086f
C48038 net168 _1052_/a_193_47# 0
C48039 _0292_ _0295_ 0
C48040 _0997_/a_891_413# net43 0.03879f
C48041 _0352_ _1006_/a_193_47# 0.03377f
C48042 _0656_/a_59_75# _0347_ 0.04609f
C48043 _0267_ _0841_/a_79_21# 0
C48044 VPWR _0995_/a_1059_315# 0.41769f
C48045 pp[1] _0988_/a_27_47# 0
C48046 output47/a_27_47# _0988_/a_891_413# 0
C48047 _0432_ clkbuf_1_1__f__0458_/a_110_47# 0.00118f
C48048 _0289_ _0296_ 0
C48049 _0284_ _0993_/a_193_47# 0.00652f
C48050 _0195_ _0245_ 0
C48051 _0983_/a_891_413# acc0.A\[18\] 0
C48052 _0212_ _0134_ 0
C48053 _0520_/a_27_297# _0179_ 0.02859f
C48054 net61 hold101/a_285_47# 0
C48055 net72 _0084_ 0
C48056 net45 _0712_/a_561_47# 0
C48057 _0384_ _0099_ 0
C48058 _0225_ _0754_/a_240_47# 0.00187f
C48059 _0433_ _0830_/a_79_21# 0
C48060 hold87/a_49_47# _0350_ 0.00136f
C48061 hold13/a_391_47# net28 0
C48062 _0511_/a_384_47# _0187_ 0
C48063 A[1] _0176_ 0
C48064 clknet_1_0__leaf__0465_ _0196_ 0
C48065 _0352_ acc0.A\[25\] 0.02963f
C48066 _1051_/a_193_47# _0525_/a_81_21# 0
C48067 hold28/a_285_47# _1048_/a_891_413# 0.00152f
C48068 hold28/a_391_47# _1048_/a_1059_315# 0
C48069 pp[16] acc0.A\[31\] 0.00131f
C48070 _0217_ clknet_1_0__leaf__0457_ 0.40645f
C48071 _0230_ _0232_ 0.16268f
C48072 _0550_/a_51_297# _0172_ 0.14086f
C48073 hold23/a_285_47# net170 0.05594f
C48074 _0550_/a_245_297# net30 0
C48075 net216 _1006_/a_561_413# 0
C48076 _0662_/a_81_21# _0275_ 0
C48077 _1013_/a_466_413# net41 0
C48078 _0104_ _1006_/a_1059_315# 0
C48079 net190 _1008_/a_1059_315# 0
C48080 _0533_/a_27_297# _0533_/a_373_47# 0.01338f
C48081 _0179_ clkbuf_0__0464_/a_110_47# 0.00119f
C48082 _0354_ _0725_/a_303_47# 0
C48083 _0355_ _0725_/a_209_47# 0.00117f
C48084 acc0.A\[12\] _1058_/a_592_47# 0.00289f
C48085 _0349_ _0730_/a_79_21# 0
C48086 hold71/a_49_47# hold71/a_285_47# 0.22264f
C48087 hold14/a_49_47# _0211_ 0.06021f
C48088 _1000_/a_891_413# _0461_ 0.00608f
C48089 _0186_ _0524_/a_373_47# 0.00246f
C48090 comp0.B\[11\] comp0.B\[10\] 0.04115f
C48091 VPWR comp0.B\[5\] 1.42985f
C48092 net168 net12 0.03125f
C48093 net187 _0352_ 0.11079f
C48094 _0608_/a_27_47# _0218_ 0
C48095 _0195_ hold9/a_285_47# 0.03192f
C48096 _0546_/a_245_297# _0546_/a_240_47# 0
C48097 _0247_ _0246_ 0.06626f
C48098 _1047_/a_27_47# clkbuf_1_1__f__0457_/a_110_47# 0.01976f
C48099 VPWR _1023_/a_634_159# 0.18293f
C48100 hold100/a_391_47# _0846_/a_51_297# 0
C48101 _1036_/a_561_413# _0175_ 0
C48102 _0746_/a_81_21# clknet_0__0460_ 0
C48103 _0534_/a_81_21# _0199_ 0.18217f
C48104 _0991_/a_634_159# _0991_/a_1059_315# 0
C48105 _0991_/a_27_47# _0991_/a_381_47# 0.06222f
C48106 _0991_/a_193_47# _0991_/a_891_413# 0.19685f
C48107 net84 _0096_ 0.16255f
C48108 _0210_ _0561_/a_51_297# 0
C48109 comp0.B\[4\] _0209_ 0
C48110 _0397_ _0394_ 0.037f
C48111 _0216_ _0178_ 0.10217f
C48112 _0243_ acc0.A\[18\] 0
C48113 _1041_/a_466_413# net22 0
C48114 hold19/a_391_47# _0184_ 0
C48115 _0747_/a_79_21# _0369_ 0.12204f
C48116 _0773_/a_117_297# _0392_ 0
C48117 _0195_ _1029_/a_193_47# 0
C48118 _0146_ clkbuf_1_0__f__0464_/a_110_47# 0
C48119 acc0.A\[12\] _0186_ 0.50473f
C48120 acc0.A\[19\] hold60/a_391_47# 0
C48121 _1052_/a_1017_47# net11 0
C48122 net101 _0526_/a_27_47# 0
C48123 _0793_/a_51_297# _0345_ 0.20904f
C48124 clknet_1_1__leaf__0459_ _0811_/a_299_297# 0.00177f
C48125 hold64/a_285_47# _0772_/a_79_21# 0
C48126 _1001_/a_634_159# _0183_ 0
C48127 hold6/a_285_47# _1040_/a_466_413# 0
C48128 clknet_1_0__leaf__0463_ _1037_/a_27_47# 0.00776f
C48129 _0399_ _0996_/a_466_413# 0.02328f
C48130 _0574_/a_109_297# acc0.A\[25\] 0.02002f
C48131 net45 _0611_/a_68_297# 0
C48132 _0282_ _0345_ 0
C48133 clknet_1_1__leaf__0460_ _0346_ 0.0277f
C48134 _0800_/a_51_297# _0297_ 0
C48135 _0226_ _0762_/a_79_21# 0
C48136 _0808_/a_81_21# _0418_ 0.22718f
C48137 _1021_/a_193_47# _0217_ 0.02828f
C48138 _1041_/a_466_413# clknet_1_0__leaf__0463_ 0.00579f
C48139 hold35/a_285_47# _0154_ 0.00315f
C48140 _0854_/a_297_297# _0347_ 0.00324f
C48141 _0573_/a_27_47# _0145_ 0
C48142 clkbuf_1_1__f__0461_/a_110_47# _0308_ 0
C48143 _0731_/a_299_297# _0326_ 0.01334f
C48144 _0840_/a_68_297# _0840_/a_150_297# 0.00477f
C48145 net130 _0085_ 0
C48146 _0125_ hold9/a_391_47# 0
C48147 acc0.A\[20\] hold40/a_391_47# 0.07318f
C48148 clknet_0__0458_ _0642_/a_27_413# 0
C48149 _0665_/a_109_297# _0298_ 0
C48150 clknet_0__0461_ _0773_/a_285_297# 0
C48151 _1058_/a_466_413# acc0.A\[10\] 0
C48152 hold44/a_391_47# _0354_ 0
C48153 _1067_/a_466_413# _0161_ 0
C48154 _0366_ _1007_/a_1017_47# 0.00118f
C48155 _0391_ _0771_/a_27_413# 0.04241f
C48156 _0446_ _0846_/a_149_47# 0.00369f
C48157 comp0.B\[10\] _0202_ 0
C48158 net223 _0771_/a_215_297# 0
C48159 _0174_ _0138_ 0
C48160 _0600_/a_103_199# _0350_ 0.00122f
C48161 _0218_ _0841_/a_297_297# 0
C48162 _0619_/a_68_297# _0435_ 0.00839f
C48163 _0478_ _0471_ 0
C48164 _0258_ _0442_ 0
C48165 _0522_/a_109_297# net13 0.01056f
C48166 clkbuf_1_1__f__0460_/a_110_47# clknet_0__0462_ 0.01649f
C48167 _0722_/a_215_47# _0352_ 0.01034f
C48168 _0800_/a_51_297# _0412_ 0.08187f
C48169 clkbuf_1_1__f__0457_/a_110_47# clknet_1_0__leaf__0461_ 0
C48170 VPWR _0601_/a_150_297# 0.00213f
C48171 _0663_/a_207_413# _0663_/a_297_47# 0.00476f
C48172 _0148_ net73 0.00229f
C48173 net216 clkbuf_0__0460_/a_110_47# 0.00169f
C48174 _0425_ _0291_ 0
C48175 clkbuf_0__0463_/a_110_47# _0176_ 0.01772f
C48176 VPWR _0697_/a_472_297# 0.00419f
C48177 _1002_/a_891_413# _0352_ 0.0024f
C48178 net167 _1068_/a_634_159# 0
C48179 _0304_ _0303_ 0.03173f
C48180 _0996_/a_1059_315# _0277_ 0
C48181 VPWR _0331_ 0.42145f
C48182 VPWR _0695_/a_300_47# 0.00101f
C48183 hold29/a_285_47# _1023_/a_891_413# 0
C48184 hold29/a_391_47# _1023_/a_1059_315# 0
C48185 _0483_ _0488_ 0.25776f
C48186 _1004_/a_466_413# net52 0.00237f
C48187 VPWR _1031_/a_1059_315# 0.40998f
C48188 _0118_ net118 0
C48189 clkbuf_0__0465_/a_110_47# _0986_/a_1059_315# 0.01586f
C48190 _0295_ _0655_/a_215_53# 0
C48191 _0216_ _1019_/a_27_47# 0
C48192 net178 _0988_/a_1017_47# 0
C48193 net39 _0648_/a_27_297# 0
C48194 _0183_ net221 0.05113f
C48195 _0296_ _0655_/a_109_93# 0
C48196 _0289_ _0811_/a_81_21# 0.00994f
C48197 _0423_ _0991_/a_891_413# 0
C48198 _0401_ _0991_/a_466_413# 0
C48199 net180 net29 0
C48200 _1043_/a_27_47# hold51/a_285_47# 0.00123f
C48201 net56 _0568_/a_27_297# 0.01159f
C48202 _0983_/a_1017_47# _0399_ 0.00161f
C48203 hold68/a_285_47# net50 0.07574f
C48204 _0248_ clknet_1_0__leaf__0457_ 0.00257f
C48205 _0515_/a_384_47# acc0.A\[11\] 0
C48206 net215 net176 0
C48207 clkbuf_1_0__f__0458_/a_110_47# _0446_ 0.00249f
C48208 clknet_0__0458_ _0848_/a_27_47# 0
C48209 _0217_ _0850_/a_68_297# 0
C48210 control0.state\[2\] clknet_1_0__leaf_clk 0
C48211 _0955_/a_32_297# _0955_/a_304_297# 0.00167f
C48212 hold76/a_391_47# _0242_ 0.0074f
C48213 hold15/a_285_47# _0336_ 0.00125f
C48214 hold15/a_391_47# _0220_ 0.02188f
C48215 net53 _0696_/a_109_297# 0.00262f
C48216 net7 _0177_ 0
C48217 hold44/a_285_47# _0569_/a_27_297# 0.00104f
C48218 _0216_ _0324_ 0.00776f
C48219 _0991_/a_27_47# _0082_ 0
C48220 _1004_/a_1059_315# clknet_1_0__leaf__0460_ 0.00377f
C48221 _0523_/a_81_21# acc0.A\[6\] 0.02183f
C48222 clknet_0__0458_ _0218_ 0.40582f
C48223 _0344_ net60 0
C48224 _1025_/a_466_413# acc0.A\[25\] 0.02307f
C48225 _0178_ net247 0.02183f
C48226 _1020_/a_27_47# _1015_/a_193_47# 0.00123f
C48227 _1020_/a_193_47# _1015_/a_27_47# 0
C48228 _0971_/a_81_21# clknet_1_0__leaf__0457_ 0.00166f
C48229 control0.reset _0565_/a_51_297# 0
C48230 hold65/a_391_47# _0252_ 0
C48231 net54 _1008_/a_193_47# 0.00927f
C48232 net39 output39/a_27_47# 0.1829f
C48233 control0.count\[1\] _0488_ 0.34756f
C48234 _1001_/a_891_413# control0.add 0.00108f
C48235 hold20/a_391_47# _1072_/a_193_47# 0
C48236 clkbuf_1_0__f__0457_/a_110_47# _1019_/a_1059_315# 0
C48237 clknet_0__0457_ _1019_/a_193_47# 0.02385f
C48238 _0709_/a_113_47# net60 0
C48239 _0243_ net211 0.00285f
C48240 _0211_ _0208_ 0.34854f
C48241 _0474_ _0215_ 0
C48242 clknet_1_1__leaf__0459_ _0091_ 0.00298f
C48243 _0080_ _0856_/a_79_21# 0.05051f
C48244 net231 _1063_/a_27_47# 0.00115f
C48245 pp[27] _0347_ 0
C48246 _0119_ _1067_/a_891_413# 0
C48247 _1021_/a_634_159# control0.add 0
C48248 hold63/a_285_47# _0572_/a_27_297# 0.00152f
C48249 _0684_/a_59_75# _1009_/a_1059_315# 0
C48250 net22 _0953_/a_32_297# 0
C48251 _1036_/a_27_47# _1036_/a_634_159# 0.14145f
C48252 _0422_ hold70/a_391_47# 0.06796f
C48253 _1047_/a_466_413# acc0.A\[15\] 0
C48254 _1012_/a_27_47# clknet_1_1__leaf__0462_ 0
C48255 _0769_/a_81_21# _0244_ 0.19845f
C48256 _0330_ clknet_1_1__leaf__0462_ 0.60508f
C48257 _0402_ _0993_/a_381_47# 0
C48258 net168 pp[5] 0
C48259 _0082_ _0350_ 0
C48260 _0217_ hold19/a_285_47# 0
C48261 _0993_/a_634_159# _0218_ 0.00135f
C48262 _1049_/a_27_47# net154 0
C48263 _0108_ _0685_/a_68_297# 0.01129f
C48264 _0191_ _0369_ 0
C48265 hold68/a_49_47# net215 0
C48266 _0523_/a_81_21# _0523_/a_384_47# 0.00138f
C48267 _0466_ clkbuf_1_0__f_clk/a_110_47# 0.12035f
C48268 comp0.B\[6\] input29/a_75_212# 0
C48269 _0662_/a_384_47# _0181_ 0
C48270 net146 net6 0.06524f
C48271 hold101/a_391_47# clkbuf_1_0__f__0465_/a_110_47# 0.01103f
C48272 hold27/a_49_47# _0498_/a_51_297# 0
C48273 net226 _0978_/a_27_297# 0.12008f
C48274 net225 _0341_ 0.12138f
C48275 net217 net67 0.03181f
C48276 _1041_/a_1059_315# _0544_/a_51_297# 0
C48277 _1041_/a_27_47# _0544_/a_240_47# 0
C48278 net189 clknet_1_1__leaf__0465_ 0.43473f
C48279 output58/a_27_47# _0369_ 0
C48280 net36 control0.sh 0
C48281 _1050_/a_891_413# _0524_/a_27_297# 0
C48282 A[15] net153 0
C48283 pp[16] net43 0.00675f
C48284 A[11] net67 0.00414f
C48285 _1059_/a_466_413# clkbuf_0__0459_/a_110_47# 0.00231f
C48286 clknet_1_0__leaf__0463_ _0953_/a_32_297# 0.03983f
C48287 _0238_ _0616_/a_78_199# 0
C48288 _1044_/a_193_47# net130 0.00337f
C48289 _1044_/a_1059_315# _1044_/a_1017_47# 0
C48290 _0403_ _0787_/a_80_21# 0.07779f
C48291 _0178_ _1048_/a_466_413# 0
C48292 _1065_/a_27_47# _0175_ 0
C48293 hold46/a_391_47# comp0.B\[12\] 0
C48294 _0529_/a_27_297# _0529_/a_373_47# 0.01338f
C48295 _0275_ _0254_ 0
C48296 hold33/a_285_47# hold46/a_49_47# 0
C48297 _0606_/a_109_53# _0383_ 0
C48298 _1038_/a_975_413# comp0.B\[6\] 0.00265f
C48299 net188 _1058_/a_27_47# 0
C48300 _0996_/a_193_47# _0345_ 0
C48301 hold49/a_285_47# _0542_/a_51_297# 0
C48302 _0460_ acc0.A\[24\] 0.00421f
C48303 _0290_ _0425_ 0.10018f
C48304 _0683_/a_113_47# _0313_ 0
C48305 net131 net130 0.01505f
C48306 _0682_/a_68_297# _1007_/a_27_47# 0
C48307 _1058_/a_1059_315# _0510_/a_27_297# 0.01884f
C48308 _0804_/a_79_21# net39 0.0211f
C48309 input20/a_75_212# input19/a_75_212# 0
C48310 _0172_ _0913_/a_27_47# 0.00334f
C48311 _0946_/a_30_53# _0978_/a_109_297# 0
C48312 net36 _1038_/a_466_413# 0.03138f
C48313 pp[0] _1038_/a_193_47# 0.00134f
C48314 clknet_1_1__leaf_clk _1065_/a_891_413# 0.04727f
C48315 _1049_/a_27_47# _0465_ 0
C48316 _0343_ hold94/a_391_47# 0
C48317 _0368_ _1007_/a_193_47# 0
C48318 _0985_/a_466_413# acc0.A\[2\] 0
C48319 _0819_/a_81_21# _0990_/a_381_47# 0
C48320 _0237_ _1005_/a_466_413# 0
C48321 _0585_/a_27_297# clkbuf_1_1__f__0457_/a_110_47# 0.00846f
C48322 VPWR B[3] 0.27647f
C48323 output55/a_27_47# _0356_ 0
C48324 pp[19] _1023_/a_1017_47# 0
C48325 _0195_ _1028_/a_381_47# 0.01652f
C48326 _0216_ _1028_/a_1059_315# 0.00243f
C48327 _1067_/a_592_47# net17 0
C48328 hold42/a_285_47# hold42/a_391_47# 0.41909f
C48329 net56 _0109_ 0
C48330 _0467_ _0880_/a_27_47# 0.00205f
C48331 hold42/a_285_47# _1057_/a_891_413# 0
C48332 net49 _0369_ 0.02298f
C48333 net57 _0723_/a_27_413# 0.00487f
C48334 _0744_/a_27_47# net67 0
C48335 _1051_/a_1017_47# _0148_ 0
C48336 _1057_/a_1059_315# _1057_/a_891_413# 0.31086f
C48337 _1057_/a_193_47# _1057_/a_975_413# 0
C48338 _1057_/a_466_413# _1057_/a_381_47# 0.03733f
C48339 VPWR _0377_ 0.26302f
C48340 acc0.A\[2\] _1049_/a_27_47# 0
C48341 _0553_/a_51_297# clknet_0__0463_ 0
C48342 B[13] _1042_/a_634_159# 0
C48343 _0269_ _0986_/a_634_159# 0
C48344 _0984_/a_193_47# _0991_/a_27_47# 0
C48345 _0984_/a_27_47# _0991_/a_193_47# 0
C48346 _0111_ _1013_/a_466_413# 0.03229f
C48347 VPWR _1064_/a_891_413# 0.19844f
C48348 _0174_ net134 0
C48349 _0454_ net206 0
C48350 net236 clkbuf_1_0__f_clk/a_110_47# 0.00196f
C48351 _0334_ hold95/a_285_47# 0.00318f
C48352 _0789_/a_75_199# _0789_/a_544_297# 0.01759f
C48353 _0501_/a_27_47# comp0.B\[15\] 0.00801f
C48354 net199 pp[24] 0
C48355 _1059_/a_466_413# _1059_/a_381_47# 0.03733f
C48356 _1059_/a_193_47# _1059_/a_975_413# 0
C48357 _1059_/a_1059_315# _1059_/a_891_413# 0.31086f
C48358 hold59/a_285_47# _0266_ 0.00102f
C48359 _1004_/a_891_413# _0576_/a_27_297# 0
C48360 _1004_/a_1059_315# _0576_/a_109_297# 0
C48361 net55 pp[28] 0
C48362 net231 _1062_/a_1059_315# 0.01136f
C48363 hold13/a_49_47# net160 0
C48364 _0528_/a_81_21# _0528_/a_384_47# 0.00138f
C48365 _0641_/a_113_47# net65 0
C48366 net36 _0851_/a_113_47# 0
C48367 _0568_/a_27_297# _0345_ 0.01474f
C48368 _0765_/a_79_21# _0381_ 0
C48369 _0586_/a_27_47# control0.add 0.19732f
C48370 _0310_ _0393_ 0
C48371 _0352_ _0103_ 0.0977f
C48372 hold101/a_285_47# _0431_ 0
C48373 net63 _0825_/a_68_297# 0
C48374 _0330_ net242 0.00866f
C48375 VPWR hold2/a_391_47# 0.18944f
C48376 net100 _0178_ 0
C48377 _0654_/a_297_47# _0345_ 0
C48378 _0820_/a_215_47# clknet_1_1__leaf__0465_ 0.00285f
C48379 _0962_/a_109_297# VPWR 0.00434f
C48380 _0328_ _0368_ 0.05262f
C48381 net193 _0540_/a_149_47# 0.01256f
C48382 hold46/a_49_47# net20 0.00233f
C48383 net36 net157 0.61058f
C48384 _0820_/a_79_21# _0088_ 0.04977f
C48385 _1058_/a_1059_315# _0181_ 0.00114f
C48386 _0210_ _0174_ 0
C48387 _0363_ _0735_/a_109_297# 0.01416f
C48388 _0312_ _0693_/a_68_297# 0
C48389 net33 control0.sh 0.10444f
C48390 _0369_ _0812_/a_297_297# 0.00204f
C48391 _1030_/a_27_47# clknet_1_1__leaf__0462_ 0.0041f
C48392 hold8/a_391_47# acc0.A\[26\] 0.07267f
C48393 comp0.B\[13\] _0138_ 0
C48394 _0337_ _0220_ 0.07157f
C48395 _0984_/a_193_47# _0350_ 0
C48396 _0284_ _0788_/a_68_297# 0
C48397 _0372_ _0748_/a_81_21# 0.11493f
C48398 net233 _0846_/a_245_297# 0
C48399 _0430_ _0443_ 0
C48400 net40 _0994_/a_1059_315# 0.00116f
C48401 hold33/a_285_47# comp0.B\[14\] 0
C48402 VPWR _1008_/a_27_47# 0.70441f
C48403 _0138_ _1046_/a_193_47# 0
C48404 clkbuf_1_0__f__0463_/a_110_47# _0546_/a_51_297# 0
C48405 _0855_/a_81_21# hold60/a_49_47# 0.00138f
C48406 hold16/a_391_47# VPWR 0.1933f
C48407 _0960_/a_27_47# control0.count\[0\] 0.10349f
C48408 hold38/a_391_47# _1062_/a_466_413# 0
C48409 net158 _1046_/a_27_47# 0.09866f
C48410 _0180_ _0528_/a_81_21# 0.00844f
C48411 hold100/a_285_47# _0448_ 0.00147f
C48412 clkbuf_1_1__f__0465_/a_110_47# _0516_/a_27_297# 0
C48413 _0857_/a_27_47# comp0.B\[0\] 0.0059f
C48414 control0.count\[2\] _0466_ 0.49687f
C48415 net187 net106 0
C48416 _0467_ _1062_/a_27_47# 0
C48417 net57 _0352_ 0
C48418 _1052_/a_381_47# _0186_ 0.00112f
C48419 hold5/a_49_47# clknet_1_1__leaf__0464_ 0
C48420 _0714_/a_51_297# acc0.A\[30\] 0.00206f
C48421 _0216_ _0347_ 0.02673f
C48422 net197 net113 0.05499f
C48423 net190 clknet_1_1__leaf__0462_ 0.17473f
C48424 net186 _1033_/a_381_47# 0
C48425 clknet_1_0__leaf__0458_ hold71/a_49_47# 0.02303f
C48426 _0244_ clknet_0__0461_ 0.00309f
C48427 _1058_/a_466_413# _0188_ 0
C48428 _1058_/a_27_47# _0155_ 0
C48429 _0343_ _0411_ 0.25478f
C48430 VPWR _0826_/a_219_297# 0.13115f
C48431 _0949_/a_59_75# _0468_ 0.19478f
C48432 _0972_/a_346_47# net17 0.00351f
C48433 _0405_ hold91/a_49_47# 0
C48434 _0305_ _1060_/a_1059_315# 0
C48435 _0307_ _0459_ 0.00658f
C48436 _0699_/a_68_297# _0699_/a_150_297# 0.00477f
C48437 _0612_/a_145_75# acc0.A\[18\] 0.00129f
C48438 _1036_/a_27_47# comp0.B\[5\] 0
C48439 _0183_ _1017_/a_27_47# 0
C48440 _0216_ _0104_ 0.24071f
C48441 _0467_ _0561_/a_51_297# 0
C48442 VPWR _0611_/a_68_297# 0.14925f
C48443 net180 _0137_ 0.40999f
C48444 _0533_/a_373_47# _0199_ 0.0022f
C48445 acc0.A\[1\] _0180_ 0.00881f
C48446 _1000_/a_193_47# _0459_ 0
C48447 comp0.B\[0\] _1062_/a_27_47# 0.00971f
C48448 pp[27] hold95/a_49_47# 0.0028f
C48449 net34 control0.count\[0\] 0
C48450 clkbuf_0__0458_/a_110_47# _0350_ 0.00181f
C48451 acc0.A\[1\] net218 0.02883f
C48452 _0183_ _1060_/a_975_413# 0
C48453 clknet_0__0458_ hold86/a_391_47# 0
C48454 clkbuf_1_0__f__0458_/a_110_47# net61 0
C48455 net66 net67 0
C48456 _0555_/a_240_47# net28 0.06002f
C48457 _0369_ clkbuf_1_0__f__0465_/a_110_47# 0.00104f
C48458 B[12] net195 0
C48459 control0.state\[1\] _1063_/a_27_47# 0.42431f
C48460 net16 input16/a_75_212# 0.1087f
C48461 clknet_1_1__leaf__0459_ net192 0
C48462 hold47/a_49_47# _0194_ 0
C48463 net105 _1014_/a_27_47# 0
C48464 VPWR hold84/a_49_47# 0.35541f
C48465 clknet_1_0__leaf__0462_ _1022_/a_1059_315# 0.01047f
C48466 _0123_ _1024_/a_1059_315# 0.00311f
C48467 _1005_/a_193_47# _1005_/a_634_159# 0.11897f
C48468 _1005_/a_27_47# _1005_/a_466_413# 0.27314f
C48469 _0978_/a_109_297# _0487_ 0
C48470 _0383_ hold3/a_285_47# 0
C48471 _0376_ hold94/a_391_47# 0.00858f
C48472 net236 control0.count\[2\] 0
C48473 net117 _1013_/a_193_47# 0
C48474 _0205_ net152 0
C48475 _0546_/a_149_47# _0139_ 0
C48476 VPWR net109 0.54114f
C48477 _0984_/a_891_413# _0849_/a_79_21# 0
C48478 _0472_ clknet_1_1__leaf__0457_ 0.01388f
C48479 clkbuf_1_1__f__0465_/a_110_47# _0399_ 0.04619f
C48480 hold45/a_391_47# VPWR 0.177f
C48481 net149 _0580_/a_373_47# 0.00247f
C48482 clknet_1_1__leaf__0459_ _0346_ 0.25184f
C48483 _0991_/a_27_47# net67 0
C48484 comp0.B\[14\] net20 0.02085f
C48485 _0991_/a_1059_315# net77 0
C48486 _0991_/a_466_413# _0089_ 0.02852f
C48487 _0210_ _0208_ 0.13193f
C48488 control0.state\[0\] _0460_ 0
C48489 _0467_ _0133_ 0
C48490 _0109_ _0345_ 0.00719f
C48491 _0355_ _0219_ 0.20554f
C48492 net78 net37 0.00177f
C48493 _0415_ _0993_/a_193_47# 0
C48494 _0297_ _0277_ 0.10198f
C48495 _0181_ net47 0.06672f
C48496 net53 hold90/a_285_47# 0.0234f
C48497 _0997_/a_381_47# clknet_1_1__leaf__0461_ 0
C48498 hold96/a_391_47# _0347_ 0
C48499 _0462_ _0743_/a_51_297# 0.00269f
C48500 _0260_ _0271_ 0
C48501 _0985_/a_193_47# _0261_ 0.01088f
C48502 _0985_/a_27_47# _0263_ 0
C48503 _0286_ _0808_/a_585_47# 0.00111f
C48504 _0286_ net79 0
C48505 net116 _0333_ 0
C48506 _0216_ _1029_/a_1017_47# 0
C48507 _0728_/a_59_75# _0355_ 0.0152f
C48508 _0603_/a_150_297# _0460_ 0
C48509 _0768_/a_27_47# _0393_ 0
C48510 clknet_1_1__leaf__0459_ _0992_/a_466_413# 0.0162f
C48511 _0730_/a_510_47# _0317_ 0
C48512 _0559_/a_51_297# net26 0.1012f
C48513 _0174_ _0542_/a_149_47# 0.01802f
C48514 VPWR _1065_/a_381_47# 0.07191f
C48515 _1038_/a_27_47# _1040_/a_27_47# 0
C48516 _1004_/a_975_413# acc0.A\[23\] 0
C48517 _1012_/a_27_47# hold92/a_49_47# 0
C48518 _0600_/a_337_297# _0600_/a_253_47# 0.00219f
C48519 _0946_/a_30_53# _0480_ 0
C48520 _0343_ clkload4/a_110_47# 0
C48521 _0247_ _0774_/a_68_297# 0.02608f
C48522 clkbuf_0__0462_/a_110_47# _0345_ 0
C48523 net123 _1037_/a_592_47# 0
C48524 _0133_ comp0.B\[0\] 0
C48525 _1038_/a_891_413# comp0.B\[4\] 0
C48526 _0995_/a_634_159# _0995_/a_1059_315# 0
C48527 _0995_/a_27_47# _0995_/a_381_47# 0.06222f
C48528 _0995_/a_193_47# _0995_/a_891_413# 0.19685f
C48529 _0529_/a_109_47# net170 0.00357f
C48530 _0412_ _0277_ 0
C48531 _0413_ _0300_ 0
C48532 _1021_/a_1017_47# _0183_ 0.00106f
C48533 _0138_ comp0.B\[9\] 0.05805f
C48534 net67 _0350_ 0
C48535 hold87/a_391_47# clknet_1_0__leaf__0458_ 0.00278f
C48536 hold59/a_285_47# _0612_/a_59_75# 0
C48537 _0216_ comp0.B\[1\] 0
C48538 net62 _0445_ 0.21462f
C48539 _1060_/a_975_413# acc0.A\[15\] 0
C48540 _0693_/a_150_297# _0219_ 0
C48541 net87 _0345_ 0
C48542 _0450_ _0445_ 0
C48543 VPWR pp[24] 0.21837f
C48544 net48 net109 0.05618f
C48545 hold9/a_285_47# _1027_/a_466_413# 0.00145f
C48546 VPWR _0819_/a_384_47# 0
C48547 _0234_ _0101_ 0
C48548 net32 _1042_/a_27_47# 0.4671f
C48549 net152 _1042_/a_193_47# 0.00137f
C48550 net76 acc0.A\[9\] 0
C48551 net53 _1007_/a_561_413# 0
C48552 _0467_ net107 0
C48553 _0227_ hold66/a_49_47# 0
C48554 _1070_/a_1059_315# _1069_/a_891_413# 0
C48555 _1070_/a_891_413# _1069_/a_1059_315# 0
C48556 hold45/a_391_47# input4/a_75_212# 0
C48557 _0292_ _0346_ 0.06518f
C48558 control0.reset _0493_/a_27_47# 0.00154f
C48559 control0.state\[1\] _1062_/a_1059_315# 0.00143f
C48560 _0243_ _0611_/a_150_297# 0
C48561 control0.state\[0\] _1062_/a_891_413# 0.04353f
C48562 net46 _0576_/a_373_47# 0
C48563 _0982_/a_27_47# _0183_ 0.02712f
C48564 _0982_/a_634_159# _0217_ 0
C48565 _1034_/a_27_47# _0473_ 0
C48566 _0461_ net104 0
C48567 hold74/a_49_47# _0115_ 0
C48568 net228 net229 0.07033f
C48569 hold25/a_391_47# input8/a_75_212# 0
C48570 _0490_ _0166_ 0
C48571 _1011_/a_1059_315# _1011_/a_891_413# 0.31086f
C48572 _1011_/a_193_47# _1011_/a_975_413# 0
C48573 _1011_/a_466_413# _1011_/a_381_47# 0.03733f
C48574 _0643_/a_253_47# net62 0.03762f
C48575 _0985_/a_193_47# _0509_/a_27_47# 0
C48576 _1016_/a_381_47# _0369_ 0
C48577 _0608_/a_109_297# _0347_ 0
C48578 net50 _1023_/a_1059_315# 0
C48579 _0935_/a_27_47# _0171_ 0.00966f
C48580 _0133_ _1034_/a_634_159# 0.00995f
C48581 _0171_ _1061_/a_193_47# 0
C48582 hold96/a_49_47# _0574_/a_27_297# 0.01494f
C48583 net97 _0350_ 0
C48584 hold29/a_49_47# acc0.A\[23\] 0.00104f
C48585 comp0.B\[1\] _1067_/a_27_47# 0
C48586 hold85/a_391_47# _0164_ 0
C48587 _0255_ _0193_ 0
C48588 clknet_0__0465_ _0986_/a_1017_47# 0
C48589 _0120_ net51 0.01297f
C48590 _0287_ _0992_/a_193_47# 0
C48591 _0289_ _0992_/a_634_159# 0
C48592 _0195_ net105 0.01876f
C48593 net45 _0997_/a_466_413# 0
C48594 _0535_/a_68_297# net22 0
C48595 net39 _0280_ 0
C48596 _0401_ _0089_ 0.00539f
C48597 _0234_ hold4/a_285_47# 0
C48598 _0992_/a_1059_315# hold81/a_391_47# 0
C48599 clkbuf_0_clk/a_110_47# _0163_ 0
C48600 _1021_/a_1059_315# hold73/a_391_47# 0.00615f
C48601 comp0.B\[0\] net107 0
C48602 _0216_ _1025_/a_27_47# 0
C48603 _1055_/a_634_159# VPWR 0.21278f
C48604 _0350_ _0986_/a_975_413# 0
C48605 _1020_/a_592_47# VPWR 0
C48606 _0266_ _0219_ 0
C48607 _1001_/a_193_47# acc0.A\[19\] 0.00193f
C48608 _1003_/a_193_47# VPWR 0.30713f
C48609 _0183_ net17 0
C48610 _0251_ _0828_/a_113_297# 0.02417f
C48611 _0982_/a_891_413# _0580_/a_109_297# 0
C48612 _0181_ _1063_/a_1059_315# 0
C48613 _0837_/a_266_297# _0218_ 0
C48614 clknet_0__0464_ _1049_/a_27_47# 0.00863f
C48615 _0827_/a_109_297# _0827_/a_27_47# 0
C48616 _0370_ clkbuf_0__0460_/a_110_47# 0.00108f
C48617 output54/a_27_47# clknet_1_1__leaf__0462_ 0.00111f
C48618 clk _0486_ 0.03386f
C48619 _0955_/a_304_297# _0474_ 0.00106f
C48620 comp0.B\[3\] comp0.B\[5\] 0.36942f
C48621 _0567_/a_109_297# _0219_ 0
C48622 _0216_ hold95/a_49_47# 0.00378f
C48623 _0195_ hold95/a_391_47# 0.00804f
C48624 hold44/a_285_47# _0127_ 0.07478f
C48625 _0298_ _0297_ 0.32653f
C48626 _0305_ _0294_ 0.38724f
C48627 _0150_ net13 0.01098f
C48628 _0794_/a_326_47# _0345_ 0.0013f
C48629 _0440_ _0186_ 0
C48630 _0733_/a_79_199# clknet_0__0462_ 0.01306f
C48631 net126 input7/a_75_212# 0
C48632 net65 _0435_ 0.02318f
C48633 _0966_/a_27_47# _0466_ 0
C48634 _1023_/a_27_47# _1023_/a_634_159# 0.14145f
C48635 A[14] _0411_ 0
C48636 clkbuf_1_0__f__0461_/a_110_47# _0616_/a_78_199# 0
C48637 _0183_ _0446_ 0
C48638 net167 _0479_ 0
C48639 net54 _0318_ 0.00411f
C48640 _0165_ _1067_/a_592_47# 0
C48641 net9 hold1/a_285_47# 0
C48642 _1042_/a_27_47# _1042_/a_1059_315# 0.04875f
C48643 _1042_/a_193_47# _1042_/a_466_413# 0.07478f
C48644 _0403_ _0402_ 0.00948f
C48645 _0181_ _1060_/a_1059_315# 0.07063f
C48646 _0583_/a_27_297# _0115_ 0
C48647 _1018_/a_27_47# net47 0
C48648 pp[17] hold61/a_49_47# 0
C48649 _0175_ _0563_/a_512_297# 0
C48650 _1037_/a_891_413# _0552_/a_68_297# 0.00123f
C48651 _1010_/a_561_413# _0347_ 0
C48652 _1010_/a_1059_315# _0352_ 0.00368f
C48653 _0815_/a_113_297# _0288_ 0
C48654 _0982_/a_27_47# acc0.A\[15\] 0
C48655 _1045_/a_1059_315# _0540_/a_51_297# 0
C48656 _0174_ net22 0.98679f
C48657 _0459_ _0507_/a_109_297# 0.00157f
C48658 _0531_/a_109_47# _0465_ 0
C48659 output43/a_27_47# net60 0
C48660 _1051_/a_561_413# clknet_1_1__leaf__0464_ 0
C48661 _0412_ _0298_ 0.24271f
C48662 _0413_ _0404_ 0.02606f
C48663 _0179_ _1050_/a_193_47# 0.021f
C48664 hold63/a_285_47# _0124_ 0.0336f
C48665 _0800_/a_245_297# _0219_ 0.00275f
C48666 pp[10] _0181_ 0
C48667 _0347_ _0841_/a_79_21# 0.11201f
C48668 _1036_/a_891_413# _1036_/a_975_413# 0.00851f
C48669 _1036_/a_381_47# _1036_/a_561_413# 0.00123f
C48670 _1039_/a_193_47# _0171_ 0
C48671 _0714_/a_512_297# _0339_ 0
C48672 _0145_ acc0.A\[15\] 0.02161f
C48673 hold69/a_49_47# net52 0.32259f
C48674 control0.sh _0563_/a_149_47# 0
C48675 pp[30] hold62/a_285_47# 0.00889f
C48676 net10 _1042_/a_27_47# 0.03382f
C48677 hold26/a_285_47# _0137_ 0
C48678 _0480_ _0487_ 0.01055f
C48679 net53 clknet_0__0462_ 0.00417f
C48680 _0526_/a_27_47# hold60/a_285_47# 0
C48681 _0767_/a_59_75# _0679_/a_150_297# 0
C48682 _0725_/a_303_47# _0353_ 0.00463f
C48683 VPWR _1040_/a_634_159# 0.18626f
C48684 _0129_ _0567_/a_27_297# 0.10909f
C48685 hold27/a_285_47# net7 0.04765f
C48686 clknet_1_0__leaf__0463_ _0174_ 0.73195f
C48687 _0966_/a_27_47# net236 0.01041f
C48688 _0176_ _0139_ 0.01765f
C48689 _0997_/a_193_47# _0793_/a_51_297# 0
C48690 net176 clknet_1_0__leaf__0460_ 0
C48691 _1041_/a_891_413# net18 0
C48692 _1041_/a_634_159# _0140_ 0
C48693 _1050_/a_891_413# _0194_ 0
C48694 _0227_ acc0.A\[22\] 0
C48695 acc0.A\[21\] _0183_ 0.47312f
C48696 _0333_ hold80/a_285_47# 0
C48697 net238 acc0.A\[15\] 0.02792f
C48698 _0410_ net42 0.02279f
C48699 pp[0] net29 0
C48700 _0238_ _0383_ 0
C48701 _1011_/a_193_47# _0334_ 0
C48702 hold13/a_391_47# clknet_0__0463_ 0
C48703 hold49/a_391_47# net19 0
C48704 acc0.A\[20\] net1 0
C48705 _0083_ _0465_ 0.003f
C48706 _0971_/a_81_21# _0160_ 0
C48707 _0163_ _1062_/a_381_47# 0
C48708 _0270_ _0444_ 0
C48709 clknet_1_0__leaf__0462_ _1024_/a_561_413# 0
C48710 _0467_ _1063_/a_561_413# 0
C48711 _1058_/a_381_47# net4 0.01447f
C48712 _1058_/a_1059_315# _0187_ 0.00273f
C48713 hold59/a_285_47# _0399_ 0.03771f
C48714 _0446_ acc0.A\[15\] 0.04545f
C48715 _1021_/a_381_47# _0181_ 0.0099f
C48716 _1032_/a_634_159# _1067_/a_27_47# 0
C48717 _0467_ _0959_/a_300_47# 0
C48718 net36 net172 0.11826f
C48719 VPWR _0471_ 0.91703f
C48720 clknet_1_0__leaf__0458_ _0264_ 0.04254f
C48721 hold30/a_391_47# _1022_/a_1059_315# 0
C48722 _0083_ acc0.A\[2\] 0.00178f
C48723 _1012_/a_891_413# net239 0.00147f
C48724 net233 _0448_ 0.2449f
C48725 _0456_ _0346_ 0.00508f
C48726 _0237_ _0103_ 0
C48727 net149 clknet_1_1__leaf__0457_ 0.67989f
C48728 _0112_ clkbuf_1_1__f__0457_/a_110_47# 0
C48729 _1054_/a_634_159# acc0.A\[7\] 0.00115f
C48730 _1054_/a_27_47# _0252_ 0
C48731 _0302_ net41 0.04505f
C48732 _0179_ _0518_/a_109_297# 0.00326f
C48733 _0195_ acc0.A\[28\] 0.93846f
C48734 _1054_/a_27_47# _0989_/a_381_47# 0
C48735 _0346_ _0655_/a_215_53# 0.00899f
C48736 net33 _0955_/a_32_297# 0.00652f
C48737 _0795_/a_299_297# net41 0.00271f
C48738 net197 hold8/a_285_47# 0
C48739 _0680_/a_80_21# _0246_ 0
C48740 _1057_/a_381_47# net189 0.12473f
C48741 VPWR _0688_/a_109_297# 0.00576f
C48742 _0626_/a_150_297# VPWR 0.00193f
C48743 B[13] net128 0.04005f
C48744 _0463_ _0498_/a_512_297# 0
C48745 net63 net148 0.00338f
C48746 _0675_/a_68_297# _0218_ 0.02694f
C48747 _0457_ _0565_/a_51_297# 0.00658f
C48748 _1053_/a_27_47# _1052_/a_466_413# 0
C48749 _1053_/a_193_47# _1052_/a_634_159# 0
C48750 _0579_/a_109_47# net211 0
C48751 _0550_/a_51_297# _1040_/a_193_47# 0
C48752 clknet_1_0__leaf__0460_ _0617_/a_68_297# 0.00318f
C48753 _0182_ _0495_/a_68_297# 0
C48754 _0195_ net209 0.19512f
C48755 _1059_/a_381_47# _0157_ 0.11485f
C48756 _0789_/a_315_47# _0299_ 0.00344f
C48757 _0251_ _0433_ 0
C48758 _0093_ _0995_/a_891_413# 0
C48759 _0181_ _0173_ 0
C48760 _0362_ _0319_ 0
C48761 _0754_/a_245_297# _0754_/a_240_47# 0
C48762 _0643_/a_103_199# _0271_ 0.00287f
C48763 _0643_/a_253_297# _0256_ 0
C48764 _0640_/a_109_53# _0433_ 0
C48765 _0421_ hold81/a_391_47# 0
C48766 _0183_ _0245_ 0.00106f
C48767 _0164_ _0160_ 0.00311f
C48768 _0196_ _0148_ 0.07242f
C48769 _0128_ _0345_ 0.00875f
C48770 clknet_1_0__leaf__0461_ _0242_ 0.16165f
C48771 _0959_/a_300_47# comp0.B\[0\] 0
C48772 input24/a_75_212# _0175_ 0
C48773 _0179_ _0145_ 0.00801f
C48774 _0673_/a_253_297# _0345_ 0
C48775 net44 clknet_1_1__leaf__0462_ 0.29688f
C48776 _0476_ net28 0
C48777 _1055_/a_891_413# clknet_1_1__leaf__0465_ 0.0016f
C48778 _0672_/a_297_297# _0345_ 0
C48779 hold11/a_285_47# clknet_1_0__leaf__0465_ 0.02859f
C48780 _0710_/a_381_47# _0342_ 0.00786f
C48781 _0341_ _0340_ 0.34474f
C48782 _0779_/a_215_47# _0352_ 0
C48783 clkbuf_0_clk/a_110_47# _1068_/a_27_47# 0.00398f
C48784 control0.reset clkbuf_1_1__f_clk/a_110_47# 0.00373f
C48785 _0673_/a_253_47# _0295_ 0.031f
C48786 clknet_1_0__leaf__0458_ net170 0
C48787 _0555_/a_245_297# _0210_ 0.00111f
C48788 _0555_/a_512_297# net160 0
C48789 _0663_/a_207_413# _0288_ 0.00399f
C48790 net14 hold83/a_391_47# 0
C48791 _1038_/a_27_47# net171 0
C48792 _0304_ _0672_/a_215_47# 0.00299f
C48793 _0328_ clknet_0__0460_ 0
C48794 _1051_/a_634_159# _0524_/a_27_297# 0
C48795 _1051_/a_193_47# _0524_/a_109_297# 0
C48796 clknet_1_0__leaf__0463_ _0208_ 0
C48797 pp[16] net40 0
C48798 _0454_ _0849_/a_215_47# 0
C48799 _0992_/a_1059_315# _0281_ 0.00176f
C48800 hold23/a_391_47# _0260_ 0
C48801 _1046_/a_1059_315# _0142_ 0.00167f
C48802 _1053_/a_634_159# net12 0.00206f
C48803 _0389_ hold76/a_49_47# 0
C48804 _0734_/a_47_47# clknet_1_1__leaf__0460_ 0.00382f
C48805 _0530_/a_299_297# _0186_ 0.00688f
C48806 net81 pp[14] 0
C48807 VPWR _0994_/a_634_159# 0.19387f
C48808 _0974_/a_448_47# _1068_/a_634_159# 0
C48809 _0852_/a_35_297# _0269_ 0
C48810 net58 _0433_ 0
C48811 clknet_1_0__leaf__0462_ _0315_ 0.29304f
C48812 _0195_ hold72/a_49_47# 0
C48813 _0229_ net150 0.00172f
C48814 clkbuf_0__0465_/a_110_47# _0841_/a_79_21# 0
C48815 _0343_ _0988_/a_1059_315# 0.00462f
C48816 _0179_ _0446_ 0.01546f
C48817 _0461_ _1015_/a_634_159# 0
C48818 _1038_/a_27_47# net24 0
C48819 _0179_ input2/a_75_212# 0.06576f
C48820 _1010_/a_27_47# _0350_ 0.09301f
C48821 _0399_ _0830_/a_79_21# 0.11953f
C48822 pp[27] _1011_/a_27_47# 0
C48823 _0646_/a_47_47# _0299_ 0
C48824 _0216_ _0106_ 0
C48825 _1034_/a_891_413# _0959_/a_80_21# 0
C48826 _0576_/a_109_297# net176 0.01209f
C48827 _0338_ hold62/a_391_47# 0
C48828 _0339_ hold62/a_285_47# 0.03548f
C48829 _1039_/a_27_47# control0.sh 0
C48830 _0697_/a_80_21# _0697_/a_472_297# 0.01636f
C48831 _0294_ _0181_ 0.68515f
C48832 _0785_/a_384_47# _0428_ 0
C48833 _0341_ _1013_/a_381_47# 0
C48834 hold16/a_49_47# _0128_ 0
C48835 _0179_ net194 0
C48836 net157 _1061_/a_27_47# 0.0059f
C48837 _0331_ _0697_/a_80_21# 0
C48838 _0151_ _1052_/a_27_47# 0.00107f
C48839 hold63/a_49_47# _1026_/a_27_47# 0.00166f
C48840 _0990_/a_27_47# clknet_1_1__leaf__0458_ 0.01039f
C48841 net56 _0331_ 0.0365f
C48842 _0995_/a_27_47# _0219_ 0.00629f
C48843 VPWR hold93/a_391_47# 0.18716f
C48844 comp0.B\[4\] _0955_/a_220_297# 0.01299f
C48845 _0521_/a_299_297# _0179_ 0.05006f
C48846 _0174_ _0544_/a_245_297# 0.0022f
C48847 acc0.A\[0\] clkbuf_0__0457_/a_110_47# 0
C48848 _0820_/a_297_297# _0399_ 0.00681f
C48849 _0670_/a_79_21# clkbuf_0__0459_/a_110_47# 0
C48850 _1009_/a_193_47# _0350_ 0.00545f
C48851 _0217_ net103 0
C48852 clknet_1_0__leaf__0462_ net150 0.05354f
C48853 _1031_/a_634_159# _1031_/a_1059_315# 0
C48854 _1031_/a_27_47# _1031_/a_381_47# 0.06222f
C48855 _1031_/a_193_47# _1031_/a_891_413# 0.19497f
C48856 net41 net6 0.04204f
C48857 _0247_ hold72/a_391_47# 0
C48858 clkbuf_1_0__f__0462_/a_110_47# _0250_ 0
C48859 B[8] net152 0
C48860 _0996_/a_466_413# _0346_ 0
C48861 _0804_/a_215_47# _0403_ 0
C48862 net23 net201 0
C48863 _1000_/a_634_159# _0218_ 0
C48864 output42/a_27_47# _0995_/a_193_47# 0
C48865 _0722_/a_79_21# _0722_/a_297_297# 0.01735f
C48866 _1005_/a_1059_315# _1005_/a_1017_47# 0
C48867 _1005_/a_193_47# net91 0.009f
C48868 _1005_/a_27_47# _0103_ 0.09891f
C48869 _0220_ _0333_ 0
C48870 _0244_ _0616_/a_215_47# 0.00136f
C48871 hold66/a_391_47# net49 0.00141f
C48872 control0.state\[0\] _0470_ 0
C48873 hold55/a_285_47# _0183_ 0
C48874 VPWR _0729_/a_150_297# 0.00223f
C48875 _0984_/a_381_47# _0082_ 0.13126f
C48876 net61 _0183_ 0
C48877 _1066_/a_27_47# _1062_/a_381_47# 0
C48878 _1066_/a_381_47# _1062_/a_27_47# 0
C48879 _1060_/a_193_47# acc0.A\[13\] 0
C48880 net15 input15/a_75_212# 0.11027f
C48881 _1013_/a_634_159# _1013_/a_592_47# 0
C48882 _0976_/a_76_199# _1069_/a_27_47# 0
C48883 net1 _1062_/a_27_47# 0
C48884 VPWR _0853_/a_150_297# 0.00123f
C48885 _1002_/a_27_47# _1002_/a_561_413# 0.0027f
C48886 _1002_/a_634_159# _1002_/a_891_413# 0.03684f
C48887 _1002_/a_193_47# _1002_/a_381_47# 0.09503f
C48888 _0836_/a_68_297# acc0.A\[6\] 0
C48889 hold68/a_285_47# _0576_/a_27_297# 0
C48890 hold68/a_49_47# _0576_/a_109_297# 0
C48891 comp0.B\[0\] _0208_ 0.09051f
C48892 comp0.B\[13\] net22 0
C48893 _0985_/a_27_47# hold28/a_391_47# 0
C48894 _0985_/a_193_47# hold28/a_285_47# 0
C48895 clknet_1_0__leaf__0465_ _0524_/a_27_297# 0.01258f
C48896 _0984_/a_466_413# clknet_1_0__leaf__0458_ 0.00343f
C48897 _0309_ _0393_ 0
C48898 net63 _0837_/a_81_21# 0.00145f
C48899 _1027_/a_891_413# _0347_ 0
C48900 net86 clknet_1_0__leaf__0461_ 0
C48901 net212 acc0.A\[6\] 0.03118f
C48902 net22 _1046_/a_193_47# 0
C48903 _0310_ _0773_/a_35_297# 0
C48904 clknet_1_1__leaf__0459_ _0997_/a_1017_47# 0
C48905 _0583_/a_27_297# net146 0
C48906 _0243_ _0461_ 0.03317f
C48907 pp[30] _0350_ 0
C48908 VPWR _0989_/a_561_413# 0.0032f
C48909 _1039_/a_27_47# net157 0
C48910 _0248_ _0246_ 0.00476f
C48911 _0183_ _0165_ 0
C48912 VPWR _0997_/a_466_413# 0.26883f
C48913 VPWR control0.reset 1.42631f
C48914 _1059_/a_193_47# _0369_ 0.02864f
C48915 _0217_ _1019_/a_1059_315# 0
C48916 _0183_ _1019_/a_634_159# 0.02155f
C48917 VPWR _0992_/a_561_413# 0.00319f
C48918 _1055_/a_27_47# acc0.A\[6\] 0
C48919 net104 _0582_/a_27_297# 0
C48920 hold35/a_285_47# net181 0
C48921 control0.state\[1\] _0958_/a_197_47# 0
C48922 control0.state\[0\] _0958_/a_303_47# 0
C48923 _1035_/a_634_159# _0175_ 0.00791f
C48924 hold20/a_285_47# _0486_ 0
C48925 VPWR _1061_/a_891_413# 0.2012f
C48926 _1011_/a_193_47# _0724_/a_113_297# 0
C48927 clknet_1_0__leaf__0463_ _1046_/a_193_47# 0
C48928 _0100_ _0382_ 0
C48929 _0375_ _0460_ 0
C48930 _0201_ _0537_/a_150_297# 0
C48931 _0350_ _0771_/a_215_297# 0
C48932 VPWR _0977_/a_75_212# 0.21833f
C48933 _1034_/a_891_413# _0173_ 0.00787f
C48934 _1034_/a_381_47# _0213_ 0
C48935 _1034_/a_27_47# _0132_ 0
C48936 acc0.A\[12\] _0512_/a_109_47# 0
C48937 hold87/a_49_47# _0081_ 0
C48938 hold9/a_285_47# net156 0.0127f
C48939 _1018_/a_592_47# _0459_ 0
C48940 net61 acc0.A\[15\] 0.00443f
C48941 _0975_/a_59_75# _0484_ 0
C48942 control0.state\[2\] _0970_/a_27_297# 0.00201f
C48943 control0.count\[1\] _1069_/a_466_413# 0.00779f
C48944 _1070_/a_466_413# control0.count\[0\] 0.00176f
C48945 _0327_ _0725_/a_209_47# 0
C48946 VPWR _1069_/a_975_413# 0.00459f
C48947 net34 _0160_ 0
C48948 net53 hold53/a_49_47# 0.0164f
C48949 output64/a_27_47# net178 0
C48950 net68 _0217_ 0
C48951 comp0.B\[2\] _0957_/a_32_297# 0
C48952 net185 _1066_/a_27_47# 0
C48953 B[13] input18/a_75_212# 0
C48954 input21/a_75_212# B[10] 0.00243f
C48955 _0399_ _0219_ 0.08181f
C48956 hold18/a_49_47# _0264_ 0
C48957 _1018_/a_27_47# _0294_ 0
C48958 _0312_ _0743_/a_51_297# 0
C48959 _1056_/a_891_413# _1058_/a_27_47# 0
C48960 _1056_/a_27_47# _1058_/a_891_413# 0
C48961 _0762_/a_79_21# _1005_/a_1059_315# 0
C48962 _1011_/a_466_413# net57 0
C48963 _0216_ _1011_/a_27_47# 0.00373f
C48964 _0985_/a_561_413# _0186_ 0.00137f
C48965 _0525_/a_81_21# _0525_/a_299_297# 0.08213f
C48966 _0399_ _0669_/a_111_297# 0
C48967 _1055_/a_1059_315# A[9] 0
C48968 _0195_ clknet_0__0461_ 0
C48969 comp0.B\[2\] net23 0
C48970 _0180_ _0198_ 0.06366f
C48971 _0179_ _0987_/a_193_47# 0
C48972 hold47/a_49_47# _1049_/a_193_47# 0
C48973 hold47/a_285_47# _1049_/a_27_47# 0
C48974 _1006_/a_634_159# _1006_/a_975_413# 0
C48975 _1006_/a_466_413# _1006_/a_561_413# 0.00772f
C48976 clkbuf_1_1__f__0462_/a_110_47# clknet_0__0462_ 0.31132f
C48977 _0201_ VPWR 0.23696f
C48978 _0286_ _0301_ 0
C48979 _0198_ net218 0.08302f
C48980 _0993_/a_27_47# net246 0.00712f
C48981 acc0.A\[1\] _1014_/a_1059_315# 0
C48982 _0476_ _0972_/a_250_297# 0
C48983 _0731_/a_81_21# acc0.A\[27\] 0
C48984 _0331_ _0345_ 0
C48985 _0116_ _0580_/a_27_297# 0
C48986 _0221_ _0725_/a_209_297# 0.08223f
C48987 _1052_/a_466_413# A[5] 0
C48988 _0984_/a_27_47# _0984_/a_561_413# 0.0027f
C48989 _0984_/a_634_159# _0984_/a_891_413# 0.03684f
C48990 _0984_/a_193_47# _0984_/a_381_47# 0.09503f
C48991 _1031_/a_27_47# _0219_ 0
C48992 net187 net220 0.00349f
C48993 _0808_/a_81_21# _0417_ 0.08333f
C48994 net141 VPWR 0.42343f
C48995 _0677_/a_47_47# _0218_ 0
C48996 clkload0/a_27_47# _0466_ 0.00237f
C48997 _0550_/a_51_297# _0207_ 0.10938f
C48998 acc0.A\[14\] net43 0
C48999 hold66/a_49_47# _0352_ 0
C49000 comp0.B\[3\] hold84/a_49_47# 0
C49001 hold69/a_391_47# _0346_ 0.05372f
C49002 net44 hold92/a_49_47# 0
C49003 net35 _1068_/a_1017_47# 0
C49004 _1039_/a_891_413# VPWR 0.18119f
C49005 _0343_ hold19/a_285_47# 0.02249f
C49006 _0664_/a_79_21# hold81/a_49_47# 0.00136f
C49007 _0712_/a_297_297# _1031_/a_891_413# 0
C49008 _0986_/a_634_159# _0986_/a_975_413# 0
C49009 _0986_/a_466_413# _0986_/a_561_413# 0.00772f
C49010 clknet_0__0458_ _0268_ 0.39491f
C49011 clkbuf_1_0__f__0458_/a_110_47# _0269_ 0.00193f
C49012 _0856_/a_297_297# _0264_ 0
C49013 _1023_/a_381_47# _1023_/a_561_413# 0.00123f
C49014 _1023_/a_27_47# net109 0.23032f
C49015 _1023_/a_891_413# _1023_/a_975_413# 0.00851f
C49016 _0990_/a_193_47# net47 0.0285f
C49017 pp[0] comp0.B\[6\] 0.00193f
C49018 hold49/a_285_47# net198 0
C49019 net1 net107 0
C49020 net22 comp0.B\[9\] 0.0087f
C49021 _1042_/a_891_413# _1042_/a_1017_47# 0.00617f
C49022 hold19/a_49_47# acc0.A\[17\] 0
C49023 _0114_ _0115_ 0
C49024 _0314_ _0216_ 0
C49025 net36 hold59/a_391_47# 0.00209f
C49026 net117 net59 0.0018f
C49027 pp[22] pp[24] 0.09033f
C49028 pp[15] _0297_ 0.00119f
C49029 clknet_1_1__leaf__0464_ _1044_/a_975_413# 0
C49030 hold9/a_285_47# acc0.A\[26\] 0.00168f
C49031 output36/a_27_47# net36 0.19073f
C49032 _1045_/a_891_413# net20 0.02068f
C49033 _1045_/a_634_159# _0142_ 0
C49034 _1037_/a_27_47# control0.sh 0.00177f
C49035 net168 _0433_ 0
C49036 net61 _0179_ 0.03708f
C49037 _0855_/a_81_21# clknet_1_0__leaf__0461_ 0.00237f
C49038 _0718_/a_47_47# hold62/a_285_47# 0.01036f
C49039 _0757_/a_68_297# _0756_/a_47_47# 0.007f
C49040 net141 output62/a_27_47# 0
C49041 comp0.B\[3\] _1065_/a_381_47# 0
C49042 _0111_ _0339_ 0.00613f
C49043 clknet_1_0__leaf__0464_ _0531_/a_109_297# 0
C49044 hold16/a_49_47# _1031_/a_1059_315# 0
C49045 hold16/a_391_47# _1031_/a_634_159# 0
C49046 hold16/a_285_47# _1031_/a_466_413# 0.0041f
C49047 _0498_/a_240_47# _0176_ 0
C49048 _0226_ net213 0.00938f
C49049 _0984_/a_381_47# net145 0
C49050 clknet_1_0__leaf__0463_ comp0.B\[9\] 0.01634f
C49051 _0710_/a_109_47# _0216_ 0.00442f
C49052 _0578_/a_27_297# _1067_/a_27_47# 0
C49053 hold22/a_49_47# net65 0
C49054 _1012_/a_27_47# _0218_ 0
C49055 hold77/a_285_47# _0219_ 0.00536f
C49056 _0752_/a_384_47# net51 0
C49057 pp[29] _1011_/a_381_47# 0
C49058 _0578_/a_109_297# _0369_ 0
C49059 _0387_ _0310_ 0.48147f
C49060 _1057_/a_27_47# _0156_ 0
C49061 _1038_/a_27_47# _1037_/a_466_413# 0
C49062 _1038_/a_466_413# _1037_/a_27_47# 0
C49063 _0732_/a_80_21# net51 0
C49064 _1056_/a_193_47# net47 0
C49065 output42/a_27_47# _0093_ 0.01427f
C49066 _0981_/a_109_297# _0488_ 0.0015f
C49067 _0981_/a_27_297# _0466_ 0.19389f
C49068 _0324_ _0319_ 0.58786f
C49069 net101 _1020_/a_634_159# 0
C49070 _0997_/a_1059_315# _0407_ 0
C49071 _0732_/a_209_297# _0105_ 0
C49072 _0855_/a_299_297# net47 0
C49073 hold46/a_285_47# hold6/a_49_47# 0
C49074 _0605_/a_109_297# clknet_1_0__leaf__0460_ 0
C49075 net194 _0141_ 0
C49076 clknet_1_0__leaf__0458_ _0856_/a_79_21# 0
C49077 _0195_ _0702_/a_113_47# 0
C49078 _0790_/a_285_297# net41 0
C49079 _0777_/a_377_297# _0394_ 0.00281f
C49080 _1002_/a_891_413# net220 0
C49081 _1002_/a_1059_315# _0385_ 0
C49082 _1054_/a_381_47# net11 0.01183f
C49083 hold30/a_285_47# _0217_ 0.06454f
C49084 hold30/a_49_47# acc0.A\[22\] 0.00502f
C49085 hold28/a_391_47# _0197_ 0
C49086 _0216_ _0180_ 0
C49087 _0259_ _0292_ 0.12106f
C49088 _0571_/a_27_297# acc0.A\[27\] 0.13564f
C49089 net53 _0687_/a_59_75# 0.00163f
C49090 _0532_/a_81_21# _0532_/a_299_297# 0.08213f
C49091 clkbuf_1_0__f__0460_/a_110_47# net51 0.00613f
C49092 acc0.A\[25\] _0364_ 0
C49093 _1033_/a_193_47# _0565_/a_51_297# 0
C49094 _1057_/a_193_47# _0992_/a_1059_315# 0
C49095 _0743_/a_245_297# _0219_ 0
C49096 _0218_ _0242_ 0.50665f
C49097 _0180_ clknet_1_1__leaf__0464_ 0.0402f
C49098 _0999_/a_592_47# _0218_ 0.00188f
C49099 _0641_/a_113_47# _0253_ 0
C49100 control0.count\[2\] _1069_/a_1059_315# 0
C49101 net140 acc0.A\[7\] 0
C49102 _0627_/a_215_53# clkbuf_0__0465_/a_110_47# 0.00687f
C49103 _0216_ _1013_/a_193_47# 0
C49104 _0195_ _1013_/a_466_413# 0.01804f
C49105 _0636_/a_59_75# _0261_ 0.00182f
C49106 _0636_/a_145_75# _0262_ 0
C49107 net33 _0474_ 0
C49108 _0250_ net51 0.09209f
C49109 _0238_ _0749_/a_81_21# 0
C49110 _0728_/a_145_75# _0353_ 0
C49111 _0455_ _0264_ 0
C49112 clkbuf_1_1__f__0463_/a_110_47# net119 0.01001f
C49113 clknet_0__0457_ clknet_1_1__leaf__0463_ 0
C49114 input26/a_75_212# net26 0.10856f
C49115 net188 A[10] 0.00149f
C49116 _0548_/a_149_47# net152 0
C49117 _0463_ _0159_ 0.0022f
C49118 net144 _0653_/a_113_47# 0
C49119 _0107_ _0219_ 0.11306f
C49120 _1000_/a_891_413# net223 0
C49121 VPWR _1035_/a_975_413# 0.00513f
C49122 _0172_ _1040_/a_193_47# 0.03283f
C49123 net180 _1040_/a_466_413# 0
C49124 acc0.A\[22\] _0352_ 0
C49125 _0217_ _0102_ 0
C49126 net236 _0981_/a_27_297# 0.01286f
C49127 _1058_/a_193_47# VPWR 0.30142f
C49128 _0788_/a_68_297# _0347_ 0.01934f
C49129 _0299_ _0219_ 0
C49130 _0345_ _0377_ 0.09358f
C49131 _0814_/a_27_47# _0814_/a_181_47# 0.00401f
C49132 _0191_ net75 0
C49133 _0305_ _0371_ 0
C49134 _0447_ _0350_ 0.13425f
C49135 _1056_/a_891_413# pp[8] 0
C49136 _1055_/a_1059_315# _0516_/a_27_297# 0
C49137 acc0.A\[27\] _0737_/a_117_297# 0
C49138 _1064_/a_634_159# _1064_/a_381_47# 0
C49139 _0234_ _0750_/a_27_47# 0
C49140 _1015_/a_193_47# net23 0
C49141 _0294_ clknet_1_1__leaf__0461_ 0.00745f
C49142 VPWR _0869_/a_27_47# 0.19708f
C49143 _1000_/a_1059_315# _0581_/a_27_297# 0
C49144 clknet_1_1__leaf_clk _1063_/a_27_47# 0.22583f
C49145 _0707_/a_75_199# _0334_ 0.24484f
C49146 _0442_ _0987_/a_27_47# 0
C49147 hold65/a_49_47# pp[3] 0
C49148 _1038_/a_1017_47# _0207_ 0
C49149 net80 net6 0
C49150 _0672_/a_79_21# _0301_ 0.0838f
C49151 _0244_ _0771_/a_215_297# 0
C49152 _0386_ _0771_/a_27_413# 0
C49153 _0279_ _0716_/a_27_47# 0
C49154 net137 _0524_/a_27_297# 0.00114f
C49155 net55 _0701_/a_80_21# 0
C49156 _0983_/a_891_413# _0582_/a_27_297# 0
C49157 _0343_ _1017_/a_634_159# 0.00194f
C49158 _1002_/a_27_47# _0369_ 0.00473f
C49159 _0081_ _0082_ 0.00192f
C49160 _0521_/a_81_21# hold83/a_285_47# 0
C49161 acc0.A\[11\] _0186_ 0.18562f
C49162 B[1] net29 0
C49163 _0845_/a_109_47# _0449_ 0.04919f
C49164 net139 net12 0.0471f
C49165 comp0.B\[14\] hold6/a_285_47# 0
C49166 hold41/a_49_47# _0512_/a_27_297# 0.00173f
C49167 _0217_ _0774_/a_68_297# 0.0011f
C49168 _0343_ _1060_/a_1017_47# 0
C49169 _0974_/a_544_297# _0166_ 0
C49170 control0.state\[1\] _0484_ 0
C49171 _0736_/a_56_297# _0318_ 0.00168f
C49172 control0.state\[0\] _0485_ 0.75449f
C49173 _0674_/a_113_47# _0347_ 0
C49174 clknet_1_0__leaf__0458_ _0454_ 0.00786f
C49175 _1017_/a_193_47# acc0.A\[17\] 0
C49176 net11 _0522_/a_27_297# 0
C49177 _0136_ _0552_/a_68_297# 0.0012f
C49178 hold25/a_391_47# net8 0.06735f
C49179 _1008_/a_27_47# _0345_ 0
C49180 _0737_/a_285_47# _0321_ 0
C49181 _0737_/a_117_297# _0364_ 0
C49182 clkbuf_1_1__f__0465_/a_110_47# _0346_ 0
C49183 net58 _0266_ 0
C49184 hold16/a_391_47# _0345_ 0
C49185 clknet_1_1__leaf__0464_ _1042_/a_466_413# 0
C49186 _0222_ _0103_ 0.47782f
C49187 hold2/a_49_47# hold2/a_391_47# 0.00188f
C49188 _0763_/a_109_47# net92 0
C49189 _0697_/a_300_47# _0329_ 0
C49190 _0287_ _0420_ 0.23237f
C49191 _0768_/a_27_47# _0387_ 0.04339f
C49192 hold74/a_285_47# _1016_/a_27_47# 0
C49193 hold74/a_49_47# _1016_/a_193_47# 0
C49194 B[13] comp0.B\[11\] 0.08803f
C49195 _0217_ _0574_/a_109_47# 0.00349f
C49196 _0989_/a_891_413# acc0.A\[6\] 0
C49197 clkbuf_1_1__f_clk/a_110_47# _1063_/a_193_47# 0.00247f
C49198 _0800_/a_149_47# _0997_/a_466_413# 0
C49199 hold36/a_285_47# net183 0.00851f
C49200 _0830_/a_215_47# _0830_/a_510_47# 0.00529f
C49201 _0787_/a_80_21# VPWR 0.15758f
C49202 _0179_ _0812_/a_215_47# 0.0097f
C49203 _0681_/a_113_47# _0324_ 0
C49204 _0429_ _0829_/a_109_297# 0.00158f
C49205 _0180_ net247 0.02595f
C49206 clknet_1_0__leaf__0465_ _1052_/a_466_413# 0.00186f
C49207 _0179_ _0514_/a_27_297# 0.01915f
C49208 _0643_/a_253_297# clknet_0__0465_ 0
C49209 _1038_/a_27_47# _0553_/a_51_297# 0
C49210 _1037_/a_891_413# VPWR 0.19129f
C49211 net61 _0441_ 0
C49212 net247 net218 0.03064f
C49213 clkbuf_1_1__f_clk/a_110_47# _0460_ 0.0079f
C49214 _0570_/a_27_297# _1028_/a_27_47# 0
C49215 net9 _1047_/a_193_47# 0
C49216 net224 _0318_ 0
C49217 VPWR _0633_/a_109_297# 0.00555f
C49218 _0255_ hold1/a_285_47# 0.06304f
C49219 _0080_ clknet_1_1__leaf__0457_ 0
C49220 _0954_/a_32_297# _0176_ 0
C49221 acc0.A\[0\] _0350_ 0
C49222 _0733_/a_448_47# _0324_ 0
C49223 _1041_/a_975_413# VPWR 0.00463f
C49224 _0489_ _0976_/a_76_199# 0.07992f
C49225 _0316_ _0319_ 0.05011f
C49226 _0098_ _0294_ 0.03454f
C49227 net86 _0218_ 0.25161f
C49228 _0722_/a_215_47# _0110_ 0.0044f
C49229 pp[15] _0995_/a_561_413# 0
C49230 _0800_/a_51_297# _0668_/a_79_21# 0
C49231 _0226_ _0603_/a_68_297# 0.00304f
C49232 net17 _0565_/a_240_47# 0.05893f
C49233 _0260_ _0529_/a_373_47# 0
C49234 hold24/a_285_47# net8 0.05331f
C49235 _0438_ _0831_/a_285_47# 0.00206f
C49236 _0226_ hold73/a_391_47# 0
C49237 control0.sh _1062_/a_27_47# 0
C49238 clknet_1_1__leaf_clk _1062_/a_1059_315# 0.00123f
C49239 _1018_/a_193_47# _0581_/a_27_297# 0.01145f
C49240 _1018_/a_27_47# _0581_/a_109_297# 0
C49241 net162 hold62/a_49_47# 0
C49242 VPWR _0831_/a_35_297# 0.17662f
C49243 _0488_ _1069_/a_27_47# 0
C49244 _0347_ _0319_ 0
C49245 _1021_/a_634_159# clknet_1_1__leaf_clk 0
C49246 hold16/a_49_47# hold16/a_391_47# 0.00188f
C49247 _0457_ clkbuf_1_1__f_clk/a_110_47# 0
C49248 hold91/a_49_47# hold91/a_285_47# 0.22264f
C49249 _1020_/a_27_47# _1020_/a_891_413# 0.03224f
C49250 _1020_/a_193_47# _1020_/a_1059_315# 0.03405f
C49251 _1020_/a_634_159# _1020_/a_466_413# 0.23992f
C49252 _1002_/a_1059_315# _0100_ 0.07031f
C49253 _1002_/a_891_413# net88 0
C49254 acc0.A\[23\] _0754_/a_149_47# 0
C49255 _0792_/a_209_297# _0406_ 0.04372f
C49256 _0408_ _0790_/a_35_297# 0.00386f
C49257 _0182_ _0844_/a_297_47# 0
C49258 hold12/a_49_47# hold12/a_285_47# 0.22264f
C49259 clknet_1_0__leaf__0465_ _0194_ 0.03999f
C49260 _0179_ net132 0.02125f
C49261 _0352_ _0379_ 0.04779f
C49262 net29 _1040_/a_1017_47# 0
C49263 _1016_/a_193_47# _0583_/a_27_297# 0
C49264 _0107_ _0746_/a_81_21# 0
C49265 _0598_/a_297_47# _0752_/a_27_413# 0
C49266 _0820_/a_79_21# net214 0.05342f
C49267 net216 _0368_ 0
C49268 _0372_ _0352_ 0.04634f
C49269 _0983_/a_466_413# net47 0.03397f
C49270 _0340_ acc0.A\[30\] 0.04429f
C49271 _1016_/a_634_159# net43 0
C49272 _0984_/a_193_47# _0081_ 0
C49273 _0984_/a_1059_315# _0454_ 0
C49274 _1028_/a_27_47# hold50/a_49_47# 0.0019f
C49275 hold35/a_285_47# net179 0
C49276 hold35/a_391_47# net141 0
C49277 _1058_/a_1059_315# clknet_1_1__leaf__0465_ 0
C49278 control0.sh _0561_/a_51_297# 0
C49279 _0259_ _0785_/a_299_297# 0.0592f
C49280 _0183_ net105 0
C49281 _0346_ _0673_/a_253_47# 0
C49282 _0180_ _1048_/a_466_413# 0.01012f
C49283 _0182_ _1048_/a_1059_315# 0.00171f
C49284 net175 _0186_ 0.00465f
C49285 _1049_/a_891_413# _0145_ 0
C49286 _1001_/a_891_413# net46 0.03939f
C49287 net14 net9 0
C49288 _0346_ _0672_/a_510_47# 0.00213f
C49289 net104 _0115_ 0.00186f
C49290 net1 _0208_ 0.05669f
C49291 _1041_/a_466_413# _0550_/a_240_47# 0
C49292 _0457_ _0584_/a_109_297# 0
C49293 _0172_ _0214_ 0
C49294 _0432_ _0825_/a_68_297# 0.10503f
C49295 _0272_ clkbuf_1_1__f__0458_/a_110_47# 0
C49296 _0217_ _1025_/a_1059_315# 0
C49297 net121 _0175_ 0.07678f
C49298 _0337_ hold95/a_49_47# 0
C49299 _1003_/a_466_413# _0466_ 0
C49300 _0430_ clknet_0__0458_ 0.05092f
C49301 _0566_/a_27_47# clknet_1_0__leaf__0461_ 0
C49302 pp[28] _1011_/a_1017_47# 0
C49303 _1039_/a_193_47# _0494_/a_27_47# 0
C49304 _0230_ _0368_ 0
C49305 clkbuf_1_1__f_clk/a_110_47# _1062_/a_891_413# 0
C49306 clkbuf_1_0__f__0465_/a_110_47# net75 0
C49307 clknet_1_0__leaf__0458_ _0846_/a_51_297# 0
C49308 _0664_/a_382_297# VPWR 0.00508f
C49309 _0113_ control0.reset 0
C49310 hold94/a_49_47# _0754_/a_51_297# 0
C49311 _0545_/a_68_297# _1040_/a_1059_315# 0
C49312 _0352_ hold40/a_49_47# 0.04524f
C49313 _0837_/a_266_47# _1051_/a_1059_315# 0
C49314 comp0.B\[2\] _0213_ 0.19636f
C49315 _0163_ _0487_ 0.11099f
C49316 _1036_/a_381_47# input24/a_75_212# 0
C49317 _0856_/a_79_21# hold18/a_49_47# 0
C49318 _0133_ control0.sh 0.02373f
C49319 _0230_ _0618_/a_215_47# 0
C49320 clknet_0__0458_ acc0.A\[5\] 0
C49321 _0176_ net173 0.19708f
C49322 _1000_/a_561_413# _0393_ 0
C49323 net86 _0775_/a_215_47# 0
C49324 _0580_/a_109_297# _0350_ 0.04259f
C49325 VPWR _0705_/a_59_75# 0.21928f
C49326 _0307_ _0347_ 0.05523f
C49327 comp0.B\[12\] _1044_/a_381_47# 0
C49328 _0371_ _0181_ 0
C49329 _0464_ _0935_/a_27_47# 0.0013f
C49330 _0924_/a_27_47# _0465_ 0.00991f
C49331 _0369_ hold70/a_391_47# 0
C49332 VPWR B[12] 0.28203f
C49333 acc0.A\[7\] input14/a_75_212# 0
C49334 _0464_ _1061_/a_193_47# 0
C49335 _0967_/a_487_297# control0.state\[2\] 0.0141f
C49336 control0.count\[1\] _0167_ 0.01653f
C49337 _0168_ control0.count\[0\] 0.05791f
C49338 _0670_/a_79_21# hold91/a_391_47# 0.00107f
C49339 net1 B[0] 0.0019f
C49340 _1000_/a_193_47# _0347_ 0.26869f
C49341 _0558_/a_68_297# control0.sh 0.01741f
C49342 _0414_ _0994_/a_381_47# 0
C49343 VPWR _1063_/a_193_47# 0.29343f
C49344 _0996_/a_27_47# _1060_/a_27_47# 0
C49345 clkbuf_1_0__f__0458_/a_110_47# _0082_ 0
C49346 hold66/a_49_47# _0237_ 0.00505f
C49347 _0762_/a_297_297# _0103_ 0
C49348 hold23/a_285_47# clknet_1_1__leaf__0457_ 0
C49349 _0195_ net97 0
C49350 _0572_/a_109_47# _0195_ 0.00145f
C49351 _0572_/a_109_297# net155 0.01052f
C49352 _0572_/a_27_297# _0216_ 0.17695f
C49353 clknet_1_0__leaf__0459_ _0869_/a_27_47# 0.00903f
C49354 _0216_ _1006_/a_381_47# 0
C49355 clknet_1_1__leaf__0458_ _0522_/a_27_297# 0
C49356 _0322_ _0219_ 0.06986f
C49357 _0719_/a_27_47# VPWR 0.28551f
C49358 _0476_ _0164_ 0.00561f
C49359 net182 net141 0
C49360 _0180_ net100 0
C49361 VPWR _0460_ 1.55552f
C49362 _0452_ _0261_ 0
C49363 net197 hold9/a_49_47# 0.03032f
C49364 _0432_ _0841_/a_79_21# 0
C49365 clknet_1_0__leaf__0460_ net241 0.00189f
C49366 _0327_ _0219_ 0.04731f
C49367 _0253_ _0435_ 0.00165f
C49368 _0579_/a_109_47# _0461_ 0
C49369 _0212_ comp0.B\[2\] 0
C49370 _1019_/a_193_47# acc0.A\[19\] 0
C49371 clkbuf_1_0__f__0459_/a_110_47# hold19/a_285_47# 0.02551f
C49372 VPWR _1060_/a_193_47# 0.32709f
C49373 net126 clknet_1_0__leaf__0463_ 0.17935f
C49374 _0242_ _0099_ 0
C49375 hold75/a_49_47# _0465_ 0.00306f
C49376 _0856_/a_79_21# _0856_/a_297_297# 0.01735f
C49377 _0474_ _0563_/a_149_47# 0
C49378 _0172_ _0207_ 0
C49379 clkbuf_1_0__f__0457_/a_110_47# _0385_ 0
C49380 VPWR _0988_/a_381_47# 0.07543f
C49381 VPWR _0553_/a_512_297# 0.00875f
C49382 _0327_ _0728_/a_59_75# 0
C49383 _0358_ VPWR 0.29824f
C49384 _1054_/a_634_159# _0186_ 0
C49385 net47 clknet_1_1__leaf__0465_ 0.03806f
C49386 _0520_/a_109_297# net140 0
C49387 _0174_ _1043_/a_193_47# 0.03026f
C49388 net157 _1047_/a_634_159# 0.02514f
C49389 _0216_ _0616_/a_292_297# 0.00272f
C49390 _0305_ _0767_/a_59_75# 0.21182f
C49391 _0457_ VPWR 0.95279f
C49392 clknet_1_0__leaf__0463_ input8/a_75_212# 0.00242f
C49393 _0260_ _0986_/a_193_47# 0
C49394 _1023_/a_1017_47# net177 0
C49395 comp0.B\[10\] _1043_/a_466_413# 0
C49396 _0476_ clknet_0__0463_ 0
C49397 _0581_/a_109_47# _0242_ 0
C49398 _0410_ net5 0.01687f
C49399 hold45/a_49_47# hold45/a_391_47# 0.00188f
C49400 _0476_ hold38/a_391_47# 0.00266f
C49401 _1044_/a_1059_315# net20 0.03392f
C49402 _0670_/a_79_21# _0670_/a_510_47# 0.00844f
C49403 _0670_/a_297_297# _0670_/a_215_47# 0
C49404 _0732_/a_80_21# _0324_ 0.04455f
C49405 _0732_/a_209_297# _0359_ 0.06078f
C49406 _0299_ _0799_/a_209_297# 0
C49407 _0298_ _0799_/a_209_47# 0
C49408 net119 _0163_ 0
C49409 hold59/a_285_47# _0346_ 0
C49410 _0457_ _1015_/a_466_413# 0.00715f
C49411 clkload0/a_27_47# clkload0/X 0.3277f
C49412 net57 _0707_/a_544_297# 0
C49413 _0195_ _0707_/a_201_297# 0
C49414 pp[9] VPWR 1.87472f
C49415 net131 _0142_ 0
C49416 _1018_/a_1059_315# _0393_ 0.00147f
C49417 _0276_ _0795_/a_81_21# 0
C49418 _1037_/a_466_413# B[6] 0
C49419 clknet_0__0458_ _0443_ 0.03684f
C49420 comp0.B\[3\] control0.reset 0
C49421 hold65/a_49_47# _0086_ 0
C49422 net48 _0460_ 0.09189f
C49423 _1001_/a_381_47# VPWR 0.07542f
C49424 hold36/a_391_47# clknet_0__0464_ 0.00779f
C49425 net45 _1017_/a_1059_315# 0.00862f
C49426 _0129_ _1031_/a_1017_47# 0
C49427 _0988_/a_193_47# pp[4] 0
C49428 _0988_/a_381_47# output62/a_27_47# 0
C49429 VPWR _1062_/a_891_413# 0.17282f
C49430 _0616_/a_493_297# _0240_ 0
C49431 _1059_/a_1017_47# net229 0
C49432 _0157_ _0506_/a_384_47# 0
C49433 _0780_/a_285_297# _0347_ 0.0016f
C49434 _0324_ clkbuf_1_0__f__0460_/a_110_47# 0
C49435 _1039_/a_1059_315# _0172_ 0
C49436 _1039_/a_634_159# _0137_ 0.03062f
C49437 _0503_/a_109_297# _0178_ 0.00136f
C49438 _1021_/a_466_413# VPWR 0.25739f
C49439 net243 acc0.A\[25\] 0
C49440 pp[29] net57 0.35522f
C49441 hold57/a_285_47# clkbuf_1_0__f__0463_/a_110_47# 0
C49442 net172 _1037_/a_27_47# 0
C49443 _1038_/a_27_47# _0135_ 0
C49444 acc0.A\[20\] _0462_ 0.05595f
C49445 _0762_/a_215_47# _0762_/a_510_47# 0.00529f
C49446 _0170_ _0466_ 0.08544f
C49447 _0998_/a_634_159# _0410_ 0
C49448 _0585_/a_109_297# _0526_/a_27_47# 0
C49449 _0211_ clknet_1_1__leaf__0463_ 0.00535f
C49450 _0324_ _0250_ 0.22386f
C49451 comp0.B\[5\] net171 0.0027f
C49452 net76 _0658_/a_113_47# 0
C49453 _0984_/a_193_47# clkbuf_1_0__f__0458_/a_110_47# 0.00555f
C49454 _1041_/a_466_413# net172 0
C49455 _0343_ _0246_ 0.02933f
C49456 _0776_/a_27_47# _0306_ 0.00471f
C49457 _0846_/a_149_47# clkbuf_0__0458_/a_110_47# 0
C49458 _0216_ _0360_ 0
C49459 hold10/a_49_47# net36 0.06026f
C49460 _0752_/a_300_297# net49 0
C49461 acc0.A\[16\] _0310_ 0
C49462 _0390_ _0719_/a_27_47# 0
C49463 _0442_ clkbuf_1_0__f__0465_/a_110_47# 0.02328f
C49464 net53 _0352_ 0.02909f
C49465 _1065_/a_466_413# _1065_/a_561_413# 0.00772f
C49466 _1065_/a_634_159# _1065_/a_975_413# 0
C49467 hold5/a_391_47# _0544_/a_51_297# 0.01217f
C49468 net207 hold40/a_49_47# 0
C49469 net105 hold40/a_285_47# 0
C49470 _0183_ _0381_ 0.03018f
C49471 net150 _0382_ 0.28889f
C49472 _0485_ _1066_/a_193_47# 0
C49473 hold66/a_49_47# _1005_/a_27_47# 0
C49474 acc0.A\[27\] _0125_ 0.2508f
C49475 _0817_/a_81_21# _0991_/a_891_413# 0
C49476 _0260_ _0845_/a_109_47# 0.01153f
C49477 _1036_/a_891_413# _1035_/a_466_413# 0.0023f
C49478 _0343_ _0747_/a_510_47# 0
C49479 _0843_/a_68_297# _0843_/a_150_297# 0.00477f
C49480 _0238_ _0618_/a_79_21# 0
C49481 net34 _0482_ 0
C49482 _1068_/a_27_47# _0487_ 0
C49483 _0985_/a_1059_315# _0271_ 0
C49484 _0985_/a_381_47# _0270_ 0
C49485 _0985_/a_891_413# _0256_ 0
C49486 _0306_ _0219_ 0.65188f
C49487 net31 _0548_/a_240_47# 0.08673f
C49488 net24 comp0.B\[5\] 0.02416f
C49489 _0251_ _0399_ 0.09307f
C49490 comp0.B\[11\] _1042_/a_634_159# 0.04526f
C49491 comp0.B\[12\] _1042_/a_193_47# 0
C49492 _0770_/a_79_21# _0241_ 0.00229f
C49493 _1014_/a_634_159# _1014_/a_1059_315# 0
C49494 _1014_/a_27_47# _1014_/a_381_47# 0.05658f
C49495 _1014_/a_193_47# _1014_/a_891_413# 0.19489f
C49496 _0452_ net47 0.05663f
C49497 _0435_ net74 0
C49498 net228 hold82/a_285_47# 0.07986f
C49499 _0269_ acc0.A\[15\] 0.01906f
C49500 VPWR _1047_/a_561_413# 0.0032f
C49501 net59 _0704_/a_68_297# 0.12502f
C49502 _0343_ net235 0
C49503 _1015_/a_27_47# _0173_ 0
C49504 _0130_ _0565_/a_51_297# 0.10389f
C49505 VPWR _0475_ 0.45832f
C49506 _0183_ hold72/a_49_47# 0
C49507 pp[9] input4/a_75_212# 0
C49508 clknet_1_0__leaf__0460_ net177 0
C49509 pp[27] net59 0
C49510 hold101/a_285_47# net248 0.00973f
C49511 _0985_/a_193_47# _0458_ 0.03979f
C49512 comp0.B\[15\] clknet_1_1__leaf__0457_ 0
C49513 VPWR _1007_/a_1017_47# 0
C49514 net180 net174 0.07746f
C49515 net236 _0170_ 0
C49516 _1021_/a_466_413# net48 0
C49517 hold87/a_49_47# _0183_ 0
C49518 clkbuf_1_0__f__0458_/a_110_47# clkbuf_0__0458_/a_110_47# 0.00443f
C49519 VPWR _0796_/a_79_21# 0.49962f
C49520 _1039_/a_634_159# comp0.B\[6\] 0
C49521 output56/a_27_47# acc0.A\[30\] 0
C49522 net120 hold56/a_391_47# 0
C49523 _1055_/a_381_47# net16 0
C49524 net55 _0330_ 0
C49525 _0435_ output61/a_27_47# 0.01206f
C49526 net65 _0830_/a_79_21# 0.05865f
C49527 _0830_/a_215_47# _0989_/a_193_47# 0
C49528 _0830_/a_79_21# _0989_/a_466_413# 0
C49529 _0089_ _0841_/a_297_297# 0
C49530 net52 pp[24] 0.01249f
C49531 hold41/a_285_47# net2 0
C49532 clkbuf_1_0__f__0459_/a_110_47# _1017_/a_634_159# 0
C49533 _0956_/a_220_297# comp0.B\[0\] 0.01255f
C49534 net44 _0218_ 0.21182f
C49535 _1018_/a_891_413# net103 0
C49536 _0802_/a_59_75# _0218_ 0.03592f
C49537 _0664_/a_79_21# _0286_ 0.00168f
C49538 _0664_/a_382_297# _0283_ 0
C49539 _0338_ _0334_ 0.06956f
C49540 _0440_ net73 0
C49541 net58 _0399_ 1.2527f
C49542 net112 _1025_/a_381_47# 0
C49543 _1026_/a_634_159# acc0.A\[25\] 0.00772f
C49544 _0317_ _0739_/a_79_21# 0
C49545 hold18/a_49_47# _0846_/a_51_297# 0
C49546 _1032_/a_27_47# _0181_ 0.03813f
C49547 _0402_ VPWR 0.61195f
C49548 hold78/a_285_47# hold78/a_391_47# 0.41909f
C49549 pp[10] clknet_1_1__leaf__0465_ 0.00131f
C49550 clkbuf_1_0__f__0463_/a_110_47# _0159_ 0
C49551 _0819_/a_81_21# _0819_/a_384_47# 0.00138f
C49552 _0274_ acc0.A\[8\] 0.21364f
C49553 _0275_ net66 0
C49554 _0959_/a_300_47# control0.sh 0
C49555 net137 _0194_ 0.01419f
C49556 _0441_ _0431_ 0
C49557 _0316_ _0333_ 0
C49558 _0343_ net103 0.0452f
C49559 net53 _0574_/a_109_297# 0
C49560 _1033_/a_27_47# _0564_/a_68_297# 0
C49561 hold47/a_49_47# VPWR 0.27859f
C49562 hold41/a_391_47# net3 0
C49563 net87 clknet_1_0__leaf__0457_ 0
C49564 net34 _0476_ 0
C49565 _0985_/a_975_413# net61 0
C49566 net17 _0171_ 0.00101f
C49567 clknet_0__0463_ clkbuf_0__0463_/a_110_47# 1.74109f
C49568 _0195_ _1010_/a_27_47# 0
C49569 _0415_ _0647_/a_47_47# 0
C49570 _0275_ _0991_/a_27_47# 0
C49571 clknet_1_0__leaf__0459_ _1060_/a_193_47# 0.00112f
C49572 net11 _0193_ 0.02121f
C49573 acc0.A\[29\] net116 0.00246f
C49574 _0387_ _0309_ 0
C49575 _1050_/a_1059_315# net135 0
C49576 _1033_/a_27_47# clknet_1_1__leaf_clk 0
C49577 _0222_ _1022_/a_381_47# 0
C49578 _0454_ _0455_ 0.29521f
C49579 net234 net149 0.10418f
C49580 _0402_ _0654_/a_27_413# 0
C49581 _0855_/a_81_21# _0112_ 0
C49582 _0174_ control0.sh 0.02179f
C49583 _1037_/a_27_47# _1036_/a_891_413# 0
C49584 _1037_/a_193_47# _1036_/a_1059_315# 0
C49585 _0481_ _1070_/a_1059_315# 0
C49586 _0963_/a_117_297# VPWR 0.00852f
C49587 _0955_/a_32_297# _1062_/a_27_47# 0
C49588 _0179_ _0269_ 0.01782f
C49589 _0836_/a_150_297# _0437_ 0
C49590 _0223_ _0741_/a_109_297# 0
C49591 _0817_/a_266_47# _0290_ 0.00115f
C49592 _0817_/a_266_297# _0425_ 0.00509f
C49593 _0300_ _0668_/a_382_297# 0
C49594 _0277_ _0668_/a_79_21# 0.04842f
C49595 _0999_/a_891_413# _0352_ 0
C49596 _0457_ clknet_1_0__leaf__0459_ 0.00463f
C49597 _1013_/a_634_159# pp[31] 0
C49598 _0498_/a_51_297# net247 0.12258f
C49599 net46 net149 0
C49600 _0470_ clkbuf_1_1__f_clk/a_110_47# 0
C49601 _0640_/a_465_297# _0255_ 0
C49602 _0820_/a_215_47# _0428_ 0.00673f
C49603 net31 net7 0.13402f
C49604 _0730_/a_215_47# acc0.A\[29\] 0
C49605 _0179_ _0189_ 0.13575f
C49606 comp0.B\[2\] _1033_/a_466_413# 0.05184f
C49607 _0680_/a_217_297# _0392_ 0
C49608 _0464_ clkbuf_0__0464_/a_110_47# 0.31602f
C49609 net150 _1005_/a_634_159# 0.00384f
C49610 acc0.A\[22\] _1005_/a_27_47# 0
C49611 _0217_ _1005_/a_193_47# 0
C49612 _0138_ net10 0
C49613 acc0.A\[29\] hold92/a_285_47# 0
C49614 net190 _1028_/a_466_413# 0.04281f
C49615 _0126_ _1028_/a_27_47# 0.15853f
C49616 _0216_ _1014_/a_1059_315# 0
C49617 _0180_ net148 0.0108f
C49618 _0955_/a_32_297# _0561_/a_51_297# 0.00187f
C49619 _0293_ _0218_ 0
C49620 _0350_ _0738_/a_150_297# 0
C49621 net71 _0465_ 0
C49622 _0275_ _0350_ 0.02736f
C49623 comp0.B\[13\] _1043_/a_193_47# 0
C49624 _0489_ _0488_ 0
C49625 _0576_/a_109_297# net177 0
C49626 _1022_/a_466_413# _0103_ 0
C49627 _0342_ net99 0
C49628 _1003_/a_634_159# clknet_1_0__leaf__0460_ 0.0098f
C49629 net34 hold89/a_285_47# 0.00364f
C49630 control0.state\[1\] hold89/a_391_47# 0.02566f
C49631 _0686_/a_219_297# _0686_/a_27_53# 0.10125f
C49632 clkbuf_0__0462_/a_110_47# hold90/a_391_47# 0.00262f
C49633 net61 _0641_/a_113_47# 0
C49634 _1059_/a_634_159# acc0.A\[15\] 0.00412f
C49635 _1019_/a_193_47# net1 0
C49636 _0643_/a_103_199# _0986_/a_193_47# 0
C49637 _0278_ clknet_1_1__leaf__0459_ 0.01876f
C49638 acc0.A\[2\] net71 0.13783f
C49639 _1018_/a_193_47# _0116_ 0.58202f
C49640 _0319_ _0106_ 0
C49641 _0366_ acc0.A\[25\] 0.17054f
C49642 A[12] _0186_ 0.03133f
C49643 B[8] A[15] 0.20439f
C49644 _1008_/a_1059_315# _1008_/a_891_413# 0.31086f
C49645 _1008_/a_193_47# _1008_/a_975_413# 0
C49646 _1008_/a_466_413# _1008_/a_381_47# 0.03733f
C49647 _1055_/a_27_47# _1055_/a_634_159# 0.14145f
C49648 _0648_/a_205_297# VPWR 0.00165f
C49649 _0505_/a_27_297# _0505_/a_109_297# 0.17136f
C49650 _0718_/a_285_47# _1011_/a_1059_315# 0
C49651 pp[27] _0335_ 0.01385f
C49652 pp[16] _0995_/a_27_47# 0
C49653 _1020_/a_634_159# _0118_ 0.04547f
C49654 net53 _1025_/a_466_413# 0.00631f
C49655 _0250_ _0347_ 0
C49656 _0133_ _0955_/a_32_297# 0
C49657 _1035_/a_975_413# comp0.B\[3\] 0
C49658 _0369_ _1009_/a_27_47# 0
C49659 _0311_ _0350_ 0
C49660 _0215_ _0173_ 0.1181f
C49661 _1016_/a_193_47# _0114_ 0
C49662 _0239_ acc0.A\[16\] 0.05977f
C49663 _0230_ _0234_ 0.06878f
C49664 VPWR _0614_/a_29_53# 0.17739f
C49665 net64 _0274_ 0.00491f
C49666 net59 _0216_ 0.44191f
C49667 pp[30] _0195_ 0.05837f
C49668 _0104_ clkbuf_1_0__f__0460_/a_110_47# 0.0035f
C49669 net216 clknet_0__0460_ 0
C49670 _0537_/a_68_297# comp0.B\[14\] 0
C49671 _0346_ _0219_ 0.03371f
C49672 acc0.A\[27\] _1009_/a_891_413# 0
C49673 clknet_0__0458_ _0986_/a_891_413# 0.00179f
C49674 hold69/a_285_47# _0748_/a_81_21# 0
C49675 _0174_ net157 0.12561f
C49676 clknet_0__0457_ _1014_/a_891_413# 0
C49677 _0183_ clknet_0__0461_ 0.0074f
C49678 _0515_/a_384_47# net181 0.0101f
C49679 acc0.A\[17\] net219 0
C49680 control0.sh _0208_ 0.07f
C49681 _0627_/a_215_53# _0432_ 0
C49682 _0104_ _0250_ 0.02606f
C49683 _1054_/a_1059_315# _0518_/a_27_297# 0
C49684 net84 _1017_/a_193_47# 0
C49685 _1032_/a_466_413# comp0.B\[0\] 0
C49686 _1041_/a_891_413# _0137_ 0
C49687 _1041_/a_561_413# _0172_ 0
C49688 _0997_/a_466_413# _0345_ 0.01316f
C49689 VPWR net27 0.60288f
C49690 net63 _0834_/a_109_297# 0.00405f
C49691 _0504_/a_27_47# _0982_/a_27_47# 0.00108f
C49692 _0101_ _0466_ 0
C49693 _0462_ _1007_/a_891_413# 0
C49694 _0846_/a_512_297# _0449_ 0.00208f
C49695 _0182_ clkbuf_1_1__f__0457_/a_110_47# 0.03552f
C49696 _0533_/a_109_47# clknet_1_1__leaf__0457_ 0
C49697 net197 _0739_/a_79_21# 0
C49698 clknet_1_1__leaf__0457_ hold71/a_285_47# 0.00222f
C49699 hold94/a_391_47# _0377_ 0
C49700 hold94/a_49_47# _0219_ 0.06992f
C49701 hold94/a_285_47# net241 0.02654f
C49702 _0991_/a_381_47# acc0.A\[15\] 0
C49703 net92 _0771_/a_215_297# 0
C49704 _0826_/a_27_53# _0434_ 0.01202f
C49705 _0217_ _0264_ 0.0302f
C49706 net66 _0510_/a_109_47# 0
C49707 _0506_/a_299_297# _0505_/a_27_297# 0
C49708 _0506_/a_81_21# _0505_/a_109_297# 0
C49709 _0473_ net29 0
C49710 _0982_/a_27_47# _0456_ 0.01054f
C49711 _0504_/a_27_47# _0145_ 0
C49712 _0982_/a_466_413# net234 0
C49713 _0559_/a_51_297# net185 0
C49714 net161 B[1] 0.00109f
C49715 comp0.B\[4\] input24/a_75_212# 0.00147f
C49716 _0294_ clknet_1_1__leaf__0465_ 0.0566f
C49717 _0305_ _0290_ 0
C49718 hold42/a_285_47# _1058_/a_381_47# 0.00206f
C49719 _1058_/a_381_47# _1057_/a_1059_315# 0
C49720 _1058_/a_1059_315# _1057_/a_381_47# 0
C49721 hold65/a_285_47# clknet_1_0__leaf__0465_ 0
C49722 _0298_ _0668_/a_79_21# 0.12955f
C49723 _0745_/a_109_47# _0250_ 0
C49724 _0210_ net8 0
C49725 _0280_ hold81/a_285_47# 0
C49726 clknet_1_0__leaf__0459_ _0796_/a_79_21# 0
C49727 net49 net1 0
C49728 _0179_ _1059_/a_634_159# 0
C49729 hold26/a_285_47# net174 0
C49730 _0343_ output41/a_27_47# 0.0063f
C49731 _0259_ clkbuf_1_1__f__0465_/a_110_47# 0.00976f
C49732 _1000_/a_592_47# _0352_ 0.00297f
C49733 _0701_/a_303_47# _0350_ 0.00241f
C49734 hold33/a_285_47# clkbuf_1_0__f__0463_/a_110_47# 0
C49735 _0315_ _0737_/a_35_297# 0
C49736 _0216_ _0124_ 0.04775f
C49737 VPWR _0470_ 0.3415f
C49738 _1016_/a_466_413# clknet_1_1__leaf__0461_ 0.03862f
C49739 clknet_1_1__leaf__0458_ _0193_ 0.00247f
C49740 _0369_ _0771_/a_27_413# 0
C49741 VPWR _1017_/a_1059_315# 0.37796f
C49742 _0504_/a_27_47# _0446_ 0
C49743 _1037_/a_466_413# comp0.B\[5\] 0
C49744 clk clknet_0_clk 0.00466f
C49745 _0563_/a_51_297# _0563_/a_149_47# 0.02487f
C49746 _0343_ _0723_/a_207_413# 0.01344f
C49747 _0506_/a_81_21# _0506_/a_299_297# 0.08213f
C49748 _0804_/a_215_47# VPWR 0.00926f
C49749 _1056_/a_891_413# A[10] 0
C49750 acc0.A\[29\] hold80/a_285_47# 0.0111f
C49751 net157 _0208_ 0.03662f
C49752 _1017_/a_634_159# clkbuf_0__0461_/a_110_47# 0
C49753 VPWR _1033_/a_193_47# 0.29864f
C49754 _0456_ _0446_ 0
C49755 _1038_/a_193_47# comp0.B\[8\] 0
C49756 VPWR _0136_ 0.37373f
C49757 clknet_1_1__leaf__0460_ _0574_/a_27_297# 0
C49758 _0243_ _0614_/a_111_297# 0.00224f
C49759 clknet_1_0__leaf__0465_ _1049_/a_193_47# 0.00336f
C49760 _0732_/a_209_297# _0325_ 0
C49761 _0251_ _0619_/a_68_297# 0.13386f
C49762 _0291_ _0181_ 0.04806f
C49763 net140 _0186_ 0
C49764 clkbuf_1_1__f__0462_/a_110_47# _0352_ 0.00256f
C49765 _0402_ _0283_ 0.1826f
C49766 _0372_ _0392_ 0
C49767 VPWR _1050_/a_891_413# 0.19134f
C49768 _0342_ _0396_ 0
C49769 _0511_/a_299_297# net192 0.05973f
C49770 comp0.B\[10\] net196 0
C49771 hold45/a_391_47# _0156_ 0.00305f
C49772 _1010_/a_634_159# _1010_/a_466_413# 0.23992f
C49773 _1010_/a_193_47# _1010_/a_1059_315# 0.03405f
C49774 _1010_/a_27_47# _1010_/a_891_413# 0.03224f
C49775 net166 _0181_ 0
C49776 clknet_1_0__leaf__0462_ _1004_/a_634_159# 0.00437f
C49777 _0644_/a_285_47# acc0.A\[15\] 0.03629f
C49778 _0717_/a_80_21# _0195_ 0
C49779 _0717_/a_209_297# net57 0
C49780 _0517_/a_81_21# net66 0
C49781 _0991_/a_634_159# _0181_ 0.02096f
C49782 net54 _1028_/a_27_47# 0
C49783 net134 net10 0
C49784 _1040_/a_27_47# _1040_/a_634_159# 0.13601f
C49785 _0329_ _0318_ 0.00244f
C49786 _0457_ _0113_ 0.03292f
C49787 _0198_ _1048_/a_891_413# 0
C49788 _0146_ _1048_/a_634_159# 0.0466f
C49789 _0432_ _0837_/a_81_21# 0
C49790 _0195_ _0339_ 0.41101f
C49791 _0238_ _0242_ 0
C49792 _1002_/a_466_413# _0217_ 0.01541f
C49793 _0472_ _0913_/a_27_47# 0.02064f
C49794 _0135_ B[6] 0
C49795 _1002_/a_1059_315# net150 0.02656f
C49796 _1002_/a_193_47# _0183_ 0.02968f
C49797 _0746_/a_81_21# _0346_ 0.19781f
C49798 B[13] input32/a_75_212# 0.00649f
C49799 input21/a_75_212# B[9] 0
C49800 _0665_/a_109_297# A[13] 0
C49801 hold54/a_285_47# _0181_ 0
C49802 _0234_ _0236_ 0.08971f
C49803 _1020_/a_381_47# _0461_ 0
C49804 _0846_/a_51_297# _0846_/a_245_297# 0.01218f
C49805 _0178_ _0526_/a_27_47# 0.22772f
C49806 net45 _1016_/a_27_47# 0.00258f
C49807 _1067_/a_27_47# _1067_/a_634_159# 0.14145f
C49808 _0174_ _0550_/a_240_47# 0.02471f
C49809 _0082_ acc0.A\[15\] 0.01848f
C49810 _0280_ _0282_ 0
C49811 net125 _0137_ 0
C49812 _0119_ VPWR 0.54634f
C49813 _0221_ _0703_/a_109_297# 0
C49814 net84 _0410_ 0
C49815 _0343_ _0102_ 0
C49816 net9 _0178_ 0.01017f
C49817 _1072_/a_27_47# _1071_/a_634_159# 0
C49818 _0575_/a_27_297# _0352_ 0
C49819 _0647_/a_47_47# _0347_ 0
C49820 _1009_/a_193_47# _1009_/a_381_47# 0.10164f
C49821 _1009_/a_634_159# _1009_/a_891_413# 0.03684f
C49822 _1009_/a_27_47# _1009_/a_561_413# 0.0027f
C49823 _0989_/a_27_47# _0989_/a_193_47# 0.96469f
C49824 hold1/a_49_47# hold1/a_285_47# 0.22264f
C49825 _0645_/a_47_47# _1059_/a_1059_315# 0
C49826 clkload2/Y net134 0
C49827 clknet_1_1__leaf__0460_ _0326_ 0.49017f
C49828 _0154_ _0186_ 0
C49829 _1065_/a_1059_315# control0.reset 0.09877f
C49830 hold5/a_49_47# _0140_ 0
C49831 acc0.A\[17\] _0352_ 0.02762f
C49832 _0982_/a_1059_315# VPWR 0.39953f
C49833 _0399_ _0831_/a_285_297# 0.04527f
C49834 _0476_ _1066_/a_466_413# 0.00638f
C49835 net213 _1005_/a_1059_315# 0
C49836 _0992_/a_27_47# _0992_/a_193_47# 0.97438f
C49837 _0817_/a_368_297# _0089_ 0
C49838 net31 _0202_ 0
C49839 _1036_/a_381_47# net121 0.00256f
C49840 comp0.B\[4\] _1035_/a_634_159# 0
C49841 _1036_/a_891_413# _0133_ 0
C49842 _0517_/a_81_21# _0350_ 0
C49843 net111 _1025_/a_381_47# 0
C49844 net7 _0548_/a_240_47# 0
C49845 net35 _0466_ 0.13841f
C49846 VPWR _1053_/a_27_47# 0.69398f
C49847 acc0.A\[27\] _1027_/a_634_159# 0
C49848 _0131_ net201 0
C49849 _1032_/a_634_159# net118 0
C49850 hold79/a_49_47# control0.count\[1\] 0.28664f
C49851 _0557_/a_512_297# _0211_ 0
C49852 comp0.B\[11\] net128 0.19809f
C49853 _1018_/a_891_413# _0774_/a_68_297# 0
C49854 _1014_/a_27_47# acc0.A\[0\] 0.00133f
C49855 _1071_/a_634_159# _1071_/a_592_47# 0
C49856 _1014_/a_1059_315# net100 0
C49857 _0996_/a_27_47# _0094_ 0.14219f
C49858 _0996_/a_634_159# _0410_ 0
C49859 _0996_/a_466_413# net238 0.04016f
C49860 _1045_/a_27_47# _1043_/a_27_47# 0
C49861 _0311_ _0244_ 0
C49862 _1015_/a_975_413# _0208_ 0.00127f
C49863 net61 _0435_ 0.03428f
C49864 _0343_ _0774_/a_68_297# 0.0099f
C49865 hold10/a_285_47# hold10/a_391_47# 0.41909f
C49866 _0178_ _0175_ 0
C49867 _1035_/a_891_413# net26 0.00278f
C49868 _0119_ net48 0.00253f
C49869 _0290_ _0181_ 0.06746f
C49870 _0113_ _0475_ 0
C49871 _0195_ _1026_/a_193_47# 0
C49872 net155 _1026_/a_27_47# 0
C49873 input23/a_75_212# B[3] 0
C49874 B[15] input26/a_75_212# 0
C49875 net157 _1046_/a_193_47# 0
C49876 _0176_ clknet_1_1__leaf__0457_ 0
C49877 _0553_/a_51_297# comp0.B\[5\] 0
C49878 _0350_ hold50/a_49_47# 0
C49879 acc0.A\[12\] acc0.A\[9\] 0
C49880 hold79/a_285_47# clkbuf_1_0__f_clk/a_110_47# 0.00193f
C49881 _0348_ _0334_ 0.03628f
C49882 _0216_ _1024_/a_466_413# 0.00195f
C49883 _0252_ _0437_ 0.02434f
C49884 acc0.A\[7\] _0087_ 0
C49885 _0087_ _0989_/a_1059_315# 0
C49886 _0437_ _0989_/a_381_47# 0.0082f
C49887 acc0.A\[24\] _1006_/a_193_47# 0
C49888 _0305_ _1059_/a_592_47# 0
C49889 _0179_ _0082_ 0
C49890 clkbuf_1_0__f__0459_/a_110_47# net103 0
C49891 _0457_ comp0.B\[3\] 0
C49892 _0479_ _0484_ 0.02616f
C49893 VPWR _0451_ 0.18475f
C49894 _1020_/a_193_47# acc0.A\[20\] 0.00477f
C49895 net2 net4 0.00111f
C49896 net112 acc0.A\[25\] 0.08778f
C49897 net36 _1039_/a_975_413# 0.00155f
C49898 net88 _1067_/a_975_413# 0
C49899 _0389_ _0391_ 0.24939f
C49900 _0243_ net223 0.04253f
C49901 _1002_/a_1059_315# control0.add 0
C49902 _1042_/a_27_47# _0203_ 0
C49903 _1012_/a_561_413# _0352_ 0
C49904 _0343_ pp[6] 0
C49905 _0555_/a_51_297# _0175_ 0
C49906 _0869_/a_27_47# _0345_ 0
C49907 acc0.A\[25\] acc0.A\[24\] 0.30403f
C49908 acc0.A\[12\] _0670_/a_79_21# 0
C49909 _0343_ _1016_/a_592_47# 0
C49910 net63 net9 0
C49911 _1033_/a_1059_315# _0215_ 0.01743f
C49912 _0172_ _0472_ 0.09551f
C49913 _0137_ _0473_ 0.03511f
C49914 _0984_/a_193_47# acc0.A\[15\] 0.01f
C49915 clknet_1_0__leaf__0459_ _1017_/a_1059_315# 0
C49916 acc0.A\[22\] _0222_ 0.31586f
C49917 hold36/a_391_47# comp0.B\[14\] 0.06703f
C49918 _1069_/a_27_47# _1069_/a_466_413# 0.26957f
C49919 _1069_/a_193_47# _1069_/a_634_159# 0.12729f
C49920 _0229_ net46 0
C49921 _0786_/a_217_297# _0295_ 0.01496f
C49922 _1052_/a_592_47# _0180_ 0
C49923 _0786_/a_80_21# _0304_ 0
C49924 _0320_ _0686_/a_219_297# 0
C49925 _0192_ VPWR 0.17362f
C49926 hold60/a_49_47# hold60/a_285_47# 0.22264f
C49927 net56 _0705_/a_59_75# 0
C49928 _0954_/a_32_297# _0954_/a_114_297# 0.01439f
C49929 _0320_ _1008_/a_1059_315# 0
C49930 _0225_ _0606_/a_392_297# 0
C49931 _0474_ _1062_/a_27_47# 0
C49932 hold66/a_285_47# _0762_/a_79_21# 0
C49933 _0334_ _0332_ 0
C49934 hold10/a_49_47# _1039_/a_27_47# 0
C49935 acc0.A\[27\] _1026_/a_891_413# 0
C49936 acc0.A\[27\] clkbuf_1_1__f__0460_/a_110_47# 0.02857f
C49937 acc0.A\[1\] _0181_ 0.60159f
C49938 output48/a_27_47# output49/a_27_47# 0
C49939 _1059_/a_27_47# hold82/a_49_47# 0.00533f
C49940 _0512_/a_109_47# acc0.A\[11\] 0.00165f
C49941 comp0.B\[7\] hold25/a_391_47# 0
C49942 _1030_/a_466_413# hold62/a_285_47# 0.0041f
C49943 _1030_/a_1059_315# hold62/a_49_47# 0
C49944 _1030_/a_634_159# hold62/a_391_47# 0
C49945 _0311_ _0731_/a_299_297# 0
C49946 net69 _0218_ 0.00309f
C49947 B[5] net28 0.00314f
C49948 _0985_/a_466_413# _0350_ 0
C49949 net22 net32 0.06891f
C49950 _0780_/a_35_297# clknet_0__0461_ 0
C49951 _0084_ _0986_/a_561_413# 0
C49952 _0445_ _0986_/a_592_47# 0
C49953 _0579_/a_373_47# _0457_ 0
C49954 clknet_1_1__leaf__0460_ acc0.A\[28\] 0.18921f
C49955 hold96/a_391_47# _1024_/a_466_413# 0
C49956 comp0.B\[2\] _0131_ 0.18762f
C49957 net172 _0174_ 0
C49958 _0577_/a_27_297# _1022_/a_27_47# 0
C49959 net150 net91 0.2251f
C49960 net14 A[7] 0.18821f
C49961 _0225_ net49 0
C49962 clknet_1_0__leaf__0462_ net46 0.04672f
C49963 clkload1/Y _0258_ 0.01209f
C49964 _0195_ acc0.A\[0\] 0
C49965 _0538_/a_51_297# _0538_/a_245_297# 0.01218f
C49966 _0462_ _0772_/a_297_297# 0
C49967 _0787_/a_80_21# _0345_ 0.00105f
C49968 clknet_1_1__leaf__0462_ _1008_/a_891_413# 0.00237f
C49969 _0474_ _0561_/a_51_297# 0.00575f
C49970 _1032_/a_1059_315# _0565_/a_240_47# 0
C49971 _0955_/a_32_297# _0208_ 0.00132f
C49972 comp0.B\[5\] _0561_/a_149_47# 0
C49973 net163 clknet_1_1__leaf__0462_ 0.00503f
C49974 net61 _0456_ 0
C49975 output67/a_27_47# net189 0.00226f
C49976 pp[9] _1057_/a_592_47# 0
C49977 net21 hold51/a_49_47# 0
C49978 VPWR _1046_/a_381_47# 0.07064f
C49979 _1022_/a_466_413# _1022_/a_381_47# 0.03733f
C49980 _1022_/a_193_47# _1022_/a_975_413# 0
C49981 _1022_/a_1059_315# _1022_/a_891_413# 0.31086f
C49982 clknet_1_0__leaf__0463_ net8 0.08217f
C49983 _0645_/a_285_47# _0644_/a_129_47# 0
C49984 hold22/a_285_47# _0518_/a_27_297# 0
C49985 _0314_ _0681_/a_113_47# 0
C49986 net89 clknet_1_0__leaf__0460_ 0.16316f
C49987 hold49/a_391_47# _0172_ 0.04453f
C49988 _0633_/a_109_297# _0345_ 0
C49989 net145 acc0.A\[15\] 0.004f
C49990 _0994_/a_27_47# _0994_/a_634_159# 0.14145f
C49991 clknet_1_0__leaf__0463_ net32 0
C49992 _0358_ net56 0
C49993 clkbuf_1_1__f__0460_/a_110_47# _0364_ 0
C49994 _0275_ _0986_/a_634_159# 0.04072f
C49995 _0779_/a_79_21# _0779_/a_297_297# 0.01735f
C49996 _0473_ comp0.B\[6\] 0.22491f
C49997 net211 _1001_/a_466_413# 0.0435f
C49998 _0292_ _0812_/a_215_47# 0.00278f
C49999 _0217_ _0385_ 0
C50000 _1055_/a_891_413# _1055_/a_975_413# 0.00851f
C50001 _1055_/a_27_47# net141 0.22831f
C50002 _1055_/a_381_47# _1055_/a_561_413# 0.00123f
C50003 _0505_/a_373_47# net6 0.00194f
C50004 _0505_/a_109_297# _0184_ 0.00339f
C50005 VPWR _0373_ 0.57683f
C50006 hold24/a_285_47# comp0.B\[7\] 0.00308f
C50007 _0718_/a_47_47# _0195_ 0
C50008 output53/a_27_47# acc0.A\[25\] 0
C50009 _0305_ _0656_/a_59_75# 0
C50010 _0467_ clknet_1_1__leaf__0463_ 0
C50011 hold88/a_49_47# VPWR 0.31537f
C50012 _0984_/a_193_47# _0179_ 0.00209f
C50013 VPWR _0758_/a_297_297# 0.0103f
C50014 _0133_ _0474_ 0.05977f
C50015 hold79/a_285_47# control0.count\[2\] 0
C50016 net157 comp0.B\[9\] 0
C50017 hold14/a_391_47# _1036_/a_466_413# 0
C50018 hold14/a_49_47# _1036_/a_891_413# 0
C50019 _1003_/a_634_159# _1003_/a_592_47# 0
C50020 _0218_ _0840_/a_150_297# 0
C50021 _1055_/a_1017_47# net181 0
C50022 hold59/a_285_47# net221 0
C50023 _1036_/a_27_47# net27 0
C50024 _1036_/a_193_47# B[4] 0
C50025 _0456_ _1019_/a_634_159# 0
C50026 net234 _1019_/a_891_413# 0
C50027 net101 clknet_1_0__leaf__0461_ 0.14945f
C50028 _0749_/a_81_21# _0384_ 0
C50029 clknet_1_0__leaf__0458_ clknet_1_1__leaf__0457_ 0
C50030 hold45/a_285_47# _1058_/a_27_47# 0
C50031 _0207_ _1040_/a_193_47# 0.00137f
C50032 comp0.B\[12\] clknet_1_1__leaf__0464_ 0.46868f
C50033 VPWR _0485_ 0.90789f
C50034 hold33/a_391_47# _0548_/a_51_297# 0.01217f
C50035 clknet_1_0__leaf__0460_ hold4/a_49_47# 0
C50036 _0343_ _0815_/a_113_297# 0
C50037 hold58/a_391_47# net205 0.1435f
C50038 _0176_ net19 0.39062f
C50039 clkbuf_0__0461_/a_110_47# _0246_ 0
C50040 hold20/a_285_47# clknet_0_clk 0.01129f
C50041 hold46/a_49_47# net180 0
C50042 hold16/a_285_47# net239 0
C50043 net22 _1042_/a_1059_315# 0
C50044 _0211_ input28/a_75_212# 0
C50045 _1054_/a_1059_315# _0191_ 0.00908f
C50046 _0217_ _0856_/a_79_21# 0
C50047 net202 comp0.B\[0\] 0
C50048 net234 net206 0.01304f
C50049 clknet_1_1__leaf__0463_ comp0.B\[0\] 0.39672f
C50050 _1004_/a_466_413# _0102_ 0.042f
C50051 _1004_/a_1059_315# _0352_ 0
C50052 _0852_/a_35_297# acc0.A\[0\] 0
C50053 _0502_/a_27_47# net133 0.00415f
C50054 _0983_/a_193_47# _0347_ 0.03711f
C50055 clknet_1_1__leaf__0461_ _0408_ 0
C50056 net67 acc0.A\[15\] 0
C50057 _0603_/a_68_297# _0765_/a_79_21# 0.01992f
C50058 net23 _1065_/a_634_159# 0.02036f
C50059 net172 _0208_ 0
C50060 VPWR _0271_ 0.47244f
C50061 _0506_/a_299_297# _0184_ 0.03118f
C50062 _1054_/a_381_47# _1053_/a_1059_315# 0
C50063 _0765_/a_79_21# hold73/a_391_47# 0
C50064 _0370_ clknet_0__0460_ 0
C50065 _0080_ net234 0
C50066 _0195_ _0580_/a_109_297# 0.00422f
C50067 _0285_ _0404_ 0
C50068 net22 net10 0.00218f
C50069 _0222_ _0379_ 0
C50070 _0664_/a_382_297# _0345_ 0
C50071 net90 _1024_/a_891_413# 0.00101f
C50072 VPWR _0987_/a_891_413# 0.20168f
C50073 _0179_ clkbuf_0__0458_/a_110_47# 0
C50074 _1024_/a_27_47# _1024_/a_1059_315# 0.04875f
C50075 _1024_/a_193_47# _1024_/a_466_413# 0.08301f
C50076 _1058_/a_561_413# net189 0.00167f
C50077 net245 _0400_ 0.00192f
C50078 hold93/a_49_47# hold93/a_391_47# 0.00188f
C50079 _0557_/a_149_47# net160 0.01062f
C50080 _0414_ _0218_ 0.025f
C50081 hold58/a_285_47# _0211_ 0.00351f
C50082 _0816_/a_68_297# _0423_ 0
C50083 net48 _0373_ 0.02495f
C50084 _0287_ _0347_ 0.06304f
C50085 _0643_/a_253_47# _0449_ 0
C50086 _1011_/a_27_47# _0333_ 0.00192f
C50087 VPWR _0727_/a_109_47# 0
C50088 _0179_ net145 0.2764f
C50089 _0985_/a_27_47# _0182_ 0
C50090 _0458_ _0636_/a_59_75# 0.01098f
C50091 acc0.A\[14\] _0266_ 0
C50092 VPWR A[5] 0.2224f
C50093 _1000_/a_891_413# _0244_ 0.00668f
C50094 _1000_/a_466_413# _0388_ 0.00288f
C50095 _1000_/a_1059_315# _0386_ 0
C50096 VPWR _1029_/a_891_413# 0.21184f
C50097 _0540_/a_51_297# _0540_/a_149_47# 0.02487f
C50098 _0982_/a_1059_315# _0453_ 0
C50099 net166 clknet_1_1__leaf__0461_ 0.09502f
C50100 _1048_/a_634_159# _1048_/a_381_47# 0
C50101 _1034_/a_634_159# clknet_1_1__leaf__0463_ 0.01108f
C50102 clkbuf_1_1__f__0460_/a_110_47# _1010_/a_193_47# 0.00119f
C50103 clknet_1_0__leaf__0463_ net10 0.00596f
C50104 net29 comp0.B\[8\] 0
C50105 _0399_ _0796_/a_215_47# 0.04593f
C50106 _0218_ net102 0
C50107 clkbuf_1_0__f__0461_/a_110_47# _0242_ 0.1289f
C50108 _0135_ comp0.B\[5\] 0.23616f
C50109 VPWR _1016_/a_27_47# 0.45538f
C50110 _0378_ _0103_ 0.04568f
C50111 _0348_ _0724_/a_113_297# 0
C50112 _0846_/a_51_297# _0448_ 0.07631f
C50113 _0501_/a_27_47# clknet_0__0463_ 0.00199f
C50114 _0556_/a_68_297# _0211_ 0.10711f
C50115 _0981_/a_109_47# clknet_1_0__leaf_clk 0.00151f
C50116 _0640_/a_215_297# _0434_ 0
C50117 clknet_0__0457_ _0580_/a_27_297# 0
C50118 _0460_ _0345_ 0.03538f
C50119 net103 clkbuf_0__0461_/a_110_47# 0.00145f
C50120 _0770_/a_79_21# _0352_ 0
C50121 _0290_ hold82/a_391_47# 0
C50122 _0313_ _0317_ 0.00103f
C50123 _0427_ _0818_/a_109_47# 0.0111f
C50124 comp0.B\[14\] net180 0
C50125 _0130_ VPWR 0.49307f
C50126 _0670_/a_79_21# net42 0.06548f
C50127 _0518_/a_373_47# acc0.A\[6\] 0
C50128 hold69/a_49_47# _0246_ 0
C50129 net36 net47 0.20097f
C50130 _0137_ _0497_/a_68_297# 0
C50131 _0217_ _0454_ 0
C50132 net32 _0544_/a_245_297# 0.00109f
C50133 net152 _0544_/a_512_297# 0
C50134 _0981_/a_27_297# _0974_/a_79_199# 0
C50135 _0179_ _0152_ 0.04698f
C50136 _0607_/a_27_297# _0677_/a_47_47# 0.00625f
C50137 net45 _0400_ 0
C50138 pp[30] hold15/a_49_47# 0.01114f
C50139 net59 hold15/a_391_47# 0
C50140 _1010_/a_466_413# net96 0
C50141 _0179_ net67 0.11403f
C50142 _0248_ _0385_ 0
C50143 _0130_ _1015_/a_466_413# 0
C50144 _0457_ _0345_ 0
C50145 net77 _0181_ 0
C50146 _0465_ _0434_ 0
C50147 _1040_/a_381_47# _1040_/a_561_413# 0.00123f
C50148 _1040_/a_891_413# _1040_/a_975_413# 0.00851f
C50149 hold74/a_391_47# acc0.A\[16\] 0.06379f
C50150 net98 _0350_ 0
C50151 hold13/a_285_47# _0137_ 0
C50152 _0795_/a_81_21# _0409_ 0.00221f
C50153 _0979_/a_27_297# net164 0.1221f
C50154 _0979_/a_109_297# _0480_ 0.01155f
C50155 _1017_/a_193_47# acc0.A\[18\] 0
C50156 _0146_ net134 0.01057f
C50157 _0322_ _0328_ 0.32483f
C50158 _0527_/a_109_47# net154 0
C50159 _1072_/a_27_47# _1072_/a_1059_315# 0.04875f
C50160 _1072_/a_193_47# _1072_/a_466_413# 0.08301f
C50161 _0841_/a_79_21# _0841_/a_215_47# 0.04584f
C50162 _0684_/a_59_75# clkbuf_0__0462_/a_110_47# 0.00568f
C50163 _0100_ _0217_ 0.02381f
C50164 _0328_ _0327_ 0.04485f
C50165 VPWR _1019_/a_381_47# 0.07064f
C50166 _0714_/a_245_297# VPWR 0.00471f
C50167 _0765_/a_215_47# _0181_ 0
C50168 hold88/a_285_47# _0088_ 0
C50169 _0640_/a_109_53# _0346_ 0
C50170 net101 _0585_/a_27_297# 0
C50171 _0314_ _0732_/a_80_21# 0
C50172 _0532_/a_299_297# clknet_1_1__leaf__0457_ 0
C50173 _0241_ acc0.A\[18\] 0
C50174 acc0.A\[14\] _0996_/a_975_413# 0.00112f
C50175 comp0.B\[3\] net27 0
C50176 _0218_ _0300_ 0.02204f
C50177 _0343_ hold72/a_391_47# 0
C50178 _1067_/a_891_413# _1067_/a_975_413# 0.00851f
C50179 _1067_/a_381_47# _1067_/a_561_413# 0.00123f
C50180 _0251_ net65 0.55766f
C50181 hold36/a_49_47# hold37/a_391_47# 0
C50182 _0251_ _0989_/a_466_413# 0.00223f
C50183 _0429_ _0989_/a_193_47# 0
C50184 _1001_/a_381_47# _0345_ 0.00445f
C50185 hold31/a_285_47# hold31/a_391_47# 0.41909f
C50186 clkbuf_1_0__f__0457_/a_110_47# control0.add 0.11503f
C50187 _0341_ _0999_/a_1059_315# 0
C50188 _1071_/a_1059_315# _0169_ 0
C50189 _1050_/a_1059_315# _0172_ 0
C50190 hold90/a_49_47# _0219_ 0.00755f
C50191 acc0.A\[17\] hold72/a_285_47# 0.00107f
C50192 _1004_/a_27_47# _0350_ 0.00261f
C50193 _0343_ hold87/a_391_47# 0
C50194 _0252_ _0989_/a_381_47# 0.01494f
C50195 net65 _0989_/a_592_47# 0
C50196 _0989_/a_466_413# _0989_/a_592_47# 0.00553f
C50197 _0989_/a_634_159# _0989_/a_1017_47# 0
C50198 _0997_/a_27_47# _0997_/a_1059_315# 0.04861f
C50199 _0997_/a_193_47# _0997_/a_466_413# 0.07482f
C50200 _1020_/a_466_413# clknet_1_0__leaf__0461_ 0
C50201 _0126_ _0350_ 0
C50202 _0129_ hold92/a_391_47# 0
C50203 _0181_ _0986_/a_1059_315# 0.00431f
C50204 _0544_/a_51_297# _1042_/a_891_413# 0.00142f
C50205 _0544_/a_240_47# _1042_/a_193_47# 0
C50206 pp[2] VPWR 0.4538f
C50207 hold30/a_49_47# pp[19] 0
C50208 _0121_ output46/a_27_47# 0
C50209 hold30/a_391_47# net46 0.00695f
C50210 _0438_ clkbuf_1_1__f__0458_/a_110_47# 0.19803f
C50211 acc0.A\[16\] _0583_/a_109_47# 0
C50212 _0992_/a_466_413# _0992_/a_592_47# 0.00553f
C50213 _0992_/a_634_159# _0992_/a_1017_47# 0
C50214 _0749_/a_384_47# _0369_ 0
C50215 comp0.B\[4\] net121 0
C50216 VPWR _1051_/a_634_159# 0.18599f
C50217 net58 _0346_ 0.02918f
C50218 net78 hold81/a_49_47# 0
C50219 _0349_ _0704_/a_68_297# 0
C50220 _0718_/a_285_47# acc0.A\[30\] 0
C50221 _0263_ _0843_/a_150_297# 0
C50222 net111 acc0.A\[25\] 0.05845f
C50223 hold6/a_49_47# _1042_/a_27_47# 0
C50224 VPWR _1045_/a_1059_315# 0.39949f
C50225 _0402_ _0808_/a_266_47# 0.00141f
C50226 _0349_ pp[27] 0.00981f
C50227 _0125_ _1027_/a_1017_47# 0
C50228 _0371_ _0693_/a_68_297# 0
C50229 clknet_0__0458_ _0841_/a_297_297# 0
C50230 _0134_ _0211_ 0.11711f
C50231 _0959_/a_300_47# _0474_ 0
C50232 hold13/a_285_47# comp0.B\[6\] 0.01526f
C50233 hold13/a_391_47# comp0.B\[5\] 0.06756f
C50234 net58 net65 0
C50235 _1027_/a_27_47# _1027_/a_193_47# 0.9705f
C50236 _0253_ _0830_/a_79_21# 0
C50237 hold46/a_49_47# hold26/a_285_47# 0.00402f
C50238 _1061_/a_634_159# _1061_/a_381_47# 0
C50239 hold54/a_49_47# net201 0
C50240 A[13] _0297_ 0
C50241 net51 _0754_/a_512_297# 0
C50242 _0291_ _0990_/a_193_47# 0
C50243 net66 _0990_/a_466_413# 0.01181f
C50244 acc0.A\[8\] _0990_/a_634_159# 0.00866f
C50245 net221 _0219_ 0
C50246 _0581_/a_27_297# _0612_/a_59_75# 0.01028f
C50247 _0225_ _0757_/a_68_297# 0
C50248 _0629_/a_145_75# _0465_ 0
C50249 _0216_ _1026_/a_1017_47# 0.00156f
C50250 _1054_/a_193_47# A[4] 0
C50251 _1007_/a_381_47# _0219_ 0
C50252 _0984_/a_27_47# net165 0
C50253 _0363_ _0362_ 0.07915f
C50254 _0319_ _0360_ 0.14551f
C50255 _0361_ _0731_/a_81_21# 0
C50256 clkbuf_0__0459_/a_110_47# acc0.A\[13\] 0.0347f
C50257 _0313_ net197 0
C50258 clkload0/X net35 0.02813f
C50259 _0216_ _0122_ 0.00738f
C50260 _0180_ hold83/a_391_47# 0.02874f
C50261 _0399_ _0833_/a_79_21# 0.17099f
C50262 _1035_/a_27_47# _1035_/a_466_413# 0.27314f
C50263 _1035_/a_193_47# _1035_/a_634_159# 0.11486f
C50264 pp[18] _0714_/a_512_297# 0
C50265 _0734_/a_47_47# _0219_ 0.01735f
C50266 net24 control0.reset 0
C50267 _0629_/a_59_75# net58 0.18158f
C50268 _0279_ _0297_ 0.00256f
C50269 _0959_/a_80_21# _1065_/a_193_47# 0
C50270 _0959_/a_217_297# _1065_/a_27_47# 0
C50271 _0559_/a_240_47# net25 0
C50272 _0217_ _1014_/a_975_413# 0
C50273 _0787_/a_209_47# _0091_ 0
C50274 _0489_ _1069_/a_466_413# 0.02105f
C50275 hold15/a_285_47# _0338_ 0
C50276 _1065_/a_381_47# clknet_1_0__leaf__0457_ 0
C50277 _0182_ _0197_ 0
C50278 _0661_/a_27_297# _0401_ 0
C50279 hold89/a_285_47# _0166_ 0
C50280 clknet_1_1__leaf__0462_ _0320_ 0.00149f
C50281 comp0.B\[1\] _0175_ 0
C50282 net140 input12/a_75_212# 0.00241f
C50283 _0402_ _0345_ 0.13739f
C50284 net76 _0990_/a_1059_315# 0
C50285 _0404_ _0218_ 0.0819f
C50286 clknet_1_0__leaf__0459_ _1016_/a_27_47# 0.03076f
C50287 VPWR _1028_/a_1017_47# 0
C50288 _1069_/a_27_47# _0167_ 0.10264f
C50289 _1069_/a_193_47# clknet_1_0__leaf_clk 0.03132f
C50290 _1069_/a_1059_315# _1069_/a_1017_47# 0
C50291 VPWR _0761_/a_113_47# 0
C50292 _1056_/a_466_413# net66 0
C50293 output44/a_27_47# net209 0
C50294 _0854_/a_297_297# _0181_ 0
C50295 net117 _1030_/a_193_47# 0
C50296 _0552_/a_150_297# _0176_ 0.00123f
C50297 clknet_0__0465_ _0990_/a_891_413# 0.01431f
C50298 _1059_/a_381_47# acc0.A\[13\] 0
C50299 _1059_/a_466_413# net5 0
C50300 _1059_/a_193_47# _0185_ 0.03415f
C50301 VPWR _0534_/a_81_21# 0.20574f
C50302 pp[8] _1055_/a_193_47# 0
C50303 _0555_/a_149_47# net29 0
C50304 _0343_ _0600_/a_337_297# 0.00172f
C50305 _0233_ _0600_/a_103_199# 0.17191f
C50306 _0460_ net52 0.24963f
C50307 VPWR hold62/a_49_47# 0.27237f
C50308 net84 _0352_ 0
C50309 _1041_/a_891_413# _1040_/a_466_413# 0
C50310 _1031_/a_975_413# _0220_ 0.00138f
C50311 comp0.B\[5\] _0160_ 0
C50312 net194 _0464_ 0.00294f
C50313 net211 _0241_ 0
C50314 clknet_1_0__leaf__0465_ VPWR 3.9918f
C50315 _0624_/a_145_75# net62 0.00298f
C50316 _0482_ _0168_ 0.00108f
C50317 hold23/a_391_47# VPWR 0.18357f
C50318 _0577_/a_27_297# _0577_/a_109_47# 0.00393f
C50319 _0433_ acc0.A\[8\] 0
C50320 _1027_/a_27_47# _1026_/a_1059_315# 0.00174f
C50321 _0399_ _0158_ 0
C50322 _0083_ _0350_ 0.00117f
C50323 _0211_ _0554_/a_68_297# 0
C50324 _1039_/a_891_413# net171 0
C50325 hold26/a_285_47# comp0.B\[14\] 0.0016f
C50326 _0361_ acc0.A\[25\] 0
C50327 net104 _0350_ 0
C50328 _0137_ comp0.B\[8\] 0
C50329 _0959_/a_80_21# net33 0.11884f
C50330 _0343_ _1011_/a_1059_315# 0.00323f
C50331 _0680_/a_80_21# _0310_ 0
C50332 _0217_ _1022_/a_1059_315# 0
C50333 _0120_ _1022_/a_27_47# 0
C50334 acc0.A\[22\] _1022_/a_466_413# 0.00125f
C50335 _0260_ _0445_ 0
C50336 clknet_1_1__leaf__0458_ _0989_/a_193_47# 0
C50337 hold57/a_285_47# net160 0.00114f
C50338 hold1/a_285_47# clknet_1_1__leaf__0458_ 0.01355f
C50339 _0123_ net50 0
C50340 _0538_/a_149_47# net183 0.01209f
C50341 hold75/a_285_47# _0451_ 0
C50342 net235 acc0.A\[6\] 0
C50343 _0561_/a_149_47# hold84/a_49_47# 0
C50344 _0545_/a_68_297# net127 0
C50345 _0474_ _0208_ 0.45047f
C50346 comp0.B\[6\] _0132_ 0.01079f
C50347 _0524_/a_27_297# _0524_/a_373_47# 0.01338f
C50348 _1022_/a_381_47# net151 0.14282f
C50349 output38/a_27_47# _0993_/a_27_47# 0
C50350 _0646_/a_285_47# _0218_ 0
C50351 output53/a_27_47# net210 0
C50352 hold22/a_285_47# _0191_ 0.09948f
C50353 _0430_ _0990_/a_27_47# 0
C50354 clknet_1_0__leaf__0459_ _1019_/a_381_47# 0.00327f
C50355 _1003_/a_27_47# _0974_/a_448_47# 0
C50356 _1003_/a_193_47# _0974_/a_544_297# 0
C50357 hold12/a_391_47# net159 0.13083f
C50358 net99 pp[31] 0
C50359 _0994_/a_891_413# _0994_/a_975_413# 0.00851f
C50360 _0994_/a_381_47# _0994_/a_561_413# 0.00123f
C50361 _0550_/a_51_297# input30/a_75_212# 0
C50362 net36 _0173_ 0
C50363 _1020_/a_592_47# clknet_1_0__leaf__0457_ 0
C50364 _0285_ _0419_ 0.03534f
C50365 _0779_/a_215_47# _0097_ 0.00187f
C50366 _1056_/a_466_413# _0350_ 0
C50367 _1055_/a_1017_47# net179 0
C50368 _0500_/a_27_47# _1048_/a_193_47# 0.00182f
C50369 _0733_/a_79_199# acc0.A\[27\] 0
C50370 _0972_/a_93_21# _0972_/a_250_297# 0.18824f
C50371 _0260_ _0643_/a_253_47# 0.01102f
C50372 net203 _0564_/a_68_297# 0
C50373 hold56/a_49_47# _0215_ 0
C50374 _1023_/a_381_47# net51 0.00987f
C50375 _0720_/a_68_297# clknet_1_1__leaf__0462_ 0.05908f
C50376 _0349_ _0216_ 0.02002f
C50377 _0835_/a_215_47# _0256_ 0.0214f
C50378 _0401_ _0990_/a_27_47# 0
C50379 hold14/a_391_47# net161 0.13105f
C50380 _0466_ _0161_ 0
C50381 _1003_/a_975_413# _0101_ 0
C50382 net36 _1047_/a_1017_47# 0.00125f
C50383 comp0.B\[11\] _0202_ 0.03021f
C50384 _0503_/a_109_297# _0180_ 0.00351f
C50385 _0993_/a_27_47# _0993_/a_1059_315# 0.04875f
C50386 _0993_/a_193_47# _0993_/a_466_413# 0.08301f
C50387 _1058_/a_193_47# _0156_ 0.18448f
C50388 _0369_ acc0.A\[10\] 0.0462f
C50389 clknet_0__0463_ _0498_/a_240_47# 0
C50390 _0235_ _0385_ 0
C50391 _1039_/a_634_159# _1039_/a_381_47# 0
C50392 _0186_ _0826_/a_27_53# 0
C50393 net203 clknet_1_1__leaf_clk 0
C50394 hold33/a_49_47# _0138_ 0.01746f
C50395 _0274_ _0369_ 0.02565f
C50396 _1020_/a_561_413# _0457_ 0
C50397 _0578_/a_109_297# net1 0.00663f
C50398 _0280_ _0672_/a_297_297# 0.00465f
C50399 acc0.A\[27\] net244 0.04109f
C50400 A[12] _0512_/a_109_47# 0.00104f
C50401 _0996_/a_27_47# _0405_ 0
C50402 _0172_ _1046_/a_891_413# 0.00153f
C50403 _1032_/a_27_47# _0215_ 0
C50404 hold14/a_391_47# net26 0.00214f
C50405 net55 _0735_/a_109_297# 0
C50406 _1049_/a_193_47# _0148_ 0
C50407 acc0.A\[14\] _0399_ 0.22886f
C50408 _1026_/a_193_47# _1026_/a_381_47# 0.09984f
C50409 _1026_/a_634_159# _1026_/a_891_413# 0.03684f
C50410 _1026_/a_27_47# _1026_/a_561_413# 0.0027f
C50411 _0733_/a_544_297# _0321_ 0.00149f
C50412 _0733_/a_448_47# _0360_ 0.08496f
C50413 _0985_/a_891_413# clknet_1_0__leaf__0458_ 0
C50414 hold10/a_391_47# _1047_/a_27_47# 0
C50415 _0234_ _1005_/a_891_413# 0.00527f
C50416 _0343_ _0341_ 0.03326f
C50417 net169 _1053_/a_561_413# 0
C50418 net140 _1053_/a_975_413# 0
C50419 _0714_/a_240_47# _0567_/a_27_297# 0
C50420 net64 _0433_ 0.00319f
C50421 _0407_ net41 0.22644f
C50422 _0195_ _0583_/a_27_297# 0
C50423 VPWR _0400_ 0.38544f
C50424 _1024_/a_634_159# net110 0
C50425 hold97/a_285_47# clkbuf_1_1__f__0460_/a_110_47# 0
C50426 _0217_ _1067_/a_381_47# 0
C50427 _0183_ _1067_/a_1059_315# 0
C50428 _1024_/a_891_413# _1024_/a_1017_47# 0.00617f
C50429 _1024_/a_193_47# _0122_ 0.22917f
C50430 _0854_/a_79_21# _1018_/a_193_47# 0
C50431 net1 net202 0
C50432 _0227_ _0605_/a_109_297# 0
C50433 _0337_ _0335_ 0
C50434 input32/a_75_212# net128 0.02251f
C50435 net1 clknet_1_1__leaf__0463_ 0
C50436 _1014_/a_634_159# _0181_ 0
C50437 _0121_ hold29/a_391_47# 0
C50438 _0278_ _0646_/a_47_47# 0.14425f
C50439 _1036_/a_466_413# net25 0
C50440 _1057_/a_27_47# net143 0.23602f
C50441 net33 _0173_ 0
C50442 output43/a_27_47# _0997_/a_1059_315# 0
C50443 _0098_ _0388_ 0
C50444 _0369_ pp[5] 0
C50445 _0540_/a_240_47# net20 0.06463f
C50446 _0540_/a_245_297# _0142_ 0
C50447 clk _1064_/a_1017_47# 0
C50448 net243 acc0.A\[22\] 0
C50449 _1048_/a_381_47# net134 0.00201f
C50450 hold78/a_285_47# _0220_ 0.01396f
C50451 net168 net65 0
C50452 _0831_/a_117_297# _0434_ 0.01089f
C50453 net242 _0720_/a_68_297# 0
C50454 _0195_ _0999_/a_193_47# 0
C50455 _1020_/a_193_47# _0208_ 0.00654f
C50456 _1068_/a_891_413# _0468_ 0.04653f
C50457 _1041_/a_27_47# _1041_/a_466_413# 0.26005f
C50458 _1041_/a_193_47# _1041_/a_634_159# 0.12497f
C50459 _0343_ _1013_/a_891_413# 0.02013f
C50460 net176 _0352_ 0
C50461 _0624_/a_59_75# _0270_ 0.01085f
C50462 hold99/a_49_47# _0993_/a_193_47# 0
C50463 hold99/a_285_47# _0993_/a_27_47# 0
C50464 B[15] B[1] 0.10313f
C50465 _0254_ _0434_ 0.00216f
C50466 _1017_/a_27_47# _0219_ 0
C50467 clknet_0__0457_ _0117_ 0
C50468 _0172_ _0256_ 0
C50469 net43 _0240_ 0
C50470 VPWR _0773_/a_117_297# 0.00986f
C50471 hold69/a_285_47# _0352_ 0
C50472 _1015_/a_1059_315# comp0.B\[15\] 0.08402f
C50473 _0369_ net43 0.00213f
C50474 _0172_ _0987_/a_1059_315# 0
C50475 net63 _0255_ 0.48579f
C50476 net76 _0439_ 0.01649f
C50477 _0302_ acc0.A\[15\] 0.31905f
C50478 _1002_/a_27_47# net1 0.00353f
C50479 _0232_ _0249_ 0.07001f
C50480 _0248_ _0771_/a_382_47# 0
C50481 hold76/a_391_47# _1001_/a_27_47# 0
C50482 _0855_/a_299_297# acc0.A\[1\] 0
C50483 input12/a_75_212# input14/a_75_212# 0
C50484 net76 VPWR 0.36298f
C50485 clknet_0__0457_ hold73/a_285_47# 0
C50486 net152 _0140_ 0.23582f
C50487 hold2/a_285_47# net149 0.0114f
C50488 clknet_0__0464_ _1061_/a_634_159# 0
C50489 _0129_ _0336_ 0.03157f
C50490 clkbuf_1_0__f__0460_/a_110_47# _1006_/a_381_47# 0
C50491 _0616_/a_78_199# _0242_ 0.00963f
C50492 net116 clknet_1_1__leaf__0462_ 0.18303f
C50493 _0130_ _0113_ 0
C50494 _1053_/a_381_47# net13 0
C50495 _1053_/a_592_47# acc0.A\[6\] 0
C50496 clknet_1_0__leaf__0465_ _1054_/a_1017_47# 0
C50497 hold44/a_391_47# _1029_/a_27_47# 0
C50498 hold44/a_49_47# _1029_/a_634_159# 0
C50499 hold44/a_285_47# _1029_/a_193_47# 0
C50500 net226 _0466_ 0.29139f
C50501 clknet_0__0458_ _0627_/a_109_93# 0.00594f
C50502 hold85/a_49_47# hold84/a_391_47# 0
C50503 hold85/a_391_47# hold84/a_49_47# 0.00139f
C50504 hold85/a_285_47# hold84/a_285_47# 0
C50505 net164 _0169_ 0.30224f
C50506 _0752_/a_27_413# _0762_/a_79_21# 0
C50507 _0267_ _0843_/a_68_297# 0
C50508 _1072_/a_891_413# _1072_/a_1017_47# 0.00617f
C50509 _0087_ _0186_ 0.02875f
C50510 _0841_/a_510_47# _0084_ 0
C50511 _0183_ net6 0.01032f
C50512 _0317_ _0321_ 0.04601f
C50513 net101 _0112_ 0
C50514 clknet_1_0__leaf__0461_ hold60/a_285_47# 0.01715f
C50515 net65 _0831_/a_285_297# 0
C50516 _0554_/a_68_297# _0210_ 0.106f
C50517 hold68/a_49_47# _0352_ 0
C50518 _1013_/a_1059_315# net60 0.09744f
C50519 _0081_ _0583_/a_27_297# 0
C50520 _1037_/a_891_413# net171 0
C50521 _1037_/a_1059_315# _0207_ 0.00244f
C50522 _0471_ _1062_/a_466_413# 0.00234f
C50523 VPWR _1025_/a_381_47# 0.076f
C50524 _0661_/a_27_297# _0089_ 0
C50525 _0244_ net104 0
C50526 clknet_1_1__leaf__0462_ hold92/a_285_47# 0.00927f
C50527 _0183_ _0447_ 0
C50528 clknet_1_1__leaf__0460_ net97 0.13965f
C50529 net183 clkbuf_0__0464_/a_110_47# 0.01317f
C50530 _0216_ _0181_ 0.55139f
C50531 _0428_ net47 0.03228f
C50532 _0476_ _0559_/a_149_47# 0.00108f
C50533 net181 _0186_ 0
C50534 _0800_/a_51_297# pp[14] 0
C50535 _0643_/a_103_199# _0445_ 0
C50536 net210 net111 0.07089f
C50537 _0190_ _0833_/a_79_21# 0
C50538 _0195_ _0570_/a_27_297# 0.11912f
C50539 _0997_/a_891_413# _0997_/a_1017_47# 0.00617f
C50540 _1053_/a_466_413# _0150_ 0
C50541 _0118_ clknet_1_0__leaf__0461_ 0
C50542 _1037_/a_891_413# net24 0
C50543 _0460_ hold93/a_49_47# 0.10545f
C50544 clknet_1_0__leaf__0457_ hold93/a_391_47# 0.00257f
C50545 _0140_ _1042_/a_466_413# 0.02129f
C50546 net198 _1042_/a_561_413# 0
C50547 VPWR _1044_/a_466_413# 0.24776f
C50548 clknet_1_0__leaf__0464_ _0527_/a_109_297# 0
C50549 VPWR net137 0.39696f
C50550 _0159_ acc0.A\[15\] 0
C50551 acc0.A\[29\] _0347_ 0
C50552 _0732_/a_80_21# _0360_ 0.0777f
C50553 clknet_0__0459_ _1059_/a_193_47# 0
C50554 net26 _0132_ 0
C50555 hold88/a_391_47# _0399_ 0.01128f
C50556 _0783_/a_510_47# _0352_ 0
C50557 _0982_/a_1059_315# _0345_ 0.02624f
C50558 _0218_ _0419_ 0.03789f
C50559 _0109_ net191 0
C50560 _0243_ _0773_/a_285_297# 0
C50561 _0316_ _0699_/a_68_297# 0
C50562 _1001_/a_466_413# _0461_ 0.00556f
C50563 net243 _0379_ 0.00485f
C50564 clkbuf_1_1__f__0465_/a_110_47# _0812_/a_215_47# 0
C50565 _0786_/a_80_21# _0421_ 0
C50566 _1035_/a_27_47# _0561_/a_51_297# 0
C50567 _1027_/a_466_413# _1027_/a_592_47# 0.00553f
C50568 _1027_/a_634_159# _1027_/a_1017_47# 0
C50569 _0643_/a_103_199# _0643_/a_253_47# 0.06061f
C50570 net44 _0710_/a_109_297# 0.00442f
C50571 net237 _0105_ 0.00125f
C50572 _0181_ _1067_/a_27_47# 0
C50573 _0315_ _0367_ 0.1146f
C50574 hold8/a_49_47# clknet_1_1__leaf__0462_ 0.00447f
C50575 VPWR _0849_/a_510_47# 0.00108f
C50576 acc0.A\[15\] net6 0.19246f
C50577 acc0.A\[16\] _0998_/a_27_47# 0
C50578 _0291_ clknet_1_1__leaf__0465_ 0.04655f
C50579 VPWR _1032_/a_975_413# 0.0049f
C50580 _1061_/a_381_47# net147 0
C50581 net205 clkbuf_1_1__f__0463_/a_110_47# 0
C50582 _0699_/a_68_297# _0347_ 0.00211f
C50583 _0462_ _0745_/a_193_47# 0
C50584 clknet_1_0__leaf__0462_ _1023_/a_193_47# 0.00475f
C50585 _0555_/a_149_47# comp0.B\[6\] 0
C50586 _0555_/a_240_47# comp0.B\[5\] 0.00121f
C50587 net66 _0088_ 0.56676f
C50588 net219 acc0.A\[18\] 0.0438f
C50589 _0116_ _0612_/a_59_75# 0.00106f
C50590 hold10/a_391_47# net133 0
C50591 _0195_ hold50/a_49_47# 0
C50592 clknet_1_0__leaf__0464_ _1061_/a_193_47# 0
C50593 _0715_/a_27_47# net47 0.01797f
C50594 net166 clknet_1_1__leaf__0465_ 0
C50595 net126 net172 0
C50596 _0340_ _1030_/a_891_413# 0
C50597 _0447_ acc0.A\[15\] 0.00344f
C50598 hold29/a_391_47# _0380_ 0
C50599 A[1] B[6] 0.00343f
C50600 _1065_/a_634_159# _0161_ 0.00133f
C50601 net232 net33 0.07678f
C50602 _1035_/a_27_47# _0133_ 0.09793f
C50603 _1035_/a_193_47# net121 0.00703f
C50604 _1035_/a_1059_315# _1035_/a_1017_47# 0
C50605 _0668_/a_382_297# _0668_/a_297_47# 0
C50606 _0250_ _0360_ 0.00124f
C50607 pp[18] _0111_ 0
C50608 _0357_ _0729_/a_68_297# 0
C50609 _0243_ _0350_ 0.08032f
C50610 hold39/a_49_47# _1034_/a_193_47# 0
C50611 hold39/a_285_47# _1034_/a_27_47# 0.01125f
C50612 net238 _0219_ 0
C50613 _0477_ comp0.B\[6\] 0
C50614 _0312_ _0747_/a_79_21# 0
C50615 _1051_/a_193_47# _0172_ 0.2396f
C50616 _0183_ acc0.A\[0\] 0.01314f
C50617 _0977_/a_75_212# control0.count\[0\] 0.00105f
C50618 _0489_ _0167_ 0.04303f
C50619 net172 input8/a_75_212# 0
C50620 control0.reset clknet_1_0__leaf__0457_ 0.00174f
C50621 _0410_ _0669_/a_29_53# 0
C50622 _0725_/a_80_21# _0723_/a_207_413# 0.00121f
C50623 _0172_ _1045_/a_466_413# 0.02179f
C50624 VPWR _0533_/a_373_47# 0
C50625 _0293_ _0401_ 0.10258f
C50626 _0287_ _0425_ 0
C50627 _0558_/a_68_297# _1035_/a_27_47# 0
C50628 hold69/a_391_47# _0326_ 0
C50629 _0151_ _0150_ 0
C50630 _0446_ _0219_ 0.15783f
C50631 _0451_ _0345_ 0
C50632 VPWR hold71/a_391_47# 0.18886f
C50633 clknet_1_1__leaf__0459_ _1013_/a_466_413# 0
C50634 _0399_ _0823_/a_109_297# 0
C50635 _0460_ hold94/a_391_47# 0
C50636 _0496_/a_27_47# _0175_ 0.22537f
C50637 VPWR _0546_/a_240_47# 0.00313f
C50638 acc0.A\[29\] _1029_/a_1017_47# 0
C50639 net44 _0607_/a_27_297# 0.17091f
C50640 _1011_/a_634_159# _0726_/a_240_47# 0
C50641 _1011_/a_466_413# _0726_/a_149_47# 0
C50642 _0343_ hold91/a_49_47# 0.00228f
C50643 _1069_/a_975_413# control0.count\[0\] 0.00107f
C50644 clknet_1_0__leaf__0465_ _0523_/a_81_21# 0.00718f
C50645 _1033_/a_193_47# _1065_/a_1059_315# 0
C50646 net32 _1043_/a_193_47# 0
C50647 _0993_/a_27_47# acc0.A\[10\] 0
C50648 _1052_/a_27_47# net148 0
C50649 acc0.A\[31\] pp[31] 0.01201f
C50650 hold78/a_391_47# _0218_ 0.00147f
C50651 _0160_ hold84/a_49_47# 0
C50652 _0231_ _0232_ 0.05461f
C50653 _0181_ net247 0.1292f
C50654 _1041_/a_891_413# net174 0
C50655 net56 _0727_/a_109_47# 0
C50656 net125 _0465_ 0.00144f
C50657 net125 _1061_/a_381_47# 0.0043f
C50658 _0734_/a_377_297# _0318_ 0.00141f
C50659 _0399_ _1016_/a_634_159# 0
C50660 _0088_ _0350_ 0
C50661 _0488_ _0162_ 0
C50662 net150 _0217_ 0.2369f
C50663 _0195_ _1018_/a_634_159# 0.01145f
C50664 net156 _1026_/a_193_47# 0
C50665 net58 _0988_/a_634_159# 0.00277f
C50666 _0640_/a_465_297# clknet_1_1__leaf__0458_ 0
C50667 _0179_ net6 0
C50668 _0467_ _1067_/a_466_413# 0
C50669 _0300_ _0792_/a_80_21# 0
C50670 _0794_/a_27_47# _0405_ 0
C50671 net208 hold62/a_285_47# 0.06144f
C50672 _0195_ _1049_/a_27_47# 0
C50673 hold15/a_285_47# acc0.A\[31\] 0.01043f
C50674 _0990_/a_193_47# _0986_/a_1059_315# 0
C50675 _0645_/a_129_47# _0302_ 0
C50676 acc0.A\[22\] net151 0.04288f
C50677 acc0.A\[27\] clkbuf_1_1__f__0462_/a_110_47# 0.02114f
C50678 _0563_/a_149_47# _0173_ 0.02257f
C50679 _0563_/a_51_297# _0208_ 0.23586f
C50680 _0132_ hold84/a_285_47# 0
C50681 net21 _0143_ 0
C50682 hold58/a_391_47# _1034_/a_193_47# 0
C50683 acc0.A\[21\] _0219_ 0.02696f
C50684 _0227_ net241 0.06193f
C50685 A[4] acc0.A\[6\] 0
C50686 _0179_ _0447_ 0.0256f
C50687 _0524_/a_373_47# _0194_ 0
C50688 acc0.A\[0\] acc0.A\[15\] 0
C50689 net9 _0528_/a_384_47# 0
C50690 _0635_/a_109_297# _0465_ 0
C50691 _1065_/a_381_47# _0160_ 0
C50692 net163 _0218_ 0
C50693 net58 _0259_ 0.03887f
C50694 _0472_ _0214_ 0
C50695 net89 _0974_/a_222_93# 0
C50696 _0101_ _0974_/a_79_199# 0
C50697 net211 _1019_/a_466_413# 0
C50698 net199 acc0.A\[25\] 0.00232f
C50699 _0995_/a_1059_315# output41/a_27_47# 0
C50700 _0995_/a_193_47# net41 0
C50701 _0800_/a_149_47# _0400_ 0
C50702 _0183_ _0580_/a_109_297# 0.00919f
C50703 _0172_ input30/a_75_212# 0
C50704 _0520_/a_27_297# net168 0.05729f
C50705 _0290_ clknet_1_1__leaf__0465_ 0.18093f
C50706 net61 _0830_/a_79_21# 0.00259f
C50707 net45 _1013_/a_561_413# 0
C50708 comp0.B\[7\] clknet_1_0__leaf__0463_ 0.05428f
C50709 _1018_/a_1059_315# _0247_ 0
C50710 VPWR clkbuf_0__0459_/a_110_47# 1.28643f
C50711 hold35/a_285_47# net66 0
C50712 _0179_ _1048_/a_561_413# 0
C50713 _0972_/a_250_297# net231 0.041f
C50714 _0972_/a_93_21# _0164_ 0.10672f
C50715 _0220_ hold61/a_391_47# 0.03141f
C50716 _0336_ hold61/a_285_47# 0.00416f
C50717 acc0.A\[23\] net51 0.67221f
C50718 _0538_/a_245_297# comp0.B\[10\] 0
C50719 _1043_/a_193_47# _1042_/a_1059_315# 0.00113f
C50720 _1043_/a_27_47# _1042_/a_891_413# 0
C50721 _1043_/a_466_413# _1042_/a_634_159# 0
C50722 _1043_/a_634_159# _1042_/a_466_413# 0
C50723 _1043_/a_891_413# _1042_/a_27_47# 0
C50724 _1043_/a_1059_315# _1042_/a_193_47# 0.00113f
C50725 _0464_ net132 0.09826f
C50726 net116 hold92/a_49_47# 0
C50727 net141 _0988_/a_1059_315# 0
C50728 net147 net174 0.00173f
C50729 clkbuf_0__0461_/a_110_47# hold72/a_391_47# 0.01029f
C50730 _1030_/a_193_47# _0704_/a_68_297# 0
C50731 _0182_ _0566_/a_27_47# 0.22207f
C50732 _0642_/a_27_413# _0989_/a_193_47# 0
C50733 _0642_/a_215_297# _0989_/a_27_47# 0
C50734 _0993_/a_891_413# _0993_/a_1017_47# 0.00617f
C50735 pp[27] _1030_/a_193_47# 0.00137f
C50736 _0373_ _0345_ 0.00141f
C50737 clkbuf_1_1__f__0465_/a_110_47# _0659_/a_68_297# 0.00201f
C50738 _0627_/a_215_53# _0627_/a_297_297# 0.00494f
C50739 hold85/a_391_47# _0471_ 0
C50740 _1039_/a_891_413# _0553_/a_51_297# 0.00728f
C50741 pp[6] acc0.A\[6\] 0
C50742 _1039_/a_381_47# net125 0
C50743 _0742_/a_299_297# _0315_ 0.07171f
C50744 _0180_ net9 0.84012f
C50745 _0199_ net175 0
C50746 _0730_/a_297_297# _0730_/a_215_47# 0
C50747 _0730_/a_79_21# _0730_/a_510_47# 0.00844f
C50748 _0751_/a_29_53# net46 0.01873f
C50749 _0535_/a_68_297# _1040_/a_891_413# 0
C50750 clknet_1_1__leaf__0460_ _1010_/a_27_47# 0.0612f
C50751 acc0.A\[29\] hold95/a_49_47# 0.01481f
C50752 _0343_ _0707_/a_208_47# 0
C50753 net10 _1043_/a_193_47# 0.0095f
C50754 _0714_/a_51_297# _1031_/a_466_413# 0
C50755 _0714_/a_149_47# _1031_/a_27_47# 0
C50756 _0399_ _0116_ 0
C50757 hold92/a_49_47# hold92/a_285_47# 0.22264f
C50758 net63 _0830_/a_215_47# 0.00747f
C50759 _0147_ net170 0
C50760 _0485_ _1064_/a_466_413# 0.00149f
C50761 _0487_ _1064_/a_634_159# 0
C50762 clknet_0__0462_ _0318_ 0.28462f
C50763 _0162_ _1064_/a_27_47# 0.0998f
C50764 _0366_ _0379_ 0
C50765 _0747_/a_297_297# _0219_ 0
C50766 _0549_/a_68_297# _0208_ 0
C50767 _1026_/a_891_413# net112 0
C50768 _1026_/a_193_47# acc0.A\[26\] 0
C50769 _1059_/a_381_47# VPWR 0.07606f
C50770 control0.count\[3\] _1005_/a_27_47# 0
C50771 _0465_ _1047_/a_1059_315# 0.01096f
C50772 _0097_ net42 0
C50773 _0473_ _0465_ 0
C50774 _1072_/a_466_413# control0.state\[2\] 0
C50775 _0375_ _0103_ 0.02342f
C50776 _0216_ _1012_/a_193_47# 0
C50777 _0472_ _1061_/a_1059_315# 0
C50778 hold25/a_49_47# _0552_/a_68_297# 0
C50779 hold14/a_49_47# _1035_/a_27_47# 0
C50780 _0817_/a_81_21# _0817_/a_585_47# 0.00695f
C50781 _0817_/a_266_297# _0817_/a_266_47# 0
C50782 acc0.A\[19\] _0771_/a_27_413# 0.01335f
C50783 clknet_1_1__leaf__0460_ _1009_/a_193_47# 0.046f
C50784 _0181_ _1009_/a_975_413# 0
C50785 _0352_ acc0.A\[18\] 0
C50786 clknet_1_1__leaf__0458_ _0988_/a_27_47# 0.0078f
C50787 _0323_ _0359_ 0.20898f
C50788 acc0.A\[2\] _1047_/a_1059_315# 0
C50789 _0081_ _1018_/a_634_159# 0
C50790 _0217_ control0.add 0.92636f
C50791 _1024_/a_592_47# acc0.A\[24\] 0
C50792 _0542_/a_512_297# net20 0
C50793 _0171_ _0560_/a_68_297# 0
C50794 clknet_1_1__leaf__0463_ control0.sh 0.03431f
C50795 net54 _0571_/a_109_297# 0
C50796 _0271_ _0345_ 0
C50797 _0121_ net50 0
C50798 _0670_/a_79_21# net5 0
C50799 hold66/a_285_47# net213 0.00853f
C50800 net100 _0181_ 0.06813f
C50801 net154 _0186_ 0.13419f
C50802 _0598_/a_297_47# _0219_ 0
C50803 _0789_/a_201_297# _0405_ 0.01314f
C50804 _0662_/a_299_297# _0259_ 0.06209f
C50805 _0343_ _0454_ 0
C50806 _0781_/a_68_297# clknet_1_1__leaf__0461_ 0
C50807 net38 net37 0
C50808 clkload2/a_110_47# VPWR 0
C50809 _0174_ _1040_/a_891_413# 0.00859f
C50810 _0136_ _1040_/a_27_47# 0
C50811 _1037_/a_634_159# _1037_/a_381_47# 0
C50812 _0602_/a_113_47# net51 0
C50813 _0218_ _0989_/a_193_47# 0
C50814 pp[16] _0997_/a_1017_47# 0
C50815 _0402_ _0992_/a_891_413# 0
C50816 acc0.A\[22\] _0378_ 0.00172f
C50817 _0255_ clkbuf_0__0465_/a_110_47# 0
C50818 _0835_/a_215_47# clknet_0__0465_ 0
C50819 _0475_ net24 0.39262f
C50820 _1029_/a_193_47# _0219_ 0
C50821 B[13] net196 0
C50822 net8 control0.sh 0
C50823 clknet_1_1__leaf__0459_ net67 0.0594f
C50824 clknet_1_0__leaf__0458_ net234 0.00118f
C50825 VPWR _1005_/a_466_413# 0.27906f
C50826 _0790_/a_285_297# acc0.A\[15\] 0.00749f
C50827 _0790_/a_285_47# net42 0.0022f
C50828 _0790_/a_35_297# _0406_ 0.17367f
C50829 _0731_/a_81_21# VPWR 0.23192f
C50830 VPWR _0519_/a_299_297# 0.28893f
C50831 _0343_ _0505_/a_27_297# 0
C50832 _0228_ hold3/a_285_47# 0.00618f
C50833 VPWR _0991_/a_1017_47# 0.00259f
C50834 net25 net26 0.0189f
C50835 _0465_ _0186_ 0
C50836 net54 _0737_/a_285_297# 0
C50837 clkbuf_1_1__f__0462_/a_110_47# _1010_/a_193_47# 0
C50838 _1054_/a_891_413# _0180_ 0.03186f
C50839 output65/a_27_47# VPWR 0.41078f
C50840 hold33/a_49_47# net22 0
C50841 _0220_ clknet_1_1__leaf__0462_ 0.00701f
C50842 hold30/a_285_47# _1023_/a_634_159# 0
C50843 hold30/a_391_47# _1023_/a_193_47# 0
C50844 _0243_ _0244_ 0.21819f
C50845 _0389_ _0386_ 0
C50846 hold64/a_285_47# _0181_ 0
C50847 pp[28] _1030_/a_27_47# 0
C50848 _1038_/a_466_413# net8 0
C50849 acc0.A\[2\] _0186_ 0.09694f
C50850 _1039_/a_381_47# _0473_ 0
C50851 hold9/a_49_47# _1008_/a_466_413# 0
C50852 _0608_/a_27_47# _0677_/a_47_47# 0
C50853 _0958_/a_109_47# _0471_ 0.00174f
C50854 clknet_0__0464_ net147 0
C50855 net61 _0219_ 0.03098f
C50856 _0216_ clknet_1_1__leaf__0461_ 0
C50857 _0335_ _0333_ 0.0664f
C50858 _0399_ _0422_ 0.0637f
C50859 _0198_ _0531_/a_27_297# 0.19321f
C50860 hold42/a_391_47# net3 0
C50861 _0869_/a_27_47# clknet_1_0__leaf__0457_ 0.20073f
C50862 _1049_/a_193_47# _1048_/a_27_47# 0.00327f
C50863 _1049_/a_27_47# _1048_/a_193_47# 0.00107f
C50864 net53 _1026_/a_634_159# 0
C50865 net189 _0512_/a_27_297# 0
C50866 _1057_/a_891_413# net3 0
C50867 clknet_1_0__leaf__0464_ clkbuf_0__0464_/a_110_47# 0.00309f
C50868 hold33/a_49_47# clknet_1_0__leaf__0463_ 0.00527f
C50869 acc0.A\[9\] acc0.A\[11\] 0.00143f
C50870 _0287_ hold70/a_285_47# 0
C50871 _0289_ hold70/a_391_47# 0
C50872 _0234_ _0369_ 0.02093f
C50873 VPWR _1011_/a_381_47# 0.07064f
C50874 hold97/a_285_47# net244 0.01067f
C50875 _0251_ _0253_ 0.12871f
C50876 input32/a_75_212# comp0.B\[11\] 0
C50877 hold88/a_391_47# _0190_ 0
C50878 VPWR _1006_/a_193_47# 0.33656f
C50879 _0476_ comp0.B\[5\] 0.00381f
C50880 _0452_ acc0.A\[1\] 0.21124f
C50881 _0751_/a_111_297# VPWR 0
C50882 net37 hold81/a_285_47# 0.02743f
C50883 _0963_/a_285_297# _1069_/a_891_413# 0
C50884 _1055_/a_193_47# A[10] 0
C50885 _0736_/a_56_297# _0350_ 0
C50886 clkload3/Y _0195_ 0.05809f
C50887 _1030_/a_1059_315# net57 0
C50888 _0195_ _1030_/a_466_413# 0.02932f
C50889 _0216_ _1030_/a_193_47# 0.00177f
C50890 clkload1/Y _0987_/a_27_47# 0
C50891 net48 _1005_/a_466_413# 0.00826f
C50892 _0118_ _0218_ 0
C50893 VPWR _0986_/a_193_47# 0.32066f
C50894 _0081_ _0114_ 0
C50895 _0471_ _0160_ 0
C50896 VPWR acc0.A\[25\] 1.24872f
C50897 _0292_ net67 0.39473f
C50898 _0293_ _0089_ 0
C50899 _0241_ _0461_ 0.02935f
C50900 hold21/a_285_47# acc0.A\[6\] 0
C50901 _0550_/a_51_297# _0176_ 0.02417f
C50902 _0714_/a_245_297# _0345_ 0
C50903 _1019_/a_381_47# _0345_ 0.01657f
C50904 _0343_ acc0.A\[30\] 0.01945f
C50905 net117 _0567_/a_27_297# 0
C50906 _0742_/a_81_21# _0742_/a_299_297# 0.08213f
C50907 _0804_/a_215_47# _0994_/a_27_47# 0
C50908 _1031_/a_193_47# hold62/a_285_47# 0
C50909 net237 _0359_ 0.20566f
C50910 net8 net157 0
C50911 acc0.A\[12\] _0403_ 0
C50912 _0715_/a_27_47# _0294_ 0
C50913 clknet_1_0__leaf__0459_ clkbuf_0__0459_/a_110_47# 0.0129f
C50914 _0500_/a_27_47# acc0.A\[15\] 0.027f
C50915 _0255_ _0824_/a_59_75# 0.03553f
C50916 _0473_ net174 0.04215f
C50917 net126 output36/a_27_47# 0
C50918 control0.state\[0\] _0972_/a_256_47# 0
C50919 control0.state\[1\] _0972_/a_250_297# 0.08798f
C50920 net213 _0183_ 0
C50921 _0195_ _0126_ 0.5264f
C50922 net23 _1062_/a_193_47# 0
C50923 net187 VPWR 0.42295f
C50924 _0487_ _1065_/a_466_413# 0
C50925 acc0.A\[3\] net10 0.10184f
C50926 net58 _0253_ 0.00406f
C50927 clknet_0__0465_ _0172_ 0
C50928 net211 _0352_ 0
C50929 _0924_/a_27_47# _0463_ 0
C50930 _0248_ control0.add 0.0313f
C50931 net125 clknet_0__0464_ 0
C50932 net224 _0350_ 0.37355f
C50933 output36/a_27_47# input8/a_75_212# 0.01193f
C50934 _0225_ _0232_ 0.22068f
C50935 _0571_/a_27_297# VPWR 0.25373f
C50936 _1001_/a_1059_315# _0869_/a_27_47# 0.00158f
C50937 net95 _1009_/a_466_413# 0
C50938 _0478_ _0979_/a_27_297# 0
C50939 _0960_/a_181_47# _0480_ 0
C50940 _0098_ _0216_ 0
C50941 _0378_ _0379_ 0.0039f
C50942 _0461_ _0772_/a_510_47# 0
C50943 net55 _0323_ 0
C50944 _1035_/a_27_47# _0208_ 0
C50945 _0606_/a_465_297# _0219_ 0
C50946 _0601_/a_150_297# _0102_ 0
C50947 _1047_/a_27_47# _1047_/a_193_47# 0.96668f
C50948 comp0.B\[8\] _1040_/a_466_413# 0.01317f
C50949 _0206_ _1040_/a_634_159# 0.01615f
C50950 VPWR _0148_ 0.40687f
C50951 _0516_/a_27_297# acc0.A\[8\] 0.01212f
C50952 _0516_/a_109_297# net66 0
C50953 _0714_/a_51_297# hold16/a_285_47# 0
C50954 net180 _0463_ 0
C50955 net53 _0366_ 0.53633f
C50956 net47 _0988_/a_193_47# 0
C50957 _1041_/a_27_47# _0174_ 0.0027f
C50958 clknet_1_0__leaf__0460_ _0758_/a_215_47# 0.00517f
C50959 hold82/a_285_47# net229 0.0102f
C50960 VPWR _0845_/a_109_47# 0.00632f
C50961 _0582_/a_109_297# net221 0.0639f
C50962 _0380_ net50 0.07068f
C50963 _0328_ hold90/a_49_47# 0
C50964 _1041_/a_634_159# comp0.B\[10\] 0
C50965 _0080_ hold2/a_285_47# 0.0012f
C50966 net68 hold2/a_391_47# 0
C50967 _0499_/a_59_75# control0.reset 0.00641f
C50968 _1052_/a_1059_315# _1052_/a_891_413# 0.31086f
C50969 _1052_/a_193_47# _1052_/a_975_413# 0
C50970 _1052_/a_466_413# _1052_/a_381_47# 0.03733f
C50971 _1001_/a_27_47# clknet_1_0__leaf__0461_ 0
C50972 _0478_ _1071_/a_561_413# 0
C50973 _0324_ _0686_/a_219_297# 0
C50974 _1007_/a_27_47# _1007_/a_561_413# 0.0027f
C50975 _1007_/a_634_159# _1007_/a_891_413# 0.03684f
C50976 _1007_/a_193_47# _1007_/a_381_47# 0.09799f
C50977 net36 net204 0
C50978 hold96/a_49_47# _1004_/a_27_47# 0.00422f
C50979 clknet_1_0__leaf__0460_ _0487_ 0.15517f
C50980 VPWR _0737_/a_117_297# 0.00858f
C50981 hold10/a_391_47# _0177_ 0
C50982 _1012_/a_1059_315# _1010_/a_1059_315# 0
C50983 _0243_ _1006_/a_634_159# 0
C50984 _0282_ net37 0.01036f
C50985 hold88/a_49_47# _1055_/a_27_47# 0
C50986 _0346_ _0158_ 0
C50987 _0837_/a_81_21# _0837_/a_368_297# 0.01485f
C50988 _1058_/a_634_159# _1058_/a_592_47# 0
C50989 _0195_ _0531_/a_109_47# 0
C50990 net186 _1034_/a_891_413# 0
C50991 _0172_ _1044_/a_634_159# 0.03574f
C50992 net187 net48 0
C50993 clkload4/Y _0459_ 0.0058f
C50994 _0477_ hold84/a_285_47# 0
C50995 _0179_ _1052_/a_634_159# 0.01614f
C50996 net228 _0419_ 0
C50997 A[8] output63/a_27_47# 0.00176f
C50998 clknet_1_0__leaf__0462_ hold52/a_391_47# 0.00981f
C50999 net24 net27 0
C51000 VPWR input31/a_75_212# 0.26531f
C51001 _0500_/a_27_47# _0179_ 0.35214f
C51002 _0172_ net184 0.00571f
C51003 net69 net222 0.00166f
C51004 _0212_ _1035_/a_1059_315# 0.01024f
C51005 net185 _1035_/a_891_413# 0
C51006 _1050_/a_634_159# net154 0.01419f
C51007 _0680_/a_472_297# _0311_ 0.00486f
C51008 net36 hold27/a_49_47# 0
C51009 VPWR _0722_/a_215_47# 0.00586f
C51010 clknet_1_0__leaf__0458_ _0630_/a_109_297# 0
C51011 _0310_ _0397_ 0.21363f
C51012 acc0.A\[12\] _0510_/a_373_47# 0
C51013 _0304_ net41 0
C51014 net47 net72 0
C51015 _0337_ _0349_ 0.00507f
C51016 net97 _0726_/a_240_47# 0
C51017 _1011_/a_1059_315# _0109_ 0.02485f
C51018 _1011_/a_592_47# _0354_ 0
C51019 net57 _0726_/a_51_297# 0
C51020 _1011_/a_975_413# _0355_ 0.00111f
C51021 clk clknet_1_0__leaf_clk 0.05316f
C51022 VPWR _1013_/a_561_413# 0.00292f
C51023 net119 _1065_/a_466_413# 0
C51024 _1002_/a_891_413# VPWR 0.19366f
C51025 _0343_ _0310_ 0
C51026 net152 net129 0
C51027 net157 net10 0
C51028 _0226_ clknet_1_0__leaf__0460_ 0
C51029 _0399_ acc0.A\[8\] 0.76812f
C51030 _0329_ _0727_/a_193_47# 0.00103f
C51031 _0742_/a_384_47# acc0.A\[24\] 0
C51032 _0656_/a_59_75# clknet_1_1__leaf__0465_ 0.01877f
C51033 _0273_ _0434_ 0.27051f
C51034 _0251_ output61/a_27_47# 0
C51035 _0538_/a_240_47# comp0.B\[14\] 0.00244f
C51036 _0312_ _0745_/a_193_47# 0
C51037 _0369_ _0828_/a_113_297# 0.00179f
C51038 clkbuf_1_0__f_clk/a_110_47# _0468_ 0
C51039 _1058_/a_634_159# _0186_ 0
C51040 _0327_ _0727_/a_277_47# 0.00597f
C51041 clkbuf_0_clk/a_110_47# _0974_/a_222_93# 0.01f
C51042 _0975_/a_59_75# _0975_/a_145_75# 0.00658f
C51043 clkbuf_0__0463_/a_110_47# comp0.B\[5\] 0
C51044 clknet_0__0464_ _0473_ 0.09427f
C51045 _0195_ net104 0.03004f
C51046 _0346_ _0391_ 0
C51047 _1027_/a_592_47# acc0.A\[26\] 0
C51048 _0136_ net171 0.13868f
C51049 net58 net74 0.20556f
C51050 _0422_ _0295_ 0
C51051 net217 _0304_ 0
C51052 _0399_ _0991_/a_193_47# 0
C51053 _1037_/a_27_47# _0173_ 0
C51054 hold80/a_49_47# hold80/a_285_47# 0.22264f
C51055 _0379_ acc0.A\[24\] 0
C51056 _1063_/a_1059_315# _0880_/a_27_47# 0.00158f
C51057 net67 _0655_/a_215_53# 0
C51058 _0324_ acc0.A\[23\] 0
C51059 hold70/a_391_47# _0418_ 0
C51060 VPWR _0525_/a_384_47# 0
C51061 _0197_ _1048_/a_1059_315# 0.00106f
C51062 net205 _1034_/a_561_413# 0
C51063 _1050_/a_27_47# hold7/a_285_47# 0
C51064 net64 _0516_/a_27_297# 0
C51065 _0265_ _0263_ 0
C51066 _0727_/a_193_47# _0221_ 0
C51067 _0984_/a_891_413# VPWR 0.18811f
C51068 net63 _0620_/a_113_47# 0
C51069 _0220_ hold92/a_49_47# 0
C51070 net63 _0989_/a_27_47# 0.03268f
C51071 _0693_/a_68_297# _1006_/a_1059_315# 0
C51072 clkbuf_1_1__f__0464_/a_110_47# clknet_0__0464_ 0.31628f
C51073 net63 hold1/a_49_47# 0.02222f
C51074 clknet_1_0__leaf__0457_ _0460_ 0.1794f
C51075 _0994_/a_561_413# _0218_ 0
C51076 _0172_ _0546_/a_149_47# 0.03122f
C51077 _0495_/a_150_297# _0175_ 0
C51078 control0.state\[1\] _0217_ 0
C51079 net138 _1052_/a_193_47# 0.01325f
C51080 acc0.A\[14\] _0346_ 0.02976f
C51081 clkbuf_1_0__f__0464_/a_110_47# _0527_/a_109_297# 0
C51082 _0459_ clknet_1_0__leaf__0461_ 0.4423f
C51083 net58 output61/a_27_47# 0
C51084 _0995_/a_1017_47# pp[14] 0.00174f
C51085 hold13/a_391_47# _1039_/a_891_413# 0
C51086 net211 net207 0
C51087 net111 _1026_/a_891_413# 0
C51088 hold44/a_285_47# acc0.A\[28\] 0.00176f
C51089 _1011_/a_27_47# acc0.A\[29\] 0.0084f
C51090 _1004_/a_27_47# net90 0.22947f
C51091 _0570_/a_109_297# _1026_/a_891_413# 0
C51092 _0369_ _0990_/a_634_159# 0
C51093 _0217_ _0583_/a_109_47# 0.00464f
C51094 _0183_ _0583_/a_27_297# 0.26879f
C51095 hold41/a_49_47# acc0.A\[10\] 0.31606f
C51096 net21 _0174_ 0
C51097 clkbuf_1_0__f__0462_/a_110_47# _1007_/a_466_413# 0.00563f
C51098 _1002_/a_891_413# net48 0.00459f
C51099 _0429_ _0642_/a_215_297# 0
C51100 _0251_ _0642_/a_382_47# 0
C51101 VPWR _1042_/a_592_47# 0
C51102 _0982_/a_381_47# _0346_ 0
C51103 net101 _0721_/a_27_47# 0.01167f
C51104 _0482_ _0962_/a_109_297# 0.00177f
C51105 hold97/a_49_47# clknet_1_1__leaf__0460_ 0.00493f
C51106 _1070_/a_27_47# _0979_/a_109_297# 0
C51107 _1070_/a_193_47# _0979_/a_27_297# 0.00104f
C51108 hold43/a_49_47# _1028_/a_27_47# 0
C51109 hold98/a_391_47# _0797_/a_207_413# 0
C51110 net231 _0164_ 0
C51111 _0578_/a_109_297# _0462_ 0
C51112 net54 _0195_ 0.05177f
C51113 _1030_/a_381_47# acc0.A\[30\] 0.00112f
C51114 _0273_ acc0.A\[7\] 0
C51115 _0273_ _0989_/a_1059_315# 0
C51116 clknet_0__0464_ _0186_ 0.0068f
C51117 _0457_ clknet_1_0__leaf__0457_ 0.24119f
C51118 clknet_1_1__leaf__0463_ _0955_/a_32_297# 0.00149f
C51119 hold56/a_285_47# _1065_/a_27_47# 0.00164f
C51120 hold16/a_49_47# hold62/a_49_47# 0
C51121 _0988_/a_466_413# _0988_/a_561_413# 0.00772f
C51122 _0988_/a_634_159# _0988_/a_975_413# 0
C51123 _0531_/a_27_297# net247 0
C51124 _0553_/a_51_297# _0553_/a_512_297# 0.0116f
C51125 _0352_ net241 0.0089f
C51126 _0313_ _0462_ 0
C51127 net187 clknet_1_0__leaf__0459_ 0.061f
C51128 output55/a_27_47# _0568_/a_27_297# 0
C51129 _1053_/a_193_47# acc0.A\[7\] 0
C51130 hold100/a_49_47# _0465_ 0.00766f
C51131 net138 net12 0.00336f
C51132 VPWR _0532_/a_384_47# 0
C51133 _0982_/a_193_47# _0465_ 0.00253f
C51134 _1063_/a_27_47# _1062_/a_1059_315# 0.00914f
C51135 _0629_/a_59_75# acc0.A\[14\] 0
C51136 acc0.A\[2\] hold100/a_49_47# 0
C51137 _0694_/a_113_47# clknet_1_0__leaf__0460_ 0
C51138 _0785_/a_81_21# acc0.A\[9\] 0.00165f
C51139 net225 _1031_/a_466_413# 0
C51140 _0111_ _1031_/a_193_47# 0
C51141 _0542_/a_245_297# net195 0
C51142 _0542_/a_149_47# _0203_ 0.00154f
C51143 _0542_/a_51_297# net19 0.10226f
C51144 net64 _0399_ 0.02853f
C51145 _0355_ _0334_ 0
C51146 hold101/a_49_47# VPWR 0.32292f
C51147 _1056_/a_634_159# _0369_ 0
C51148 net243 _0575_/a_27_297# 0.0012f
C51149 _0959_/a_80_21# _1062_/a_27_47# 0
C51150 A[13] _0994_/a_891_413# 0
C51151 _0432_ _0840_/a_68_297# 0.00504f
C51152 _0443_ _0840_/a_150_297# 0
C51153 _0982_/a_193_47# acc0.A\[2\] 0
C51154 _0179_ A[8] 0.00651f
C51155 _0768_/a_27_47# _0397_ 0
C51156 _0999_/a_891_413# _0097_ 0
C51157 _1003_/a_381_47# net240 0
C51158 _0316_ _0686_/a_219_297# 0.12812f
C51159 _0640_/a_215_297# net62 0
C51160 hold79/a_49_47# _0489_ 0.00357f
C51161 _0961_/a_113_297# _0978_/a_27_297# 0.01922f
C51162 _1021_/a_193_47# _0460_ 0.00813f
C51163 _0399_ _0423_ 0
C51164 _0118_ _0099_ 0
C51165 _1021_/a_466_413# clknet_1_0__leaf__0457_ 0.00573f
C51166 output67/a_27_47# pp[10] 0.01469f
C51167 pp[9] output37/a_27_47# 0.08034f
C51168 _0316_ _1008_/a_1059_315# 0
C51169 net167 _0484_ 0.00741f
C51170 _0244_ _0612_/a_145_75# 0.00149f
C51171 _0769_/a_299_297# acc0.A\[18\] 0
C51172 input23/a_75_212# net27 0
C51173 net23 input27/a_75_212# 0.10967f
C51174 net133 _1047_/a_193_47# 0.016f
C51175 _0081_ net104 0
C51176 net46 _0247_ 0.05866f
C51177 _0265_ clknet_1_0__leaf__0461_ 0
C51178 hold22/a_391_47# _0180_ 0
C51179 _0141_ net20 0.04735f
C51180 comp0.B\[9\] _1040_/a_891_413# 0
C51181 _0626_/a_68_297# _0256_ 0.228f
C51182 _0433_ _0369_ 0.00391f
C51183 _0580_/a_27_297# acc0.A\[19\] 0.10747f
C51184 _0583_/a_27_297# acc0.A\[15\] 0
C51185 output44/a_27_47# pp[30] 0.01905f
C51186 _0279_ _0994_/a_891_413# 0
C51187 _0795_/a_384_47# net5 0
C51188 clkbuf_1_0__f__0457_/a_110_47# net46 0.00111f
C51189 _0400_ _0345_ 0.27435f
C51190 _0792_/a_303_47# _0219_ 0.00401f
C51191 _0107_ _0370_ 0
C51192 _0959_/a_80_21# _0561_/a_51_297# 0
C51193 _0285_ _0420_ 0
C51194 _0144_ _1061_/a_27_47# 0
C51195 _0536_/a_51_297# net147 0
C51196 _0557_/a_245_297# _0175_ 0.00305f
C51197 _0228_ _0760_/a_285_47# 0
C51198 _0605_/a_109_297# _0237_ 0.0148f
C51199 _0254_ _0186_ 0.16915f
C51200 _0347_ _1008_/a_1059_315# 0
C51201 _1037_/a_891_413# _0135_ 0.04513f
C51202 _0531_/a_27_297# _1048_/a_466_413# 0
C51203 _0531_/a_109_297# _1048_/a_634_159# 0
C51204 _0996_/a_193_47# hold91/a_49_47# 0
C51205 _0996_/a_27_47# hold91/a_285_47# 0
C51206 hold97/a_285_47# clkbuf_1_1__f__0462_/a_110_47# 0.00119f
C51207 _0235_ control0.add 0
C51208 net62 _0465_ 0.01356f
C51209 hold38/a_285_47# hold38/a_391_47# 0.41909f
C51210 clknet_1_0__leaf__0462_ _0576_/a_373_47# 0
C51211 _0465_ _0450_ 0.00966f
C51212 pp[30] _1030_/a_975_413# 0
C51213 hold34/a_49_47# hold34/a_391_47# 0.00188f
C51214 clkload1/Y clkbuf_1_0__f__0465_/a_110_47# 0.00274f
C51215 hold13/a_49_47# _0957_/a_32_297# 0.00281f
C51216 _0239_ _0397_ 0
C51217 net44 pp[28] 0
C51218 clknet_0__0463_ clknet_1_1__leaf__0457_ 0.01086f
C51219 VPWR _0103_ 0.51406f
C51220 _0642_/a_27_413# _0988_/a_27_47# 0
C51221 _0513_/a_299_297# acc0.A\[10\] 0
C51222 _0343_ _0184_ 0
C51223 net58 _0446_ 0.20621f
C51224 _0133_ _0959_/a_80_21# 0
C51225 VPWR hold91/a_391_47# 0.18237f
C51226 hold18/a_285_47# VPWR 0.29385f
C51227 _0985_/a_891_413# _0448_ 0
C51228 net234 _0455_ 0
C51229 _0218_ _0668_/a_297_47# 0.00847f
C51230 hold30/a_49_47# net177 0.00116f
C51231 _1001_/a_634_159# _1001_/a_975_413# 0
C51232 _1001_/a_466_413# _1001_/a_561_413# 0.00772f
C51233 _0422_ _0811_/a_299_297# 0.00182f
C51234 acc0.A\[21\] _0594_/a_113_47# 0
C51235 net172 net8 0.07132f
C51236 _0305_ _0307_ 0.0184f
C51237 net60 output60/a_27_47# 0.18973f
C51238 _1062_/a_634_159# _1062_/a_381_47# 0
C51239 _0708_/a_68_297# pp[31] 0
C51240 _0342_ _0567_/a_109_297# 0.02406f
C51241 _1011_/a_1059_315# _0725_/a_80_21# 0
C51242 _0992_/a_193_47# net228 0
C51243 acc0.A\[5\] _0193_ 0.00372f
C51244 _0831_/a_285_297# _0253_ 0.00749f
C51245 _1021_/a_193_47# _1021_/a_466_413# 0.07593f
C51246 _1021_/a_27_47# _1021_/a_1059_315# 0.04875f
C51247 pp[27] _0354_ 0.00796f
C51248 _1003_/a_1059_315# net49 0.10321f
C51249 _0575_/a_27_297# _1024_/a_381_47# 0
C51250 _0430_ _0827_/a_27_47# 0.04133f
C51251 _0086_ _0434_ 0
C51252 _0347_ acc0.A\[23\] 0
C51253 net53 net112 0
C51254 _0590_/a_113_47# net50 0
C51255 _0642_/a_215_297# clknet_1_1__leaf__0458_ 0
C51256 net210 VPWR 0.5156f
C51257 VPWR net57 1.83723f
C51258 net179 net62 0
C51259 _0476_ hold84/a_49_47# 0.03177f
C51260 control0.state\[0\] _0971_/a_299_297# 0
C51261 control0.state\[1\] _0971_/a_81_21# 0
C51262 _0459_ _1060_/a_891_413# 0.00817f
C51263 net53 acc0.A\[24\] 0
C51264 _0222_ net176 0
C51265 net115 _1008_/a_193_47# 0
C51266 net191 _1008_/a_27_47# 0
C51267 _1029_/a_193_47# net94 0
C51268 _0267_ _0263_ 0.43573f
C51269 _1000_/a_891_413# _0183_ 0
C51270 hold87/a_49_47# hold59/a_285_47# 0.00189f
C51271 _0963_/a_117_297# control0.count\[0\] 0.00795f
C51272 net194 net183 0.00277f
C51273 VPWR _0548_/a_51_297# 0.47699f
C51274 _0856_/a_215_47# VPWR 0.00191f
C51275 net34 _0975_/a_59_75# 0.06609f
C51276 _0968_/a_109_297# _0486_ 0.01204f
C51277 net48 _0103_ 0.02944f
C51278 clknet_1_0__leaf__0465_ _0836_/a_68_297# 0.00133f
C51279 clknet_1_1__leaf__0464_ _1043_/a_1059_315# 0.09041f
C51280 acc0.A\[18\] _0392_ 0
C51281 _0234_ _0756_/a_47_47# 0
C51282 clknet_1_1__leaf__0459_ _0302_ 0.00391f
C51283 _0216_ _1015_/a_27_47# 0
C51284 _0104_ acc0.A\[23\] 0
C51285 _0372_ _0610_/a_59_75# 0
C51286 clknet_1_1__leaf__0459_ _0795_/a_299_297# 0
C51287 _0172_ _0176_ 0.47148f
C51288 _0317_ _0685_/a_68_297# 0.10751f
C51289 _0817_/a_81_21# _0816_/a_68_297# 0.00157f
C51290 net45 _0779_/a_215_47# 0
C51291 _0326_ _0219_ 0.04312f
C51292 A[13] _0668_/a_79_21# 0
C51293 _0585_/a_109_297# clknet_1_0__leaf__0461_ 0
C51294 VPWR _0670_/a_510_47# 0.00135f
C51295 clknet_1_0__leaf__0465_ net212 0
C51296 _0092_ _0994_/a_466_413# 0
C51297 hold55/a_391_47# _0461_ 0
C51298 _1034_/a_193_47# clkbuf_1_1__f__0463_/a_110_47# 0.00641f
C51299 _1020_/a_466_413# _0721_/a_27_47# 0.00575f
C51300 _0951_/a_296_53# comp0.B\[0\] 0
C51301 _0257_ net63 0.00716f
C51302 hold38/a_49_47# _1034_/a_27_47# 0
C51303 hold40/a_391_47# hold73/a_285_47# 0
C51304 net216 _0346_ 0.03044f
C51305 _1004_/a_592_47# _0216_ 0.00112f
C51306 _0224_ _1022_/a_1059_315# 0
C51307 _0714_/a_512_297# _0344_ 0
C51308 _0589_/a_113_47# acc0.A\[28\] 0
C51309 _0561_/a_51_297# _0173_ 0.11557f
C51310 control0.state\[1\] _0164_ 0.00142f
C51311 _0983_/a_891_413# _0195_ 0
C51312 _0717_/a_80_21# output44/a_27_47# 0
C51313 _1072_/a_891_413# _1068_/a_891_413# 0
C51314 _0476_ _1065_/a_381_47# 0
C51315 _0219_ hold95/a_391_47# 0
C51316 _0359_ _0320_ 0
C51317 acc0.A\[12\] acc0.A\[13\] 0
C51318 net181 _0514_/a_109_297# 0
C51319 _0146_ acc0.A\[3\] 0
C51320 _0221_ hold62/a_285_47# 0
C51321 _0760_/a_47_47# clknet_1_0__leaf__0460_ 0.00316f
C51322 _0200_ net174 0.0021f
C51323 hold20/a_285_47# clknet_1_0__leaf_clk 0
C51324 _0125_ VPWR 1.04392f
C51325 comp0.B\[13\] net21 0
C51326 _1036_/a_891_413# clknet_1_1__leaf__0463_ 0.01734f
C51327 _1036_/a_466_413# net122 0
C51328 _1052_/a_634_159# hold83/a_49_47# 0.00168f
C51329 _1052_/a_27_47# hold83/a_391_47# 0.00285f
C51330 _1052_/a_193_47# hold83/a_285_47# 0.00241f
C51331 _0770_/a_297_47# _0771_/a_27_413# 0
C51332 _0478_ _0169_ 0.00165f
C51333 hold68/a_49_47# _0222_ 0
C51334 _0343_ _0315_ 0.09977f
C51335 _0461_ _1019_/a_466_413# 0.00442f
C51336 _0101_ acc0.A\[21\] 0.02486f
C51337 _0201_ _1046_/a_1059_315# 0
C51338 clknet_0__0458_ _0990_/a_27_47# 0.00109f
C51339 _1001_/a_27_47# _0218_ 0
C51340 _0133_ _0173_ 0.42113f
C51341 _0343_ output47/a_27_47# 0
C51342 hold67/a_285_47# hold67/a_391_47# 0.41909f
C51343 _1041_/a_27_47# comp0.B\[9\] 0
C51344 _1041_/a_466_413# net153 0.01475f
C51345 _1041_/a_1059_315# net127 0
C51346 _1047_/a_466_413# _1047_/a_592_47# 0.00553f
C51347 _1047_/a_634_159# _1047_/a_1017_47# 0
C51348 A[12] acc0.A\[9\] 0
C51349 comp0.B\[8\] net174 0.69582f
C51350 _0307_ _0675_/a_150_297# 0
C51351 _0190_ acc0.A\[8\] 0
C51352 _0305_ _0780_/a_285_297# 0.00183f
C51353 _0423_ _0295_ 0
C51354 hold25/a_49_47# VPWR 0.28223f
C51355 _0131_ _0563_/a_240_47# 0.03331f
C51356 comp0.B\[1\] _0563_/a_245_297# 0
C51357 _0285_ _0284_ 0.56122f
C51358 net185 _0561_/a_512_297# 0
C51359 output53/a_27_47# net53 0.1789f
C51360 _0230_ hold94/a_49_47# 0.09114f
C51361 pp[18] _0195_ 0
C51362 _0985_/a_466_413# _0183_ 0
C51363 net40 pp[31] 0
C51364 _0343_ _0718_/a_129_47# 0.00107f
C51365 _0461_ net219 0
C51366 hold41/a_49_47# _0188_ 0.00715f
C51367 _0217_ _1018_/a_1059_315# 0.00272f
C51368 _0567_/a_27_297# _0704_/a_68_297# 0
C51369 _0354_ _0724_/a_199_47# 0.00261f
C51370 net178 _0153_ 0.05554f
C51371 _1007_/a_891_413# net93 0
C51372 _0243_ _0195_ 0
C51373 hold22/a_49_47# _0152_ 0.36572f
C51374 _0536_/a_51_297# _0473_ 0.02751f
C51375 net243 _1004_/a_1059_315# 0.05435f
C51376 net12 hold83/a_285_47# 0.03649f
C51377 _0525_/a_81_21# acc0.A\[6\] 0
C51378 _0432_ _0255_ 0.45259f
C51379 _0837_/a_266_47# _0442_ 0.04093f
C51380 _0172_ net130 0.04536f
C51381 _1020_/a_1017_47# _0352_ 0.00226f
C51382 _0446_ _0262_ 0.02123f
C51383 net197 _1027_/a_975_413# 0
C51384 _0570_/a_27_297# net156 0.00655f
C51385 net23 net17 0.02561f
C51386 hold7/a_285_47# _0987_/a_27_47# 0.00104f
C51387 hold7/a_49_47# _0987_/a_193_47# 0
C51388 control0.sh input28/a_75_212# 0
C51389 _1057_/a_27_47# net37 0
C51390 hold98/a_285_47# acc0.A\[31\] 0
C51391 _0234_ hold66/a_391_47# 0
C51392 _0752_/a_27_413# net213 0.00176f
C51393 _0268_ _0843_/a_150_297# 0
C51394 net180 clkbuf_1_0__f__0463_/a_110_47# 0.14513f
C51395 _0251_ net61 0.13373f
C51396 clknet_1_1__leaf__0459_ net6 0.01782f
C51397 net44 _0608_/a_27_47# 0.03899f
C51398 _0682_/a_68_297# acc0.A\[26\] 0
C51399 _0971_/a_384_47# _0163_ 0
C51400 comp0.B\[12\] _0140_ 0.00143f
C51401 _0195_ net227 0
C51402 hold58/a_49_47# _0175_ 0
C51403 _0216_ _0354_ 0.0369f
C51404 VPWR _0505_/a_109_47# 0
C51405 _0269_ _0219_ 0.02311f
C51406 _0558_/a_150_297# _0212_ 0
C51407 _1061_/a_975_413# comp0.B\[9\] 0
C51408 _1057_/a_634_159# net67 0.01321f
C51409 net61 _0989_/a_592_47# 0
C51410 pp[15] pp[14] 0.26822f
C51411 net193 net174 0
C51412 _0438_ _0825_/a_68_297# 0
C51413 _0179_ _0517_/a_81_21# 0.00101f
C51414 acc0.A\[28\] _0219_ 0.00543f
C51415 _0983_/a_891_413# _0081_ 0
C51416 net69 _0854_/a_215_47# 0
C51417 acc0.A\[17\] _0097_ 0
C51418 net169 _0152_ 0
C51419 _0666_/a_113_47# clknet_1_1__leaf__0459_ 0
C51420 _0389_ _0369_ 0
C51421 clknet_1_1__leaf__0460_ _0685_/a_150_297# 0
C51422 _1063_/a_634_159# _1063_/a_592_47# 0
C51423 _0494_/a_27_47# _0560_/a_68_297# 0.00124f
C51424 net144 _0186_ 0
C51425 _0833_/a_79_21# _0988_/a_634_159# 0
C51426 _0833_/a_215_47# _0988_/a_27_47# 0
C51427 _0307_ _0181_ 0.0323f
C51428 hold58/a_285_47# control0.sh 0.00808f
C51429 _0195_ _0407_ 0
C51430 _0573_/a_27_47# _0584_/a_27_297# 0
C51431 net157 _0492_/a_27_47# 0.06229f
C51432 _0219_ net209 0
C51433 hold75/a_391_47# clknet_1_0__leaf__0458_ 0.00117f
C51434 _0305_ _0507_/a_109_297# 0.00718f
C51435 _0326_ _0746_/a_81_21# 0.00885f
C51436 _0400_ _0791_/a_113_297# 0.05206f
C51437 _0405_ _0791_/a_199_47# 0
C51438 _0959_/a_217_297# _0959_/a_472_297# 0.00517f
C51439 _0959_/a_80_21# _0959_/a_300_47# 0.00997f
C51440 net63 net11 0
C51441 hold27/a_49_47# _1061_/a_27_47# 0.01003f
C51442 _0218_ _0459_ 0.12195f
C51443 _0429_ net63 0.04243f
C51444 _0585_/a_27_297# _0585_/a_109_297# 0.17136f
C51445 B[9] B[14] 0.16965f
C51446 _0121_ _0576_/a_27_297# 0.11664f
C51447 net61 net58 0.1271f
C51448 clknet_1_0__leaf__0464_ _1050_/a_193_47# 0.00212f
C51449 _1049_/a_27_47# acc0.A\[15\] 0
C51450 net36 _0632_/a_113_47# 0
C51451 VPWR _1048_/a_27_47# 0.66771f
C51452 net232 _1062_/a_27_47# 0.00668f
C51453 net64 _0190_ 0
C51454 _0200_ clknet_0__0464_ 0.00112f
C51455 hold11/a_391_47# _0147_ 0
C51456 _1028_/a_1059_315# clknet_1_1__leaf__0462_ 0.00485f
C51457 VPWR _0506_/a_384_47# 0
C51458 hold46/a_49_47# _0473_ 0.00179f
C51459 control0.count\[3\] _1071_/a_1059_315# 0
C51460 net214 net66 0.02597f
C51461 _0530_/a_81_21# clknet_1_1__leaf__0457_ 0
C51462 _0556_/a_68_297# control0.sh 0
C51463 _0237_ net241 0
C51464 _0381_ _0219_ 0.03862f
C51465 _0819_/a_299_297# clknet_0__0465_ 0.04283f
C51466 hold47/a_285_47# _0186_ 0
C51467 _0515_/a_384_47# net66 0
C51468 _0349_ _0333_ 0
C51469 _0195_ _0569_/a_109_297# 0.04505f
C51470 net178 _0990_/a_27_47# 0
C51471 hold101/a_391_47# _0835_/a_78_199# 0
C51472 _0570_/a_27_297# acc0.A\[26\] 0.01798f
C51473 _0183_ _0114_ 0.02678f
C51474 VPWR _1010_/a_1059_315# 0.43246f
C51475 _0183_ _0615_/a_109_297# 0.00175f
C51476 clkbuf_1_0__f__0462_/a_110_47# _0105_ 0.00803f
C51477 _1000_/a_193_47# _1000_/a_466_413# 0.07379f
C51478 _1000_/a_27_47# _1000_/a_1059_315# 0.04875f
C51479 _1060_/a_634_159# _1060_/a_592_47# 0
C51480 _0513_/a_299_297# _0188_ 0.00863f
C51481 _1051_/a_891_413# _0527_/a_27_297# 0
C51482 hold57/a_49_47# control0.sh 0.04326f
C51483 _1070_/a_193_47# _0169_ 0
C51484 VPWR _0979_/a_27_297# 0.19282f
C51485 hold48/a_391_47# net18 0.00178f
C51486 _1051_/a_1059_315# _0346_ 0
C51487 _0192_ _0520_/a_109_47# 0
C51488 net230 _0520_/a_109_297# 0.00199f
C51489 _0462_ _0616_/a_493_297# 0
C51490 net196 net128 0
C51491 _1053_/a_891_413# net11 0.02052f
C51492 _0236_ _0346_ 0.17831f
C51493 net53 _0691_/a_68_297# 0
C51494 _0343_ control0.add 0.09953f
C51495 VPWR _0846_/a_512_297# 0.00729f
C51496 clknet_1_1__leaf__0463_ _0474_ 0.0366f
C51497 _0343_ _0742_/a_81_21# 0.1693f
C51498 _0568_/a_27_297# acc0.A\[30\] 0
C51499 _0553_/a_51_297# _0136_ 0.14109f
C51500 _0805_/a_27_47# VPWR 0.23051f
C51501 _0399_ _0986_/a_466_413# 0.01453f
C51502 net53 _0682_/a_150_297# 0.00181f
C51503 _0329_ _0350_ 0.58264f
C51504 control0.state\[1\] net34 0.21109f
C51505 _0476_ _0471_ 0.19538f
C51506 VPWR _1009_/a_891_413# 0.19678f
C51507 hold36/a_49_47# clknet_1_1__leaf__0464_ 0
C51508 hold14/a_49_47# _0173_ 0
C51509 _0579_/a_373_47# net187 0.00197f
C51510 _0625_/a_59_75# _0186_ 0.01725f
C51511 _0857_/a_27_47# _1033_/a_1059_315# 0
C51512 clknet_1_0__leaf__0460_ _0350_ 0.3084f
C51513 _0216_ _0452_ 0
C51514 acc0.A\[21\] net35 0.00293f
C51515 _0655_/a_215_53# _0302_ 0
C51516 _0375_ acc0.A\[22\] 0
C51517 _0161_ _1062_/a_193_47# 0.00834f
C51518 _0316_ clknet_1_1__leaf__0462_ 0.00284f
C51519 _1071_/a_561_413# VPWR 0.00314f
C51520 _0973_/a_109_47# _0460_ 0
C51521 clkbuf_1_1__f__0465_/a_110_47# net67 0
C51522 _0309_ _0397_ 0.51178f
C51523 _1056_/a_27_47# net178 0.00394f
C51524 hold37/a_285_47# clkbuf_0__0464_/a_110_47# 0.00235f
C51525 _0330_ _0701_/a_80_21# 0.17687f
C51526 _0195_ _0567_/a_109_47# 0.00195f
C51527 _0216_ _0567_/a_27_297# 0.17291f
C51528 _0276_ _0399_ 0.26149f
C51529 _0985_/a_466_413# _0179_ 0.02313f
C51530 _0984_/a_1059_315# hold75/a_391_47# 0.01554f
C51531 net42 acc0.A\[13\] 0.10267f
C51532 _0948_/a_109_297# _0477_ 0
C51533 net214 _0350_ 0.06576f
C51534 _0254_ net62 0
C51535 _0179_ _1049_/a_27_47# 0.05774f
C51536 clknet_1_1__leaf__0462_ _0347_ 0.05886f
C51537 _0221_ _0350_ 0
C51538 _1059_/a_634_159# _0219_ 0
C51539 _0119_ clknet_1_0__leaf__0457_ 0.04255f
C51540 _0701_/a_209_297# _0333_ 0.00231f
C51541 net193 clknet_0__0464_ 0
C51542 net36 acc0.A\[1\] 0.28899f
C51543 output36/a_27_47# net8 0
C51544 _0573_/a_27_47# _1015_/a_634_159# 0
C51545 _0461_ _0352_ 0.02012f
C51546 _0117_ acc0.A\[19\] 0.00182f
C51547 clknet_0__0464_ _1046_/a_466_413# 0.0336f
C51548 _0114_ acc0.A\[15\] 0
C51549 _0997_/a_27_47# net41 0.42275f
C51550 clknet_1_1__leaf__0460_ _0738_/a_150_297# 0
C51551 _0154_ acc0.A\[9\] 0.0016f
C51552 clkbuf_1_1__f__0463_/a_110_47# _0565_/a_240_47# 0
C51553 comp0.B\[14\] _0473_ 0.12735f
C51554 _0462_ clkbuf_0__0460_/a_110_47# 0.0788f
C51555 _1071_/a_27_47# clknet_0_clk 0.00528f
C51556 _1071_/a_466_413# clkbuf_1_0__f_clk/a_110_47# 0.00322f
C51557 output54/a_27_47# _1027_/a_381_47# 0
C51558 net54 _1027_/a_466_413# 0.02044f
C51559 _1008_/a_1059_315# _0106_ 0.01156f
C51560 _1008_/a_381_47# _0365_ 0.00737f
C51561 _0177_ _1047_/a_193_47# 0
C51562 _0959_/a_80_21# _0208_ 0
C51563 VPWR _0954_/a_220_297# 0.01167f
C51564 hold13/a_49_47# _0213_ 0.08612f
C51565 _0337_ _1030_/a_193_47# 0
C51566 _0178_ _1047_/a_27_47# 0.0302f
C51567 hold89/a_285_47# _0471_ 0
C51568 _0313_ _0312_ 0
C51569 comp0.B\[11\] _1043_/a_466_413# 0
C51570 _0346_ _0422_ 0.00459f
C51571 _0958_/a_27_47# _1062_/a_381_47# 0
C51572 _1020_/a_193_47# _0578_/a_109_297# 0
C51573 net53 net111 0.00325f
C51574 _1000_/a_27_47# _1018_/a_193_47# 0
C51575 clkbuf_1_0__f__0459_/a_110_47# _0184_ 0
C51576 net183 _1045_/a_27_47# 0.00533f
C51577 clknet_1_0__leaf__0465_ _0527_/a_373_47# 0
C51578 _0134_ control0.sh 0
C51579 pp[8] A[10] 0.02945f
C51580 hold13/a_391_47# _0475_ 0.00139f
C51581 VPWR _1022_/a_381_47# 0.07542f
C51582 clknet_1_1__leaf__0460_ _0311_ 0.0524f
C51583 _1034_/a_193_47# _0163_ 0
C51584 _0637_/a_56_297# _0465_ 0.00157f
C51585 _0174_ _0173_ 0.33002f
C51586 VPWR _0779_/a_215_47# 0.00684f
C51587 _0852_/a_117_297# _0266_ 0.00142f
C51588 net85 net42 0
C51589 clknet_1_1__leaf__0459_ _0993_/a_891_413# 0
C51590 _0284_ _0218_ 0
C51591 _0993_/a_561_413# net38 0
C51592 net22 hold6/a_49_47# 0
C51593 B[14] hold6/a_285_47# 0
C51594 _0999_/a_193_47# _0999_/a_381_47# 0.09799f
C51595 _0999_/a_634_159# _0999_/a_891_413# 0.03684f
C51596 _0999_/a_27_47# _0999_/a_561_413# 0.0027f
C51597 _0854_/a_79_21# _0399_ 0.12339f
C51598 net17 _1063_/a_466_413# 0.02794f
C51599 _0992_/a_193_47# _0090_ 0.23108f
C51600 _1017_/a_193_47# _0115_ 0.25034f
C51601 _0972_/a_250_297# clknet_1_1__leaf_clk 0.04168f
C51602 _1001_/a_27_47# _0099_ 0.07952f
C51603 net2 _0992_/a_27_47# 0
C51604 hold26/a_285_47# clkbuf_1_0__f__0463_/a_110_47# 0
C51605 comp0.B\[7\] control0.sh 0
C51606 _0342_ _1031_/a_27_47# 0
C51607 _1001_/a_466_413# net223 0.00459f
C51608 _0341_ _1031_/a_1059_315# 0.00912f
C51609 _0340_ _1031_/a_466_413# 0
C51610 _1001_/a_634_159# _0391_ 0
C51611 clknet_1_0__leaf__0465_ _0989_/a_891_413# 0
C51612 net63 clknet_1_1__leaf__0458_ 0.18048f
C51613 net120 _1034_/a_891_413# 0
C51614 net121 input25/a_75_212# 0.01082f
C51615 net61 _0262_ 0
C51616 _1062_/a_891_413# _0160_ 0
C51617 net23 B[2] 0.04282f
C51618 B[15] net25 0
C51619 _0118_ _1032_/a_193_47# 0
C51620 _1020_/a_193_47# net202 0.00542f
C51621 _0310_ clkbuf_0__0461_/a_110_47# 0.00109f
C51622 comp0.B\[14\] _0186_ 0
C51623 net67 _0673_/a_253_47# 0
C51624 _0600_/a_103_199# _0219_ 0.0065f
C51625 B[9] _0544_/a_51_297# 0
C51626 clknet_1_0__leaf__0465_ _1061_/a_466_413# 0.00505f
C51627 hold49/a_49_47# comp0.B\[14\] 0
C51628 _1021_/a_193_47# _0119_ 0.43347f
C51629 _1021_/a_891_413# _1021_/a_1017_47# 0.00617f
C51630 _0181_ _0507_/a_109_297# 0.02317f
C51631 _0233_ net213 0
C51632 _0575_/a_373_47# _0122_ 0
C51633 _1017_/a_975_413# _0459_ 0
C51634 _0147_ _1048_/a_592_47# 0
C51635 _1049_/a_1017_47# net134 0
C51636 _0576_/a_27_297# _0380_ 0
C51637 _0180_ _0830_/a_215_47# 0
C51638 hold41/a_285_47# _0187_ 0
C51639 clkload3/a_268_47# net43 0
C51640 hold55/a_285_47# net23 0.0224f
C51641 net242 _0347_ 0
C51642 _0648_/a_27_297# _0648_/a_205_297# 0.00412f
C51643 clknet_1_1__leaf__0459_ _0790_/a_285_297# 0
C51644 _0510_/a_27_297# net4 0.18073f
C51645 VPWR _0540_/a_149_47# 0.00197f
C51646 _0135_ net27 0
C51647 hold17/a_285_47# _0979_/a_27_297# 0.00104f
C51648 net162 net60 0
C51649 _0257_ clkbuf_0__0465_/a_110_47# 0
C51650 _0733_/a_79_199# _0361_ 0.11143f
C51651 _1056_/a_1059_315# acc0.A\[12\] 0.02108f
C51652 net62 _0988_/a_561_413# 0
C51653 _1043_/a_27_47# net20 0
C51654 _0456_ _0447_ 0
C51655 net245 net42 0.00117f
C51656 _1011_/a_634_159# _0219_ 0
C51657 _1011_/a_381_47# _0345_ 0
C51658 net126 _1041_/a_27_47# 0
C51659 _0178_ clknet_1_0__leaf__0461_ 0.01127f
C51660 net48 _1022_/a_381_47# 0.00579f
C51661 pp[26] _1026_/a_1059_315# 0
C51662 _1031_/a_891_413# _1013_/a_1059_315# 0
C51663 _1006_/a_193_47# _0345_ 0
C51664 clknet_0__0461_ _0219_ 0
C51665 _0375_ _0379_ 0
C51666 _0195_ net208 0.42246f
C51667 net150 _0224_ 0
C51668 control0.count\[1\] _0978_/a_27_297# 0
C51669 _0168_ _0978_/a_373_47# 0.00236f
C51670 _0673_/a_103_199# _0288_ 0
C51671 _0118_ _0721_/a_27_47# 0
C51672 net23 _0165_ 0.11022f
C51673 _0986_/a_193_47# _0345_ 0
C51674 hold46/a_391_47# _0535_/a_68_297# 0.01241f
C51675 acc0.A\[25\] _0345_ 0
C51676 net9 comp0.B\[12\] 0
C51677 _0833_/a_79_21# _0253_ 0.00997f
C51678 control0.count\[2\] _1071_/a_466_413# 0.03157f
C51679 _0111_ _0344_ 0
C51680 _0642_/a_27_413# _0642_/a_215_297# 0.14121f
C51681 _1055_/a_1059_315# _0189_ 0
C51682 clkbuf_1_0__f__0457_/a_110_47# _0902_/a_27_47# 0.00542f
C51683 hold37/a_391_47# _0143_ 0
C51684 _0173_ _0208_ 0.35595f
C51685 _0462_ _1009_/a_27_47# 0
C51686 VPWR _1067_/a_975_413# 0.00499f
C51687 _0222_ _1023_/a_466_413# 0.00149f
C51688 _1050_/a_381_47# _0186_ 0
C51689 _0554_/a_68_297# control0.sh 0.00456f
C51690 net53 _0361_ 0.01382f
C51691 _1033_/a_381_47# clknet_1_0__leaf__0461_ 0
C51692 _0267_ _0848_/a_27_47# 0.04859f
C51693 _0582_/a_27_297# net219 0.09877f
C51694 _1019_/a_1059_315# _0869_/a_27_47# 0
C51695 net187 _0345_ 0
C51696 _0359_ _1007_/a_1059_315# 0
C51697 _0753_/a_79_21# _0753_/a_381_47# 0.00247f
C51698 hold34/a_285_47# _0153_ 0
C51699 _0762_/a_79_21# _0754_/a_51_297# 0
C51700 acc0.A\[14\] net221 0
C51701 _0111_ _0709_/a_113_47# 0
C51702 _0618_/a_297_297# _0250_ 0
C51703 net154 net73 0.09525f
C51704 net186 _0215_ 0
C51705 _0218_ _0267_ 0.50779f
C51706 net161 net122 0.00253f
C51707 _0780_/a_35_297# _0677_/a_285_47# 0
C51708 net4 _0181_ 0.12016f
C51709 net180 _0548_/a_245_297# 0
C51710 _0461_ net207 0.00612f
C51711 VPWR _1027_/a_634_159# 0.202f
C51712 net183 net132 0
C51713 net204 _1037_/a_27_47# 0
C51714 _0218_ _0772_/a_79_21# 0.06908f
C51715 _0346_ _0370_ 0.00549f
C51716 _0210_ comp0.B\[2\] 0.00229f
C51717 clknet_0__0457_ _0713_/a_27_47# 0.00585f
C51718 net44 _0678_/a_68_297# 0
C51719 _0640_/a_109_53# _0431_ 0
C51720 comp0.B\[15\] _0214_ 0
C51721 _0258_ clkbuf_1_1__f__0458_/a_110_47# 0
C51722 net45 net42 0.00525f
C51723 _0135_ _0136_ 0
C51724 _1000_/a_634_159# _0242_ 0
C51725 pp[17] pp[31] 0.00841f
C51726 net118 _0181_ 0.1988f
C51727 _0805_/a_27_47# _0283_ 0.027f
C51728 hold46/a_391_47# _0174_ 0.00133f
C51729 clknet_1_1__leaf__0462_ hold95/a_49_47# 0
C51730 _0338_ _0568_/a_373_47# 0
C51731 _0698_/a_113_297# clkbuf_1_1__f__0462_/a_110_47# 0
C51732 output51/a_27_47# pp[23] 0.15655f
C51733 _0982_/a_1059_315# _0850_/a_68_297# 0.00125f
C51734 clkload0/a_27_47# _0468_ 0
C51735 clk _0970_/a_27_297# 0.00874f
C51736 _0346_ acc0.A\[8\] 0.00718f
C51737 _0459_ _0581_/a_109_47# 0
C51738 hold61/a_49_47# net209 0
C51739 _0167_ _0162_ 0
C51740 _0343_ hold74/a_391_47# 0.00782f
C51741 _1042_/a_27_47# hold51/a_285_47# 0
C51742 net185 _0132_ 0.06482f
C51743 _0082_ _0219_ 0.11642f
C51744 _0105_ net51 0
C51745 hold85/a_49_47# _0161_ 0
C51746 net86 _0675_/a_68_297# 0
C51747 _0083_ _0183_ 0
C51748 clknet_1_0__leaf__0457_ _0373_ 0
C51749 net122 net26 0
C51750 VPWR _0764_/a_81_21# 0.2097f
C51751 hold86/a_391_47# _0265_ 0
C51752 _0399_ _1014_/a_193_47# 0
C51753 _0546_/a_149_47# _1040_/a_193_47# 0
C51754 _1019_/a_27_47# clknet_1_0__leaf__0461_ 0
C51755 _0456_ acc0.A\[0\] 0.17915f
C51756 _0183_ net104 0
C51757 _0257_ _0824_/a_59_75# 0
C51758 _0645_/a_377_297# acc0.A\[13\] 0
C51759 _1004_/a_193_47# _0379_ 0.00101f
C51760 _1004_/a_1059_315# _0378_ 0
C51761 net65 acc0.A\[8\] 0.41978f
C51762 net55 _0730_/a_215_47# 0.05575f
C51763 acc0.A\[8\] _0989_/a_466_413# 0.029f
C51764 _0460_ _0246_ 0
C51765 VPWR _0700_/a_113_47# 0
C51766 hold74/a_285_47# acc0.A\[17\] 0.00143f
C51767 _0307_ clknet_1_1__leaf__0461_ 0.24068f
C51768 pp[17] hold15/a_285_47# 0.04361f
C51769 _0123_ _1007_/a_381_47# 0
C51770 net200 _1007_/a_1059_315# 0
C51771 _0346_ _0991_/a_193_47# 0.02945f
C51772 _0768_/a_27_47# clkbuf_0__0461_/a_110_47# 0
C51773 _0974_/a_222_93# _0487_ 0.0319f
C51774 _0712_/a_465_47# _0340_ 0.00444f
C51775 _0126_ net156 0.27005f
C51776 clknet_1_0__leaf__0464_ _0987_/a_193_47# 0
C51777 hold88/a_49_47# _0988_/a_1059_315# 0.00621f
C51778 _0345_ _0737_/a_117_297# 0.00221f
C51779 _0180_ _0843_/a_68_297# 0
C51780 _0273_ _0186_ 0
C51781 input17/a_75_212# B[0] 0.19279f
C51782 _0730_/a_297_297# _0347_ 0.00562f
C51783 _0747_/a_510_47# _0460_ 0
C51784 VPWR _0524_/a_373_47# 0
C51785 net133 _0178_ 0.04537f
C51786 B[5] B[6] 0.10414f
C51787 _0461_ _0613_/a_109_297# 0
C51788 _1034_/a_634_159# _1034_/a_381_47# 0
C51789 _0536_/a_149_47# _0536_/a_240_47# 0.06872f
C51790 _0536_/a_51_297# _0200_ 0.11551f
C51791 hold6/a_285_47# _0544_/a_51_297# 0
C51792 _0796_/a_215_47# net238 0.05555f
C51793 _0462_ _0771_/a_27_413# 0
C51794 VPWR input34/a_27_47# 0.28476f
C51795 net59 acc0.A\[29\] 0
C51796 _1021_/a_891_413# acc0.A\[21\] 0.00342f
C51797 _0559_/a_51_297# net205 0.10604f
C51798 _0621_/a_35_297# _0434_ 0
C51799 hold75/a_49_47# _0852_/a_35_297# 0
C51800 clknet_1_0__leaf__0458_ hold2/a_285_47# 0.00947f
C51801 _0428_ _0291_ 0.01945f
C51802 hold25/a_285_47# net180 0.00228f
C51803 _0982_/a_592_47# clknet_1_0__leaf__0461_ 0
C51804 _0217_ net234 0.31006f
C51805 _0398_ _0781_/a_68_297# 0.11317f
C51806 _0660_/a_113_47# _0291_ 0
C51807 _1013_/a_466_413# _0219_ 0.00379f
C51808 _0587_/a_27_47# net42 0
C51809 _0343_ _0583_/a_109_47# 0
C51810 clknet_0__0464_ _1045_/a_193_47# 0.00205f
C51811 clkbuf_0__0464_/a_110_47# _1045_/a_381_47# 0
C51812 _1063_/a_975_413# _0161_ 0
C51813 _0086_ _0988_/a_466_413# 0
C51814 net235 _0988_/a_381_47# 0
C51815 _0833_/a_79_21# net74 0.01143f
C51816 _0239_ clkbuf_0__0461_/a_110_47# 0
C51817 control0.state\[0\] _1068_/a_1059_315# 0
C51818 _0981_/a_27_297# _0468_ 0.00205f
C51819 _0252_ clknet_0__0465_ 0
C51820 hold16/a_285_47# _0340_ 0
C51821 _0359_ clkbuf_1_0__f__0462_/a_110_47# 0.02333f
C51822 VPWR _1026_/a_891_413# 0.19136f
C51823 _0535_/a_68_297# net153 0
C51824 _0585_/a_27_297# _0178_ 0
C51825 _0483_ _1072_/a_1059_315# 0
C51826 control0.count\[3\] _1072_/a_381_47# 0.0166f
C51827 VPWR clkbuf_1_1__f__0460_/a_110_47# 1.2557f
C51828 acc0.A\[12\] VPWR 2.28061f
C51829 hold96/a_285_47# net50 0.05263f
C51830 net48 _0764_/a_81_21# 0.02078f
C51831 _0217_ net46 0.03101f
C51832 output43/a_27_47# net41 0.06238f
C51833 net78 _0992_/a_381_47# 0
C51834 _0750_/a_181_47# net51 0
C51835 _0218_ _0638_/a_109_297# 0.00175f
C51836 net243 net176 0
C51837 VPWR _1024_/a_592_47# 0
C51838 _0083_ acc0.A\[15\] 0.00106f
C51839 _0585_/a_109_297# _0112_ 0.0063f
C51840 hold66/a_49_47# VPWR 0.31396f
C51841 net135 _0142_ 0
C51842 net203 _0214_ 0.07062f
C51843 net242 hold95/a_49_47# 0
C51844 hold64/a_285_47# _0452_ 0
C51845 hold64/a_49_47# _0266_ 0
C51846 _1018_/a_193_47# acc0.A\[19\] 0
C51847 clknet_1_0__leaf__0460_ _1005_/a_1059_315# 0
C51848 net18 net195 0.20766f
C51849 net198 net19 0
C51850 net1 hold73/a_285_47# 0
C51851 hold52/a_285_47# acc0.A\[25\] 0.05974f
C51852 _0519_/a_81_21# _0437_ 0
C51853 net114 net113 0
C51854 _0350_ hold94/a_285_47# 0
C51855 _1017_/a_634_159# _1017_/a_1059_315# 0
C51856 _1017_/a_27_47# _1017_/a_381_47# 0.05761f
C51857 _1017_/a_193_47# _1017_/a_891_413# 0.19226f
C51858 _0487_ _1062_/a_634_159# 0.02111f
C51859 clkbuf_1_1__f__0461_/a_110_47# net43 0.21087f
C51860 _1058_/a_1059_315# _0512_/a_27_297# 0
C51861 net64 _0346_ 0
C51862 clknet_1_1__leaf__0460_ hold50/a_49_47# 0
C51863 _0516_/a_27_297# _0369_ 0
C51864 _1052_/a_27_47# net9 0.05649f
C51865 pp[27] _0353_ 0.00579f
C51866 hold47/a_391_47# net194 0.13575f
C51867 pp[6] net141 0
C51868 _0420_ net228 0.00104f
C51869 hold24/a_49_47# net180 0
C51870 _0473_ _1046_/a_561_413# 0
C51871 _0984_/a_193_47# _0219_ 0
C51872 _0472_ _1046_/a_891_413# 0
C51873 clkbuf_0__0463_/a_110_47# control0.reset 0.02443f
C51874 output64/a_27_47# _0988_/a_27_47# 0
C51875 _0126_ acc0.A\[26\] 0.00447f
C51876 _1006_/a_193_47# net52 0.00481f
C51877 _1000_/a_193_47# _0098_ 0.18107f
C51878 _1000_/a_891_413# _1000_/a_1017_47# 0.00617f
C51879 _1000_/a_634_159# net86 0
C51880 _0715_/a_27_47# _0291_ 0
C51881 _1056_/a_27_47# hold34/a_285_47# 0
C51882 _1056_/a_193_47# hold34/a_49_47# 0
C51883 net64 net65 0
C51884 _0822_/a_109_297# _0252_ 0
C51885 _0993_/a_381_47# _0281_ 0
C51886 _0388_ _0308_ 0
C51887 acc0.A\[28\] net94 0
C51888 _0195_ _0096_ 0.02618f
C51889 _0129_ _1013_/a_634_159# 0
C51890 net163 _1013_/a_27_47# 0
C51891 VPWR _0169_ 0.23572f
C51892 net230 _0186_ 0.06547f
C51893 _0346_ _0423_ 0.08471f
C51894 _0459_ net228 0
C51895 _0174_ net153 0
C51896 _0130_ clknet_1_0__leaf__0457_ 0
C51897 _1072_/a_592_47# VPWR 0
C51898 hold46/a_49_47# _0200_ 0.04614f
C51899 output45/a_27_47# acc0.A\[31\] 0.03715f
C51900 pp[18] hold15/a_49_47# 0
C51901 _0804_/a_79_21# _0804_/a_215_47# 0.04584f
C51902 VPWR _0445_ 0.199f
C51903 clknet_1_1__leaf__0463_ _0563_/a_51_297# 0
C51904 _0263_ _0347_ 0
C51905 clkbuf_0__0463_/a_110_47# _1061_/a_891_413# 0
C51906 clkbuf_1_1__f__0463_/a_110_47# _0171_ 0
C51907 _0556_/a_68_297# net172 0
C51908 _0536_/a_149_47# _1046_/a_27_47# 0
C51909 _0536_/a_51_297# _1046_/a_466_413# 0.00183f
C51910 _0461_ net106 0
C51911 acc0.A\[25\] net52 0
C51912 _0985_/a_27_47# _0197_ 0.00564f
C51913 _0520_/a_109_47# clknet_1_0__leaf__0465_ 0
C51914 _0128_ acc0.A\[30\] 0
C51915 acc0.A\[5\] hold1/a_285_47# 0.071f
C51916 _0287_ _0817_/a_266_47# 0
C51917 _0528_/a_81_21# _0527_/a_27_297# 0
C51918 net240 _1063_/a_381_47# 0
C51919 _0973_/a_27_297# _0161_ 0.18722f
C51920 net56 net57 0.00255f
C51921 hold96/a_49_47# net215 0.00631f
C51922 net243 hold68/a_49_47# 0
C51923 hold82/a_49_47# hold82/a_391_47# 0.00188f
C51924 hold46/a_49_47# comp0.B\[8\] 0
C51925 _0401_ _0992_/a_193_47# 0.00136f
C51926 _0347_ _1007_/a_466_413# 0
C51927 _0352_ _1007_/a_27_47# 0.00358f
C51928 clknet_1_0__leaf__0460_ _1006_/a_634_159# 0
C51929 _0195_ _1031_/a_193_47# 0.12829f
C51930 _0963_/a_285_297# _0481_ 0.07201f
C51931 acc0.A\[20\] _1032_/a_27_47# 0
C51932 _0457_ _1033_/a_1017_47# 0
C51933 _0751_/a_183_297# clknet_1_0__leaf__0460_ 0
C51934 _0231_ _0618_/a_215_47# 0.04931f
C51935 _0234_ _0374_ 0.1176f
C51936 hold70/a_49_47# _0419_ 0
C51937 VPWR _0650_/a_68_297# 0.15191f
C51938 _0480_ clkbuf_1_0__f_clk/a_110_47# 0.0125f
C51939 _1072_/a_634_159# clknet_0_clk 0.01256f
C51940 _1050_/a_634_159# _1050_/a_381_47# 0
C51941 _0643_/a_253_47# VPWR 0.00168f
C51942 _0470_ _0160_ 0.08767f
C51943 _1019_/a_381_47# clknet_1_0__leaf__0457_ 0
C51944 _0083_ _0179_ 0.67493f
C51945 _0399_ _0369_ 1.15682f
C51946 hold85/a_285_47# _0946_/a_30_53# 0
C51947 _1024_/a_27_47# net50 0.04252f
C51948 clknet_1_1__leaf__0462_ _0106_ 0.00496f
C51949 clknet_0__0457_ _0399_ 0.01247f
C51950 _0221_ _1011_/a_561_413# 0.00276f
C51951 _0551_/a_27_47# _0465_ 0.00125f
C51952 _0820_/a_79_21# acc0.A\[9\] 0.00404f
C51953 _0280_ _0402_ 0
C51954 _0427_ _0401_ 0.31491f
C51955 _0428_ _0290_ 0.02417f
C51956 hold26/a_391_47# _0548_/a_51_297# 0.01261f
C51957 _0335_ acc0.A\[29\] 0.19394f
C51958 _0465_ _0849_/a_79_21# 0.00208f
C51959 _1036_/a_193_47# net28 0
C51960 _0565_/a_51_297# _0565_/a_149_47# 0.02487f
C51961 _0660_/a_113_47# _0290_ 0
C51962 _0241_ net223 0
C51963 _0680_/a_217_297# VPWR 0.22542f
C51964 _0461_ _0769_/a_299_297# 0
C51965 _0222_ net241 0.3051f
C51966 _0998_/a_1059_315# net43 0.11648f
C51967 _0640_/a_109_53# _0269_ 0.00322f
C51968 _1054_/a_193_47# _1052_/a_1059_315# 0
C51969 _1054_/a_27_47# _1052_/a_891_413# 0.00437f
C51970 _0971_/a_81_21# clknet_1_1__leaf_clk 0.0013f
C51971 net54 net156 0.10741f
C51972 hold88/a_285_47# _0186_ 0.0399f
C51973 _0795_/a_81_21# _0297_ 0
C51974 _0982_/a_466_413# net149 0
C51975 _0176_ _1040_/a_193_47# 0.02526f
C51976 _0620_/a_113_47# _0180_ 0
C51977 _1039_/a_634_159# _0463_ 0.00633f
C51978 _0180_ _0989_/a_27_47# 0
C51979 pp[11] VPWR 0.31611f
C51980 acc0.A\[22\] VPWR 0.97202f
C51981 comp0.B\[12\] net129 0
C51982 comp0.B\[11\] net196 0
C51983 _0566_/a_27_47# clkbuf_1_1__f__0457_/a_110_47# 0.00183f
C51984 _1056_/a_466_413# _0179_ 0.03968f
C51985 clkbuf_0__0465_/a_110_47# clknet_1_1__leaf__0458_ 0
C51986 _0533_/a_109_297# control0.reset 0
C51987 _0195_ net71 0.04136f
C51988 _0477_ _1062_/a_381_47# 0.00707f
C51989 hold46/a_391_47# comp0.B\[13\] 0.0015f
C51990 hold46/a_49_47# net193 0.00377f
C51991 clknet_1_1__leaf__0461_ _0507_/a_109_297# 0
C51992 _0975_/a_59_75# _0166_ 0
C51993 _0486_ _1068_/a_975_413# 0.00184f
C51994 _0200_ comp0.B\[14\] 0.08867f
C51995 net46 _0248_ 0.26709f
C51996 clknet_1_0__leaf__0461_ _0347_ 0.00786f
C51997 _0353_ _0724_/a_199_47# 0
C51998 _0555_/a_245_297# _0173_ 0
C51999 _0999_/a_27_47# _0998_/a_1059_315# 0
C52000 input5/a_75_212# A[13] 0.20019f
C52001 hold46/a_391_47# _1046_/a_193_47# 0
C52002 _0533_/a_27_297# _0465_ 0.00335f
C52003 hold10/a_285_47# _0180_ 0.00605f
C52004 hold10/a_49_47# net8 0.00142f
C52005 clkload4/Y _1016_/a_891_413# 0
C52006 net123 _0209_ 0
C52007 _0574_/a_27_297# _1007_/a_193_47# 0
C52008 _0343_ _1000_/a_561_413# 0
C52009 _1033_/a_1059_315# _0208_ 0
C52010 _0292_ _0275_ 0.24373f
C52011 _0317_ clknet_0__0460_ 0.00719f
C52012 net39 _0801_/a_113_47# 0
C52013 _0999_/a_891_413# net85 0
C52014 net17 _0161_ 0.41715f
C52015 _0412_ _0795_/a_81_21# 0
C52016 _1050_/a_193_47# clkbuf_1_0__f__0464_/a_110_47# 0
C52017 _0345_ _0103_ 0.00142f
C52018 _0772_/a_79_21# _0099_ 0.05029f
C52019 _0772_/a_215_47# _0391_ 0.00549f
C52020 clkbuf_1_1__f__0458_/a_110_47# _0988_/a_193_47# 0
C52021 _0772_/a_510_47# net223 0.00245f
C52022 _0164_ clknet_1_1__leaf_clk 0.00745f
C52023 _0086_ _0186_ 0.02168f
C52024 comp0.B\[14\] comp0.B\[8\] 0
C52025 _0310_ _0777_/a_377_297# 0
C52026 VPWR _0993_/a_592_47# 0
C52027 _1016_/a_634_159# net221 0.01584f
C52028 _0752_/a_300_297# _0234_ 0.00308f
C52029 net58 _0269_ 0.2269f
C52030 net201 comp0.B\[0\] 0.09243f
C52031 clknet_1_0__leaf__0462_ _1007_/a_592_47# 0.00151f
C52032 _0732_/a_80_21# _0732_/a_209_47# 0.01013f
C52033 _0715_/a_27_47# _0290_ 0
C52034 hold91/a_391_47# _0345_ 0.00736f
C52035 _0971_/a_299_297# clkbuf_1_1__f_clk/a_110_47# 0
C52036 hold18/a_285_47# _0345_ 0.00464f
C52037 _0207_ _0546_/a_149_47# 0
C52038 hold31/a_285_47# acc0.A\[6\] 0.00135f
C52039 _0983_/a_891_413# _0183_ 0
C52040 VPWR _0542_/a_245_297# 0.00684f
C52041 _0775_/a_215_47# _0775_/a_510_47# 0.00529f
C52042 _0305_ _0287_ 0.00955f
C52043 _0186_ _0987_/a_381_47# 0
C52044 _0996_/a_891_413# _0790_/a_35_297# 0
C52045 clknet_0__0463_ _0564_/a_68_297# 0
C52046 _0216_ _0353_ 0
C52047 _0433_ net75 0
C52048 acc0.A\[1\] hold60/a_391_47# 0
C52049 _1043_/a_193_47# _0203_ 0
C52050 _0312_ clkbuf_0__0460_/a_110_47# 0.04437f
C52051 hold20/a_285_47# hold20/a_391_47# 0.41909f
C52052 clkbuf_1_0__f__0458_/a_110_47# hold75/a_49_47# 0.01845f
C52053 _0327_ _0334_ 0.00125f
C52054 comp0.B\[7\] net172 0
C52055 net185 net25 0.12221f
C52056 _1001_/a_891_413# net206 0
C52057 _0212_ B[2] 0
C52058 hold32/a_391_47# _0153_ 0.00339f
C52059 _0479_ _0975_/a_145_75# 0
C52060 _1016_/a_1059_315# _0459_ 0.00593f
C52061 _0174_ _0144_ 0
C52062 hold88/a_391_47# _0253_ 0
C52063 _0648_/a_205_297# _0280_ 0
C52064 _0195_ _0395_ 0
C52065 acc0.A\[22\] net48 0.02028f
C52066 output66/a_27_47# net3 0
C52067 net4 _0187_ 0.01429f
C52068 clknet_0__0464_ net73 0
C52069 hold17/a_285_47# _0169_ 0.00934f
C52070 control0.count\[2\] _0480_ 0.12914f
C52071 clknet_1_1__leaf__0459_ _0999_/a_193_47# 0
C52072 hold38/a_391_47# clknet_1_1__leaf_clk 0
C52073 _0147_ clknet_1_1__leaf__0457_ 0
C52074 VPWR net42 1.47742f
C52075 net196 _0202_ 0.0121f
C52076 net57 _0345_ 0.03198f
C52077 net97 _0219_ 0.00994f
C52078 _1002_/a_381_47# clknet_1_0__leaf__0460_ 0.00247f
C52079 net54 acc0.A\[26\] 0.91338f
C52080 clknet_0__0458_ _0840_/a_150_297# 0
C52081 _1006_/a_975_413# _0219_ 0
C52082 _0234_ _0249_ 0
C52083 _0136_ _0206_ 0
C52084 acc0.A\[12\] _0283_ 0.31648f
C52085 _0415_ _0218_ 0.02931f
C52086 net39 _0286_ 0
C52087 pp[12] A[13] 0.01138f
C52088 _0413_ net81 0.00103f
C52089 net185 _0477_ 0
C52090 _0614_/a_29_53# _0246_ 0.16741f
C52091 net10 _0541_/a_68_297# 0.01314f
C52092 hold86/a_49_47# _0446_ 0.03529f
C52093 _0461_ _0392_ 0.00184f
C52094 _0559_/a_51_297# net160 0
C52095 _0712_/a_297_297# _0195_ 0
C52096 _0985_/a_634_159# _0985_/a_592_47# 0
C52097 _0728_/a_59_75# net97 0.00115f
C52098 hold39/a_285_47# comp0.B\[6\] 0.02145f
C52099 net193 comp0.B\[14\] 0.45347f
C52100 clknet_1_0__leaf__0464_ net132 0.00441f
C52101 _0563_/a_149_47# _0562_/a_68_297# 0
C52102 _0326_ _1007_/a_193_47# 0
C52103 clknet_1_1__leaf__0458_ _0824_/a_59_75# 0.0096f
C52104 _1018_/a_1059_315# _1018_/a_891_413# 0.31086f
C52105 _1018_/a_193_47# _1018_/a_975_413# 0
C52106 _1018_/a_466_413# _1018_/a_381_47# 0.03733f
C52107 _0982_/a_1059_315# hold100/a_285_47# 0
C52108 net36 _1014_/a_634_159# 0
C52109 hold85/a_285_47# _0967_/a_109_93# 0.00145f
C52110 _0956_/a_114_297# clknet_1_0__leaf__0461_ 0
C52111 hold85/a_391_47# _0485_ 0.00168f
C52112 hold19/a_285_47# _1016_/a_27_47# 0.01366f
C52113 hold19/a_49_47# _1016_/a_193_47# 0.00127f
C52114 hold11/a_49_47# _0464_ 0.00334f
C52115 _0243_ _0183_ 0.03105f
C52116 comp0.B\[14\] _1046_/a_466_413# 0
C52117 _0596_/a_145_75# _0228_ 0
C52118 _0279_ pp[12] 0
C52119 pp[1] clknet_1_1__leaf__0465_ 0
C52120 _0222_ net177 0.03607f
C52121 _0982_/a_193_47# _0982_/a_891_413# 0.1937f
C52122 _0982_/a_27_47# _0982_/a_381_47# 0.06222f
C52123 _0982_/a_634_159# _0982_/a_1059_315# 0
C52124 acc0.A\[4\] _0186_ 0.01958f
C52125 _0592_/a_68_297# clknet_1_0__leaf__0460_ 0.00208f
C52126 VPWR _0742_/a_384_47# 0
C52127 _1011_/a_27_47# clknet_1_1__leaf__0462_ 0
C52128 _1049_/a_634_159# _1049_/a_466_413# 0.23992f
C52129 _1049_/a_193_47# _1049_/a_1059_315# 0.03405f
C52130 _1049_/a_27_47# _1049_/a_891_413# 0.03224f
C52131 _0343_ _1018_/a_1059_315# 0.02765f
C52132 _0285_ _0347_ 0
C52133 _0983_/a_891_413# acc0.A\[15\] 0.00235f
C52134 comp0.B\[1\] clknet_1_0__leaf__0461_ 0.16182f
C52135 _0524_/a_109_297# acc0.A\[6\] 0
C52136 _0115_ net219 0.00154f
C52137 _1019_/a_1017_47# _0459_ 0
C52138 _0324_ _0105_ 0
C52139 net180 _0540_/a_240_47# 0
C52140 _0753_/a_561_47# _0233_ 0.00175f
C52141 _0753_/a_465_47# _0231_ 0.00184f
C52142 _0965_/a_47_47# _0486_ 0
C52143 _0762_/a_79_21# _0219_ 0
C52144 clkbuf_0__0462_/a_110_47# _0315_ 0.04123f
C52145 _0465_ _0529_/a_27_297# 0
C52146 VPWR _0379_ 0.45333f
C52147 _1054_/a_466_413# A[8] 0
C52148 _1019_/a_27_47# _0218_ 0.00225f
C52149 _0362_ _0359_ 0
C52150 hold56/a_49_47# _0133_ 0
C52151 hold98/a_285_47# net40 0.00378f
C52152 hold46/a_391_47# comp0.B\[9\] 0
C52153 hold79/a_285_47# net226 0.02979f
C52154 _0369_ _0295_ 0.07015f
C52155 _1066_/a_634_159# _1066_/a_466_413# 0.23992f
C52156 _1066_/a_193_47# _1066_/a_1059_315# 0.03405f
C52157 _1066_/a_27_47# _1066_/a_891_413# 0.03206f
C52158 _0473_ _1045_/a_891_413# 0
C52159 VPWR _0372_ 1.62248f
C52160 hold37/a_391_47# _1050_/a_27_47# 0
C52161 hold37/a_285_47# _1050_/a_193_47# 0
C52162 clkbuf_1_0__f__0459_/a_110_47# hold74/a_391_47# 0
C52163 net56 _1010_/a_1059_315# 0.08707f
C52164 pp[10] _0512_/a_27_297# 0
C52165 net63 _0218_ 0.02732f
C52166 net193 _0543_/a_68_297# 0
C52167 acc0.A\[14\] net238 0.02782f
C52168 comp0.B\[2\] comp0.B\[0\] 0.02549f
C52169 net53 net199 0
C52170 net89 _0237_ 0.00228f
C52171 _0101_ _0381_ 0
C52172 net86 _0242_ 0.12904f
C52173 net45 _0999_/a_891_413# 0.00863f
C52174 _1001_/a_27_47# _0721_/a_27_47# 0
C52175 VPWR _1052_/a_381_47# 0.07064f
C52176 _1031_/a_1059_315# acc0.A\[30\] 0
C52177 _1023_/a_634_159# _1022_/a_1059_315# 0.00187f
C52178 _1023_/a_193_47# _1022_/a_891_413# 0.00445f
C52179 _0328_ _0326_ 0.12523f
C52180 _0833_/a_215_47# _0833_/a_510_47# 0.00529f
C52181 clknet_1_1__leaf__0460_ net98 0.00265f
C52182 _0967_/a_487_297# clk 0
C52183 _1068_/a_634_159# _1068_/a_466_413# 0.23992f
C52184 _1068_/a_193_47# _1068_/a_1059_315# 0.03405f
C52185 _1068_/a_27_47# _1068_/a_891_413# 0.03089f
C52186 clkload3/a_110_47# clkload3/Y 0.00568f
C52187 input1/a_27_47# A[0] 0.20312f
C52188 _0176_ _0214_ 0
C52189 _1056_/a_381_47# hold67/a_285_47# 0
C52190 acc0.A\[14\] _0446_ 0.00214f
C52191 _0134_ _1036_/a_891_413# 0.00122f
C52192 _0487_ _1063_/a_592_47# 0
C52193 VPWR _0971_/a_299_297# 0.28528f
C52194 _0655_/a_109_93# acc0.A\[10\] 0
C52195 _0283_ _0650_/a_68_297# 0.02763f
C52196 clkbuf_1_1__f__0464_/a_110_47# _1045_/a_891_413# 0
C52197 hold58/a_285_47# _0474_ 0
C52198 pp[9] _0512_/a_373_47# 0
C52199 VPWR hold40/a_49_47# 0.31928f
C52200 _0797_/a_297_47# _0297_ 0
C52201 _0312_ _1009_/a_27_47# 0
C52202 _1032_/a_1059_315# net23 0
C52203 _1035_/a_27_47# clknet_1_1__leaf__0463_ 0.01495f
C52204 _0992_/a_27_47# hold70/a_285_47# 0.00287f
C52205 _0818_/a_193_47# _0401_ 0
C52206 comp0.B\[10\] hold5/a_49_47# 0.32524f
C52207 _0204_ net18 0
C52208 net71 _1048_/a_193_47# 0
C52209 _0519_/a_81_21# _0252_ 0.01999f
C52210 _0519_/a_384_47# acc0.A\[7\] 0
C52211 net248 _0830_/a_79_21# 0
C52212 hold47/a_49_47# _1051_/a_27_47# 0
C52213 _0269_ _0262_ 0
C52214 _1051_/a_466_413# _0186_ 0.00291f
C52215 _0557_/a_240_47# net26 0.00346f
C52216 _1034_/a_634_159# comp0.B\[2\] 0.01617f
C52217 hold6/a_391_47# net18 0.00125f
C52218 output65/a_27_47# _0989_/a_891_413# 0
C52219 pp[7] _0989_/a_27_47# 0
C52220 acc0.A\[27\] _1008_/a_193_47# 0.02894f
C52221 _0710_/a_109_47# clknet_1_1__leaf__0462_ 0
C52222 _0275_ _0785_/a_299_297# 0.09358f
C52223 _0442_ _0433_ 0.02848f
C52224 _0413_ _0797_/a_207_413# 0
C52225 _0979_/a_373_47# _0488_ 0.00211f
C52226 _0983_/a_193_47# _0181_ 0
C52227 _0464_ _0159_ 0.00186f
C52228 clknet_1_1__leaf__0460_ _0126_ 0
C52229 hold64/a_49_47# _0399_ 0
C52230 net48 _0372_ 0
C52231 clknet_0__0464_ _1044_/a_27_47# 0.00238f
C52232 _1072_/a_27_47# _0466_ 0.00807f
C52233 net43 _0793_/a_149_47# 0.02927f
C52234 _0816_/a_68_297# _0426_ 0.113f
C52235 net36 _0216_ 0
C52236 _0967_/a_109_93# _0958_/a_27_47# 0.0012f
C52237 acc0.A\[12\] net182 0
C52238 _0225_ _0618_/a_215_47# 0
C52239 _0958_/a_27_47# _0487_ 0.00642f
C52240 _0228_ _0383_ 0.1748f
C52241 hold34/a_49_47# clknet_1_1__leaf__0465_ 0
C52242 _0787_/a_303_47# net246 0
C52243 net34 clknet_1_1__leaf_clk 0
C52244 _0534_/a_299_297# _1047_/a_1059_315# 0
C52245 _0346_ _1006_/a_466_413# 0.03397f
C52246 hold57/a_391_47# comp0.B\[6\] 0.00442f
C52247 hold57/a_49_47# _0474_ 0
C52248 _0170_ _0468_ 0
C52249 _0369_ _0619_/a_68_297# 0
C52250 _0756_/a_47_47# net50 0.09169f
C52251 control0.state\[1\] _0166_ 0
C52252 _0112_ _0178_ 0
C52253 _0287_ _0181_ 0
C52254 _0427_ _0089_ 0
C52255 _0207_ _0176_ 0.12639f
C52256 pp[30] _1031_/a_381_47# 0
C52257 _1032_/a_634_159# clknet_1_0__leaf__0461_ 0.01688f
C52258 _0257_ _0432_ 0.09708f
C52259 _0973_/a_109_297# _0487_ 0.0113f
C52260 hold41/a_285_47# clknet_1_1__leaf__0465_ 0
C52261 _0805_/a_27_47# _0808_/a_266_47# 0
C52262 _1071_/a_592_47# _0466_ 0
C52263 _1071_/a_1017_47# _0488_ 0
C52264 _0343_ _0998_/a_27_47# 0.00431f
C52265 _1021_/a_1059_315# _0352_ 0.01094f
C52266 _0390_ _0372_ 0
C52267 hold8/a_285_47# _0365_ 0
C52268 _0403_ _0281_ 0.00247f
C52269 _0993_/a_975_413# _0286_ 0
C52270 _0853_/a_150_297# _0264_ 0
C52271 _0481_ _0946_/a_30_53# 0
C52272 _0645_/a_47_47# _0996_/a_27_47# 0
C52273 _1017_/a_1059_315# net103 0
C52274 _0357_ _0356_ 0.21776f
C52275 _1017_/a_27_47# _1016_/a_634_159# 0.00954f
C52276 _1017_/a_634_159# _1016_/a_27_47# 0.00275f
C52277 _1017_/a_193_47# _1016_/a_193_47# 0
C52278 _0231_ _0234_ 0.05123f
C52279 clknet_1_0__leaf__0459_ net42 0.00136f
C52280 _0190_ _0369_ 0
C52281 acc0.A\[8\] _0988_/a_634_159# 0
C52282 _0181_ _0526_/a_27_47# 0.06492f
C52283 _0966_/a_27_47# _0480_ 0.00122f
C52284 _0276_ _0346_ 0.02819f
C52285 net10 _1040_/a_891_413# 0
C52286 net153 comp0.B\[9\] 0
C52287 VPWR input19/a_75_212# 0.19073f
C52288 acc0.A\[13\] net5 0.48849f
C52289 net34 _0479_ 0
C52290 _0390_ hold40/a_49_47# 0
C52291 _0645_/a_377_297# VPWR 0.00505f
C52292 _0733_/a_79_199# VPWR 0.31248f
C52293 _0804_/a_510_47# _0092_ 0
C52294 _1067_/a_27_47# _1065_/a_193_47# 0
C52295 _1067_/a_193_47# _1065_/a_27_47# 0
C52296 A[11] _0186_ 0.00354f
C52297 _1010_/a_27_47# _0219_ 0
C52298 net204 _0174_ 0.02911f
C52299 _0404_ _0797_/a_27_413# 0
C52300 net36 _0852_/a_285_297# 0
C52301 _0521_/a_384_47# net230 0.00908f
C52302 _0521_/a_81_21# _0151_ 0.17578f
C52303 _0144_ _1046_/a_193_47# 0.00188f
C52304 _1033_/a_634_159# _1033_/a_592_47# 0
C52305 hold3/a_285_47# net51 0
C52306 _0283_ net42 0
C52307 _0798_/a_113_297# _0410_ 0
C52308 _0195_ _0329_ 0.23795f
C52309 _0259_ acc0.A\[8\] 0.04843f
C52310 clknet_0__0458_ _0827_/a_27_47# 0
C52311 net55 _0362_ 0.0132f
C52312 net194 hold37/a_285_47# 0.03977f
C52313 _1012_/a_634_159# _1012_/a_592_47# 0
C52314 _1039_/a_1059_315# _0176_ 0.01262f
C52315 _0196_ net154 0
C52316 _0148_ _0527_/a_373_47# 0
C52317 hold55/a_49_47# _1033_/a_1059_315# 0
C52318 _0165_ _0161_ 0.03255f
C52319 _0115_ _0352_ 0.00201f
C52320 hold79/a_391_47# _0487_ 0
C52321 _0347_ _0105_ 0
C52322 clknet_1_0__leaf__0460_ net92 0.29325f
C52323 net76 _0988_/a_1059_315# 0
C52324 _0805_/a_27_47# _0345_ 0.00196f
C52325 _0399_ _0409_ 0.02918f
C52326 _0476_ _0475_ 0.0216f
C52327 hold27/a_49_47# _0174_ 0
C52328 _1019_/a_891_413# net149 0
C52329 _0749_/a_384_47# _0462_ 0
C52330 acc0.A\[23\] _0360_ 0
C52331 clknet_1_0__leaf__0458_ _0853_/a_68_297# 0.00275f
C52332 _1009_/a_193_47# _0219_ 0.09816f
C52333 hold86/a_49_47# net61 0.28592f
C52334 VPWR net244 0.16457f
C52335 _0259_ _0991_/a_193_47# 0
C52336 _1050_/a_634_159# acc0.A\[4\] 0.0372f
C52337 _0241_ clkbuf_0__0457_/a_110_47# 0
C52338 net44 _0677_/a_47_47# 0.42627f
C52339 _0744_/a_27_47# _0186_ 0
C52340 _0343_ _1030_/a_891_413# 0.00796f
C52341 _0990_/a_1017_47# _0181_ 0
C52342 hold47/a_391_47# net132 0
C52343 net35 _0381_ 0
C52344 _1055_/a_466_413# acc0.A\[9\] 0
C52345 hold26/a_285_47# _0540_/a_240_47# 0
C52346 _1041_/a_193_47# net152 0
C52347 _1041_/a_27_47# net32 0.00471f
C52348 net53 VPWR 2.17742f
C52349 _0967_/a_215_297# net17 0
C52350 hold88/a_285_47# net62 0.02106f
C52351 _0854_/a_79_21# _0346_ 0.0017f
C52352 clknet_0_clk _0951_/a_109_93# 0.01057f
C52353 _0195_ _0221_ 0.1288f
C52354 _0746_/a_299_297# clkbuf_0__0460_/a_110_47# 0
C52355 net36 net247 0
C52356 VPWR _0440_ 0.49498f
C52357 _0508_/a_81_21# _0508_/a_384_47# 0.00138f
C52358 net181 acc0.A\[9\] 0
C52359 _0180_ net11 0.20589f
C52360 comp0.B\[14\] _1045_/a_193_47# 0
C52361 _0218_ _0347_ 0.55593f
C52362 net149 net206 0.08738f
C52363 VPWR _1034_/a_27_47# 0.39352f
C52364 hold16/a_391_47# acc0.A\[30\] 0.03448f
C52365 _0960_/a_109_47# VPWR 0
C52366 _1004_/a_27_47# _0575_/a_109_297# 0
C52367 _1004_/a_193_47# _0575_/a_27_297# 0
C52368 comp0.B\[13\] hold37/a_391_47# 0
C52369 net140 _1052_/a_466_413# 0.00375f
C52370 net58 _0082_ 0.00292f
C52371 _1017_/a_27_47# _0116_ 0
C52372 _0217_ _0902_/a_27_47# 0.03623f
C52373 _0513_/a_384_47# clknet_1_1__leaf__0465_ 0.00123f
C52374 hold65/a_49_47# _0435_ 0
C52375 hold24/a_391_47# net36 0.06102f
C52376 _0080_ net149 0.00389f
C52377 _0715_/a_27_47# _0986_/a_1059_315# 0.00242f
C52378 hold6/a_49_47# _1043_/a_193_47# 0
C52379 _1053_/a_193_47# input12/a_75_212# 0.00485f
C52380 net125 _0463_ 0
C52381 _0179_ _1054_/a_592_47# 0
C52382 net21 _1044_/a_592_47# 0
C52383 _0537_/a_68_297# _0141_ 0
C52384 _0998_/a_27_47# _0998_/a_193_47# 0.96205f
C52385 _0086_ net62 0
C52386 net64 _0988_/a_634_159# 0.02056f
C52387 _0430_ _0988_/a_27_47# 0
C52388 net126 _0547_/a_150_297# 0
C52389 pp[30] _0219_ 0.11643f
C52390 _0108_ hold95/a_391_47# 0
C52391 _1031_/a_381_47# _0339_ 0.00622f
C52392 hold58/a_49_47# comp0.B\[4\] 0.4459f
C52393 _0635_/a_109_297# _0350_ 0
C52394 _1020_/a_891_413# clknet_0__0457_ 0.01081f
C52395 net204 _0208_ 0.08663f
C52396 _0734_/a_47_47# _0370_ 0
C52397 _0199_ _0465_ 0.04277f
C52398 net54 clknet_1_1__leaf__0460_ 0.01004f
C52399 net119 _0132_ 0
C52400 _0443_ _0640_/a_465_297# 0.00152f
C52401 _0779_/a_510_47# _0395_ 0.00182f
C52402 _1001_/a_466_413# _0350_ 0
C52403 net44 _1012_/a_27_47# 0
C52404 _1046_/a_466_413# _1046_/a_561_413# 0.00772f
C52405 _1046_/a_634_159# _1046_/a_975_413# 0
C52406 net245 net5 0
C52407 _1019_/a_27_47# _0099_ 0.00114f
C52408 _0481_ _0487_ 0
C52409 _1056_/a_27_47# _0153_ 0.0118f
C52410 _1032_/a_975_413# clknet_1_0__leaf__0457_ 0
C52411 net64 _0259_ 0
C52412 _0753_/a_465_47# _0225_ 0
C52413 _1051_/a_891_413# _1050_/a_27_47# 0
C52414 _1051_/a_634_159# _1050_/a_466_413# 0
C52415 _1051_/a_1059_315# _1050_/a_193_47# 0.00596f
C52416 _1051_/a_466_413# _1050_/a_634_159# 0
C52417 _1051_/a_27_47# _1050_/a_891_413# 0
C52418 _1051_/a_193_47# _1050_/a_1059_315# 0.00596f
C52419 net45 acc0.A\[17\] 0.08844f
C52420 _0985_/a_193_47# net9 0
C52421 _0985_/a_1059_315# net175 0
C52422 clknet_1_0__leaf__0462_ hold53/a_391_47# 0.01794f
C52423 hold9/a_391_47# _1028_/a_27_47# 0
C52424 _0227_ _0487_ 0
C52425 _0982_/a_193_47# clkbuf_0__0457_/a_110_47# 0
C52426 _0996_/a_592_47# acc0.A\[15\] 0
C52427 hold91/a_285_47# _0301_ 0
C52428 clknet_1_0__leaf__0463_ _1038_/a_561_413# 0
C52429 _0144_ comp0.B\[9\] 0
C52430 net175 _1049_/a_193_47# 0
C52431 _0183_ _0612_/a_145_75# 0
C52432 _0272_ _0840_/a_68_297# 0
C52433 _0998_/a_891_413# clknet_1_1__leaf__0461_ 0
C52434 _0259_ _0423_ 0.034f
C52435 _0289_ _0816_/a_68_297# 0
C52436 _0131_ net17 0
C52437 _0554_/a_68_297# _0474_ 0
C52438 _0775_/a_215_47# _0347_ 0.06136f
C52439 net63 net15 0
C52440 _0457_ _1032_/a_381_47# 0.00422f
C52441 net66 _0186_ 0.02679f
C52442 _1016_/a_891_413# _0218_ 0
C52443 _0179_ hold35/a_285_47# 0
C52444 _1024_/a_193_47# output52/a_27_47# 0
C52445 VPWR _0999_/a_891_413# 0.20666f
C52446 hold27/a_391_47# _0536_/a_149_47# 0
C52447 hold27/a_285_47# _0536_/a_240_47# 0
C52448 _1052_/a_1059_315# acc0.A\[6\] 0.16544f
C52449 _0359_ _0324_ 0.65128f
C52450 _1052_/a_193_47# net13 0
C52451 _0614_/a_111_297# _0352_ 0
C52452 _0501_/a_27_47# control0.reset 0.18342f
C52453 _0983_/a_1059_315# net165 0
C52454 net45 net60 0.17859f
C52455 _0230_ acc0.A\[21\] 0
C52456 _0226_ _0227_ 0.13671f
C52457 _0316_ _0690_/a_150_297# 0
C52458 acc0.A\[4\] net62 0.32681f
C52459 _0697_/a_80_21# clkbuf_1_1__f__0460_/a_110_47# 0
C52460 _0464_ net20 0
C52461 _0344_ _0195_ 0.09394f
C52462 _0985_/a_975_413# _0083_ 0
C52463 _0984_/a_193_47# net58 0.00109f
C52464 _0240_ _0306_ 0.04335f
C52465 _0924_/a_27_47# acc0.A\[15\] 0.02567f
C52466 _0172_ _0542_/a_51_297# 0.15185f
C52467 net36 net100 0.0181f
C52468 _0369_ _0306_ 0
C52469 _0463_ _0473_ 0.06831f
C52470 clkbuf_0__0463_/a_110_47# _0475_ 0
C52471 _0985_/a_634_159# acc0.A\[3\] 0
C52472 _0346_ _1014_/a_193_47# 0.00663f
C52473 clknet_1_0__leaf__0460_ net90 0.09783f
C52474 _0302_ _0219_ 0
C52475 _0970_/a_114_47# _0162_ 0.00429f
C52476 _0299_ _0409_ 0.00779f
C52477 net216 _0245_ 0
C52478 output45/a_27_47# _0708_/a_68_297# 0.00128f
C52479 _1053_/a_891_413# net15 0.00133f
C52480 _1053_/a_466_413# _0191_ 0
C52481 hold101/a_391_47# _0346_ 0.06732f
C52482 _0982_/a_466_413# _0080_ 0.00648f
C52483 _0982_/a_1059_315# net68 0
C52484 hold88/a_49_47# net235 0
C52485 _1049_/a_634_159# _0147_ 0.04169f
C52486 _1049_/a_466_413# net135 0
C52487 clknet_1_1__leaf__0459_ _0653_/a_113_47# 0
C52488 clkbuf_0__0465_/a_110_47# _0218_ 0
C52489 _0459_ clkbuf_1_0__f__0461_/a_110_47# 0.00338f
C52490 hold25/a_49_47# _1040_/a_27_47# 0
C52491 _1011_/a_27_47# hold80/a_49_47# 0
C52492 net12 net13 0.03807f
C52493 _0172_ _0142_ 0.17044f
C52494 _0226_ _0759_/a_113_47# 0
C52495 _0747_/a_297_297# net216 0.00359f
C52496 _0747_/a_79_21# _0371_ 0.12457f
C52497 hold96/a_285_47# _0576_/a_27_297# 0
C52498 _0598_/a_382_297# hold3/a_49_47# 0
C52499 _0985_/a_466_413# _0504_/a_27_47# 0
C52500 _0606_/a_215_297# _0606_/a_392_297# 0.00419f
C52501 _0606_/a_109_53# _0606_/a_297_297# 0
C52502 _0473_ _1044_/a_1059_315# 0
C52503 _0748_/a_81_21# _0350_ 0
C52504 VPWR _0530_/a_299_297# 0.2927f
C52505 _1070_/a_634_159# _1070_/a_466_413# 0.23992f
C52506 _1070_/a_193_47# _1070_/a_1059_315# 0.03405f
C52507 _1070_/a_27_47# _1070_/a_891_413# 0.03224f
C52508 _1052_/a_891_413# _0523_/a_299_297# 0
C52509 _0399_ _0084_ 0.18304f
C52510 _1053_/a_1059_315# _1053_/a_891_413# 0.31086f
C52511 _1053_/a_193_47# _1053_/a_975_413# 0
C52512 _1053_/a_466_413# _1053_/a_381_47# 0.03733f
C52513 _0575_/a_27_297# net199 0.11535f
C52514 hold42/a_49_47# acc0.A\[10\] 0
C52515 net44 _1030_/a_27_47# 0.08503f
C52516 _0268_ _0267_ 0.00877f
C52517 _0647_/a_47_47# _0647_/a_129_47# 0.00369f
C52518 net169 A[8] 0
C52519 _1057_/a_466_413# acc0.A\[10\] 0.00612f
C52520 clknet_1_0__leaf__0465_ _1050_/a_466_413# 0.00207f
C52521 _1015_/a_27_47# net118 0
C52522 _0578_/a_109_47# net23 0
C52523 _0180_ clknet_1_1__leaf__0458_ 0.08132f
C52524 _0329_ _1010_/a_891_413# 0
C52525 net45 _0998_/a_634_159# 0.00431f
C52526 _0217_ _1023_/a_193_47# 0
C52527 acc0.A\[22\] _1023_/a_27_47# 0
C52528 _0198_ _1061_/a_27_47# 0.00139f
C52529 _1032_/a_27_47# _0208_ 0
C52530 net186 _1065_/a_193_47# 0
C52531 hold43/a_49_47# _0195_ 0
C52532 _1066_/a_466_413# clknet_1_1__leaf_clk 0
C52533 _0186_ _0350_ 0
C52534 _0238_ net51 0
C52535 _0253_ acc0.A\[8\] 0.075f
C52536 hold75/a_49_47# acc0.A\[15\] 0.00511f
C52537 _0339_ _0219_ 0.06083f
C52538 _0314_ _1007_/a_466_413# 0
C52539 _1037_/a_1059_315# _0176_ 0
C52540 hold64/a_285_47# net36 0
C52541 _1034_/a_891_413# _0175_ 0
C52542 hold32/a_285_47# clknet_1_1__leaf__0465_ 0.00162f
C52543 net21 _1042_/a_1059_315# 0
C52544 net58 clkbuf_0__0458_/a_110_47# 0.00994f
C52545 acc0.A\[23\] _1022_/a_27_47# 0
C52546 _1068_/a_634_159# _0166_ 0.00105f
C52547 _0401_ _0420_ 0
C52548 _1030_/a_634_159# _1030_/a_592_47# 0
C52549 clkbuf_1_1__f__0464_/a_110_47# _1044_/a_1059_315# 0.02112f
C52550 _1038_/a_193_47# _0552_/a_68_297# 0
C52551 _0200_ _1045_/a_891_413# 0
C52552 clknet_1_0__leaf__0458_ _0631_/a_109_297# 0
C52553 clkbuf_1_1__f__0463_/a_110_47# _0494_/a_27_47# 0
C52554 clknet_1_0__leaf__0462_ _0758_/a_79_21# 0.00367f
C52555 _0270_ _0271_ 0.0993f
C52556 _0476_ _0470_ 0
C52557 _0234_ _0225_ 0.67309f
C52558 _0432_ clknet_1_1__leaf__0458_ 0.24992f
C52559 hold27/a_285_47# _1046_/a_27_47# 0
C52560 hold27/a_49_47# _1046_/a_193_47# 0
C52561 _0251_ _0152_ 0
C52562 _1014_/a_1059_315# hold60/a_49_47# 0.00621f
C52563 acc0.A\[12\] _0808_/a_266_47# 0
C52564 net148 _0150_ 0
C52565 _0621_/a_35_297# _0186_ 0
C52566 _0764_/a_81_21# _0345_ 0
C52567 _1035_/a_592_47# net122 0
C52568 _0992_/a_561_413# net37 0
C52569 clknet_0__0463_ _0913_/a_27_47# 0.03152f
C52570 _0343_ net46 0.05249f
C52571 net21 net10 0.0246f
C52572 _0389_ acc0.A\[19\] 0.06137f
C52573 net122 B[15] 0.01215f
C52574 _0458_ _0639_/a_109_297# 0
C52575 _0598_/a_297_47# _0230_ 0.00119f
C52576 _1015_/a_592_47# _0181_ 0
C52577 output49/a_27_47# net49 0.21914f
C52578 _0987_/a_634_159# _0987_/a_381_47# 0
C52579 _0349_ acc0.A\[29\] 0.02672f
C52580 _0151_ _0191_ 0.00164f
C52581 net194 _1051_/a_1059_315# 0
C52582 _0354_ _0333_ 0.36683f
C52583 acc0.A\[27\] _0318_ 0.38802f
C52584 _0149_ _0186_ 0.16279f
C52585 _0263_ net218 0.00139f
C52586 clknet_0__0462_ _0350_ 0
C52587 hold49/a_49_47# _1044_/a_1059_315# 0
C52588 net194 _1045_/a_381_47# 0
C52589 _0182_ _1047_/a_193_47# 0.01778f
C52590 _0180_ _1047_/a_27_47# 0.00321f
C52591 acc0.A\[1\] _1047_/a_634_159# 0
C52592 _0713_/a_27_47# hold40/a_391_47# 0
C52593 _0608_/a_109_297# _0308_ 0
C52594 acc0.A\[20\] _0765_/a_215_47# 0.03909f
C52595 _0992_/a_592_47# net67 0
C52596 clknet_1_0__leaf__0465_ _0518_/a_373_47# 0
C52597 _1000_/a_592_47# VPWR 0
C52598 _1004_/a_27_47# _1004_/a_891_413# 0.03206f
C52599 _1004_/a_193_47# _1004_/a_1059_315# 0.03405f
C52600 _1004_/a_634_159# _1004_/a_466_413# 0.23992f
C52601 net126 net153 0
C52602 _0342_ _0778_/a_68_297# 0
C52603 _0129_ _0338_ 0
C52604 _1027_/a_27_47# _1008_/a_27_47# 0
C52605 _0410_ net41 0.44417f
C52606 _0151_ _1053_/a_381_47# 0.11656f
C52607 clkload4/a_268_47# acc0.A\[16\] 0
C52608 _0486_ clknet_0_clk 0.07416f
C52609 _1059_/a_27_47# _1060_/a_891_413# 0
C52610 _0967_/a_109_93# _0477_ 0.01427f
C52611 _0476_ _0958_/a_303_47# 0.00527f
C52612 _0219_ net6 0.32953f
C52613 _0477_ _0487_ 0
C52614 rst _1064_/a_27_47# 0
C52615 pp[29] _0703_/a_109_297# 0.00238f
C52616 _0633_/a_109_297# _0264_ 0
C52617 _1029_/a_634_159# _1029_/a_381_47# 0
C52618 hold75/a_49_47# _0179_ 0
C52619 net40 output45/a_27_47# 0
C52620 _0462_ hold73/a_285_47# 0.01643f
C52621 hold37/a_285_47# _1045_/a_27_47# 0.00104f
C52622 _0352_ net223 0.28799f
C52623 VPWR _0565_/a_149_47# 0
C52624 _0389_ _0249_ 0
C52625 comp0.B\[15\] _0499_/a_145_75# 0
C52626 _0447_ _0219_ 0.12594f
C52627 _0195_ _0997_/a_27_47# 0
C52628 _0136_ A[1] 0
C52629 _0318_ _0364_ 0
C52630 clkbuf_1_1__f__0460_/a_110_47# _0345_ 0
C52631 acc0.A\[12\] _0345_ 0.07417f
C52632 clkbuf_1_0__f__0464_/a_110_47# net132 0
C52633 net4 clknet_1_1__leaf__0465_ 0.1687f
C52634 VPWR clkbuf_1_1__f__0462_/a_110_47# 1.32032f
C52635 clkload0/a_27_47# _1072_/a_891_413# 0.0041f
C52636 clkload0/X _1072_/a_27_47# 0
C52637 net64 _0253_ 0.20419f
C52638 _0275_ clkbuf_1_1__f__0465_/a_110_47# 0.00449f
C52639 comp0.B\[15\] net149 0
C52640 _0621_/a_117_297# _0253_ 0.00127f
C52641 acc0.A\[4\] _0987_/a_634_159# 0.01978f
C52642 net213 _0754_/a_51_297# 0
C52643 _0359_ _0347_ 0
C52644 net35 _0468_ 0.16918f
C52645 net103 _1016_/a_27_47# 0.02985f
C52646 _0661_/a_205_297# _0289_ 0.00311f
C52647 _0661_/a_27_297# _0293_ 0.10108f
C52648 net178 net16 0.04042f
C52649 _0661_/a_109_297# _0287_ 0.0013f
C52650 _0760_/a_285_47# net51 0
C52651 acc0.A\[8\] net74 0
C52652 _0346_ _0369_ 0.04054f
C52653 _0272_ _0255_ 0.00135f
C52654 _0222_ hold4/a_49_47# 0.03345f
C52655 control0.count\[3\] _1068_/a_193_47# 0
C52656 clknet_0__0457_ _0346_ 0.55558f
C52657 _1037_/a_975_413# clknet_1_1__leaf__0463_ 0
C52658 _0378_ _1023_/a_466_413# 0
C52659 hold81/a_49_47# hold81/a_285_47# 0.22264f
C52660 _0555_/a_245_297# net204 0
C52661 _1028_/a_193_47# _1028_/a_381_47# 0.09799f
C52662 _1028_/a_634_159# _1028_/a_891_413# 0.03684f
C52663 _1028_/a_27_47# _1028_/a_561_413# 0.00163f
C52664 hold41/a_391_47# hold42/a_391_47# 0.0141f
C52665 _0180_ clknet_1_0__leaf__0461_ 0
C52666 net118 _0215_ 0
C52667 _0343_ _0996_/a_27_47# 0.0043f
C52668 net65 _0369_ 0.1433f
C52669 _0369_ _0989_/a_466_413# 0.0023f
C52670 _0266_ net165 0.11014f
C52671 _0441_ _0835_/a_292_297# 0.00105f
C52672 _0837_/a_368_297# _0255_ 0
C52673 _0440_ _0835_/a_493_297# 0
C52674 _0442_ _0835_/a_78_199# 0
C52675 _0115_ hold72/a_285_47# 0.00704f
C52676 _0216_ hold60/a_391_47# 0
C52677 _0394_ _1009_/a_891_413# 0
C52678 _1033_/a_891_413# comp0.B\[1\] 0.00363f
C52679 _0369_ _0992_/a_466_413# 0.00147f
C52680 _0852_/a_117_297# _0346_ 0.00409f
C52681 _0985_/a_561_413# VPWR 0.0032f
C52682 hold27/a_49_47# comp0.B\[9\] 0
C52683 pp[30] hold61/a_49_47# 0.00818f
C52684 _0445_ _0345_ 0.00425f
C52685 control0.count\[3\] _0478_ 0.29879f
C52686 acc0.A\[8\] output61/a_27_47# 0
C52687 VPWR _1018_/a_381_47# 0.07101f
C52688 clknet_1_1__leaf__0459_ _0651_/a_113_47# 0
C52689 A[13] pp[14] 0.0151f
C52690 clknet_1_1__leaf__0460_ net227 0.00293f
C52691 clknet_0__0463_ _0172_ 0.005f
C52692 net10 _0261_ 0.00102f
C52693 VPWR _1049_/a_1059_315# 0.39863f
C52694 _0179_ _0516_/a_109_297# 0
C52695 _0743_/a_240_47# _0367_ 0.01379f
C52696 net200 _0347_ 0
C52697 _0812_/a_79_21# net228 0
C52698 _0100_ hold93/a_391_47# 0
C52699 _1041_/a_634_159# net31 0.0402f
C52700 _0575_/a_27_297# VPWR 0.20197f
C52701 _0376_ net46 0
C52702 _0693_/a_68_297# _0250_ 0
C52703 hold97/a_391_47# _1008_/a_27_47# 0
C52704 hold97/a_285_47# _1008_/a_193_47# 0.01463f
C52705 VPWR _1066_/a_1059_315# 0.42725f
C52706 net136 acc0.A\[4\] 0.09414f
C52707 _0981_/a_27_297# _0480_ 0
C52708 _0266_ acc0.A\[19\] 0
C52709 _0650_/a_68_297# _0345_ 0
C52710 VPWR _1068_/a_1059_315# 0.37998f
C52711 net179 acc0.A\[9\] 0
C52712 VPWR A[0] 0.4056f
C52713 _0455_ _0853_/a_68_297# 0.10689f
C52714 _0454_ _0853_/a_150_297# 0
C52715 VPWR acc0.A\[17\] 0.83381f
C52716 hold13/a_285_47# _0463_ 0
C52717 _0337_ _0353_ 0
C52718 comp0.B\[14\] _1044_/a_27_47# 0
C52719 _0241_ _0350_ 0
C52720 _0277_ _0406_ 0
C52721 _1051_/a_891_413# _0987_/a_27_47# 0.00302f
C52722 net101 clkbuf_1_1__f__0457_/a_110_47# 0
C52723 VPWR net18 0.71609f
C52724 _0993_/a_27_47# _0091_ 0.11455f
C52725 _0993_/a_634_159# _0419_ 0.00194f
C52726 _0993_/a_1059_315# _0417_ 0
C52727 _0518_/a_109_297# acc0.A\[8\] 0.0015f
C52728 _0828_/a_113_297# _0436_ 0.09847f
C52729 _0828_/a_199_47# _0435_ 0
C52730 net1 _1015_/a_193_47# 0.01349f
C52731 hold32/a_49_47# A[9] 0.02997f
C52732 _0140_ _1043_/a_1059_315# 0
C52733 net198 _1043_/a_975_413# 0
C52734 net18 _1043_/a_561_413# 0.00133f
C52735 hold76/a_49_47# _0771_/a_215_297# 0.01107f
C52736 hold76/a_285_47# _0771_/a_27_413# 0.00495f
C52737 _0642_/a_382_47# acc0.A\[8\] 0
C52738 clknet_1_0__leaf__0465_ _1046_/a_1059_315# 0.00177f
C52739 _0465_ _0449_ 0.00851f
C52740 _0531_/a_27_297# net9 0.17238f
C52741 _0170_ _1071_/a_466_413# 0
C52742 _1016_/a_193_47# net219 0
C52743 hold25/a_49_47# net171 0.09036f
C52744 net187 clknet_1_0__leaf__0457_ 0.066f
C52745 _0136_ clkbuf_0__0463_/a_110_47# 0
C52746 clkbuf_1_0__f_clk/a_110_47# _1068_/a_27_47# 0
C52747 _0227_ _0760_/a_47_47# 0
C52748 acc0.A\[21\] _0760_/a_377_297# 0
C52749 _0662_/a_81_21# acc0.A\[9\] 0.01868f
C52750 _0710_/a_109_297# _0220_ 0.01051f
C52751 net45 _0793_/a_245_297# 0
C52752 _1019_/a_466_413# clkbuf_0__0457_/a_110_47# 0.00789f
C52753 _0998_/a_466_413# _0998_/a_592_47# 0.00553f
C52754 _0998_/a_634_159# _0998_/a_1017_47# 0
C52755 _0803_/a_68_297# _0403_ 0.00594f
C52756 _1009_/a_634_159# _0318_ 0
C52757 net64 net74 0.00523f
C52758 clknet_1_1__leaf__0459_ _0806_/a_199_47# 0
C52759 _0621_/a_117_297# net74 0.00129f
C52760 net10 _0509_/a_27_47# 0
C52761 _0101_ _0762_/a_79_21# 0.05937f
C52762 net247 _1061_/a_27_47# 0
C52763 _1024_/a_466_413# acc0.A\[23\] 0
C52764 VPWR net60 1.06863f
C52765 net203 _1033_/a_27_47# 0.03047f
C52766 hold56/a_285_47# _1033_/a_381_47# 0
C52767 _0404_ _0788_/a_150_297# 0
C52768 _0984_/a_27_47# net47 0.03082f
C52769 _0282_ hold81/a_49_47# 0.00222f
C52770 _0346_ _0844_/a_79_21# 0
C52771 hold38/a_49_47# comp0.B\[6\] 0
C52772 hold38/a_285_47# comp0.B\[5\] 0
C52773 VPWR net5 0.84437f
C52774 _1019_/a_193_47# _1019_/a_592_47# 0.00135f
C52775 _1019_/a_466_413# _1019_/a_561_413# 0.00772f
C52776 _1019_/a_634_159# _1019_/a_975_413# 0
C52777 _1058_/a_193_47# net37 0.01203f
C52778 _0123_ _0574_/a_27_297# 0.11026f
C52779 _0347_ net228 0.02644f
C52780 hold42/a_49_47# _0188_ 0.02283f
C52781 _1057_/a_466_413# _0188_ 0
C52782 clknet_1_1__leaf__0463_ _0959_/a_80_21# 0
C52783 hold89/a_49_47# _0946_/a_30_53# 0.04532f
C52784 _0469_ clkbuf_0_clk/a_110_47# 0.00716f
C52785 _0420_ hold70/a_49_47# 0
C52786 clknet_1_1__leaf__0458_ _0986_/a_381_47# 0
C52787 net72 _0986_/a_1059_315# 0
C52788 net133 _0180_ 0.08945f
C52789 VPWR _1012_/a_561_413# 0.00372f
C52790 net133 net218 0
C52791 hold54/a_285_47# _0208_ 0.03742f
C52792 net22 _0545_/a_68_297# 0.0248f
C52793 _0398_ _0307_ 0.17362f
C52794 _0849_/a_79_21# net146 0
C52795 net55 _0316_ 0.08028f
C52796 net64 output61/a_27_47# 0.00103f
C52797 _0472_ _0176_ 0.04124f
C52798 _0726_/a_51_297# _0726_/a_149_47# 0.02487f
C52799 _1050_/a_1059_315# net184 0
C52800 _1050_/a_891_413# net131 0
C52801 acc0.A\[4\] _1045_/a_193_47# 0
C52802 _0217_ hold2/a_285_47# 0
C52803 net59 clknet_1_1__leaf__0462_ 0.10199f
C52804 hold9/a_49_47# net114 0.0028f
C52805 net66 net62 0
C52806 _1058_/a_466_413# net67 0.00975f
C52807 _1013_/a_27_47# _0220_ 0
C52808 _0325_ _0324_ 0.20844f
C52809 clknet_1_0__leaf__0458_ _1060_/a_27_47# 0
C52810 hold55/a_49_47# _1032_/a_27_47# 0.00166f
C52811 _0717_/a_80_21# hold61/a_49_47# 0
C52812 net55 _0347_ 0.0441f
C52813 control0.sh net201 0.00757f
C52814 _0718_/a_285_47# hold16/a_285_47# 0
C52815 _1050_/a_27_47# _0528_/a_81_21# 0
C52816 clknet_1_0__leaf__0465_ _0270_ 0
C52817 hold26/a_49_47# net22 0.04546f
C52818 _0982_/a_193_47# _0350_ 0
C52819 _0182_ _0585_/a_109_297# 0
C52820 _0180_ _0585_/a_27_297# 0
C52821 net162 _1031_/a_891_413# 0.00413f
C52822 _0629_/a_59_75# _0844_/a_79_21# 0.00355f
C52823 VPWR _0998_/a_634_159# 0.18061f
C52824 hold3/a_285_47# hold3/a_391_47# 0.41909f
C52825 net149 hold71/a_285_47# 0
C52826 _0335_ hold61/a_391_47# 0
C52827 _0338_ hold61/a_285_47# 0.05758f
C52828 clknet_1_0__leaf__0465_ _0987_/a_466_413# 0.00559f
C52829 clknet_1_0__leaf__0463_ _0545_/a_68_297# 0
C52830 _0991_/a_27_47# _0450_ 0
C52831 _0991_/a_193_47# _0446_ 0
C52832 _0758_/a_297_297# _0102_ 0
C52833 _0758_/a_215_47# _0352_ 0.00137f
C52834 _1024_/a_592_47# net52 0
C52835 _0991_/a_1059_315# _0218_ 0
C52836 _0294_ _0991_/a_891_413# 0.02199f
C52837 _0990_/a_634_159# _0990_/a_592_47# 0
C52838 _0461_ _0771_/a_298_297# 0
C52839 net50 _0374_ 0
C52840 net42 _0345_ 0.18086f
C52841 _0790_/a_285_297# _0219_ 0.00352f
C52842 _0267_ net222 0
C52843 _0546_/a_51_297# net127 0
C52844 _1002_/a_466_413# _0460_ 0.00998f
C52845 _1002_/a_891_413# clknet_1_0__leaf__0457_ 0.00179f
C52846 net46 _0224_ 0
C52847 net168 _0152_ 0.01847f
C52848 _0949_/a_59_75# _0958_/a_27_47# 0.01546f
C52849 _0430_ _0642_/a_215_297# 0.01553f
C52850 _0537_/a_68_297# _1043_/a_27_47# 0
C52851 clknet_1_0__leaf__0463_ hold26/a_49_47# 0
C52852 _0179_ net71 0.06884f
C52853 _0556_/a_68_297# _1035_/a_27_47# 0
C52854 _0304_ acc0.A\[15\] 0.08007f
C52855 _0174_ _0205_ 0.18223f
C52856 _0564_/a_68_297# _0564_/a_150_297# 0.00477f
C52857 _0433_ _0436_ 0
C52858 _0476_ _0485_ 0.11529f
C52859 hold49/a_391_47# _0176_ 0.00299f
C52860 _1065_/a_27_47# _0951_/a_109_93# 0.0014f
C52861 _0393_ _0774_/a_150_297# 0
C52862 _0488_ control0.state\[2\] 0
C52863 hold24/a_391_47# _1039_/a_27_47# 0
C52864 comp0.B\[10\] net152 0.13959f
C52865 _0251_ net248 0
C52866 hold66/a_285_47# clknet_1_0__leaf__0460_ 0.01605f
C52867 net200 _1025_/a_27_47# 0.09285f
C52868 _0216_ net113 0.1917f
C52869 net135 _0147_ 0
C52870 _0743_/a_51_297# _0319_ 0
C52871 net62 _0350_ 0.50872f
C52872 hold9/a_49_47# _0365_ 0
C52873 _1051_/a_27_47# _1051_/a_634_159# 0.14145f
C52874 _0450_ _0350_ 0.08276f
C52875 VPWR acc0.A\[11\] 1.44211f
C52876 _0083_ _0504_/a_27_47# 0
C52877 _0606_/a_465_297# _0236_ 0
C52878 _0612_/a_59_75# acc0.A\[19\] 0
C52879 _1070_/a_634_159# _0168_ 0.00281f
C52880 _1070_/a_1059_315# VPWR 0.4108f
C52881 net106 _1033_/a_634_159# 0
C52882 _0226_ _0352_ 0
C52883 _1045_/a_634_159# _1045_/a_1059_315# 0
C52884 _1045_/a_27_47# _1045_/a_381_47# 0.06222f
C52885 _1045_/a_193_47# _1045_/a_891_413# 0.19685f
C52886 net189 acc0.A\[10\] 0.02826f
C52887 net45 net84 0.00433f
C52888 net150 net109 0
C52889 clknet_1_0__leaf__0462_ hold30/a_391_47# 0.01705f
C52890 net157 net201 0
C52891 _1066_/a_1017_47# control0.sh 0
C52892 _1014_/a_561_413# _0465_ 0
C52893 _0552_/a_68_297# net29 0.02257f
C52894 _1062_/a_561_413# _0468_ 0
C52895 _0473_ clkbuf_1_0__f__0463_/a_110_47# 0.03777f
C52896 VPWR _1030_/a_561_413# 0.00306f
C52897 clknet_1_1__leaf__0463_ _0173_ 0.49414f
C52898 _0314_ _0105_ 0.0451f
C52899 _0783_/a_297_297# _0397_ 0
C52900 _1029_/a_27_47# _0365_ 0
C52901 _0378_ net241 0
C52902 _0733_/a_79_199# _0697_/a_80_21# 0.0013f
C52903 _1043_/a_634_159# _1043_/a_1059_315# 0
C52904 _1043_/a_27_47# _1043_/a_381_47# 0.06222f
C52905 _1043_/a_193_47# _1043_/a_891_413# 0.19489f
C52906 clknet_1_0__leaf__0459_ acc0.A\[17\] 0.00163f
C52907 net177 net151 0
C52908 _0372_ _0345_ 0.14736f
C52909 _0654_/a_27_413# acc0.A\[11\] 0
C52910 _1038_/a_891_413# _0209_ 0.03377f
C52911 hold52/a_391_47# _0217_ 0
C52912 _1004_/a_1059_315# VPWR 0.40386f
C52913 _1021_/a_466_413# _1002_/a_466_413# 0
C52914 comp0.B\[2\] control0.sh 0
C52915 _0216_ _0720_/a_150_297# 0
C52916 _1021_/a_27_47# _1002_/a_381_47# 0.00112f
C52917 _1021_/a_891_413# _1002_/a_193_47# 0
C52918 hold89/a_391_47# _0484_ 0
C52919 hold89/a_49_47# _0487_ 0.04985f
C52920 _1054_/a_27_47# _1054_/a_193_47# 0.96668f
C52921 _0736_/a_56_297# clknet_1_1__leaf__0460_ 0.0026f
C52922 _1071_/a_27_47# clknet_1_0__leaf_clk 0.23748f
C52923 _0363_ _0181_ 0.11889f
C52924 _0174_ _1042_/a_193_47# 0.00433f
C52925 acc0.A\[14\] _0269_ 0.1477f
C52926 hold65/a_391_47# acc0.A\[6\] 0.02811f
C52927 _0783_/a_79_21# acc0.A\[17\] 0
C52928 net8 _0173_ 0
C52929 _1032_/a_1017_47# net17 0.00117f
C52930 _0227_ _0350_ 0
C52931 hold28/a_391_47# _0180_ 0.00673f
C52932 comp0.B\[10\] _1042_/a_466_413# 0
C52933 _0425_ _0218_ 0
C52934 net194 _1044_/a_891_413# 0
C52935 hold28/a_391_47# net218 0
C52936 _0792_/a_80_21# _0792_/a_209_297# 0.06257f
C52937 _0467_ _0466_ 0.11899f
C52938 _0987_/a_891_413# _0085_ 0.05681f
C52939 _0987_/a_381_47# net73 0
C52940 _0241_ _0244_ 0.00403f
C52941 A[4] A[5] 0.21305f
C52942 net53 _0697_/a_80_21# 0
C52943 control0.state\[2\] _1064_/a_27_47# 0
C52944 input4/a_75_212# acc0.A\[11\] 0
C52945 _0219_ _0685_/a_150_297# 0
C52946 _0823_/a_109_297# _0431_ 0.01129f
C52947 _0207_ net28 0
C52948 VPWR hold81/a_391_47# 0.18794f
C52949 _0972_/a_93_21# _0471_ 0.08492f
C52950 _0343_ _0794_/a_27_47# 0
C52951 clknet_0__0461_ _0775_/a_79_21# 0.00126f
C52952 clknet_1_0__leaf__0459_ net5 0.05387f
C52953 _0352_ clkbuf_0__0457_/a_110_47# 0
C52954 _0134_ _1035_/a_27_47# 0
C52955 _0557_/a_51_297# net121 0
C52956 hold47/a_285_47# _0196_ 0
C52957 _0642_/a_27_413# _0432_ 0
C52958 hold78/a_49_47# acc0.A\[31\] 0.01553f
C52959 _1059_/a_634_159# _0158_ 0
C52960 net145 _1060_/a_466_413# 0
C52961 _0983_/a_193_47# _0983_/a_466_413# 0.08015f
C52962 _0983_/a_27_47# _0983_/a_1059_315# 0.04875f
C52963 _0820_/a_79_21# hold67/a_49_47# 0.00163f
C52964 pp[17] output45/a_27_47# 0
C52965 hold34/a_285_47# net16 0
C52966 clknet_1_0__leaf__0465_ _1051_/a_27_47# 0.01151f
C52967 net224 clknet_1_1__leaf__0460_ 0.02621f
C52968 clknet_1_0__leaf__0465_ _1045_/a_634_159# 0.00208f
C52969 _1029_/a_381_47# net115 0
C52970 _1029_/a_891_413# net191 0
C52971 hold98/a_49_47# _0995_/a_193_47# 0.00405f
C52972 hold98/a_285_47# _0995_/a_27_47# 0
C52973 _0201_ _0954_/a_32_297# 0.06524f
C52974 _0538_/a_51_297# comp0.B\[12\] 0
C52975 _0399_ _0507_/a_27_297# 0
C52976 _0325_ _0347_ 0
C52977 _0258_ _0825_/a_68_297# 0.17674f
C52978 _0183_ clknet_1_0__leaf__0460_ 0.02346f
C52979 _0770_/a_79_21# VPWR 0.27636f
C52980 net55 hold95/a_49_47# 0.00832f
C52981 _0769_/a_81_21# _0391_ 0.00144f
C52982 _0244_ _0772_/a_510_47# 0
C52983 VPWR net175 0.30365f
C52984 net236 _0467_ 0
C52985 _0180_ _0218_ 0.00194f
C52986 clknet_1_0__leaf__0462_ _0574_/a_373_47# 0.00141f
C52987 _1015_/a_27_47# _0526_/a_27_47# 0
C52988 _0346_ _0409_ 0.01344f
C52989 net213 _0219_ 0
C52990 acc0.A\[4\] net73 0
C52991 _0399_ net165 0.044f
C52992 net39 _0301_ 0
C52993 _0113_ _0565_/a_149_47# 0
C52994 acc0.A\[10\] _0417_ 0
C52995 clknet_0__0465_ _0256_ 0
C52996 _1020_/a_381_47# _0183_ 0
C52997 _1003_/a_27_47# _0217_ 0.00413f
C52998 _0956_/a_32_297# _0956_/a_114_297# 0.01439f
C52999 net216 _0326_ 0.00347f
C53000 _0806_/a_113_297# _0418_ 0.09755f
C53001 acc0.A\[31\] _0129_ 0.00347f
C53002 _1013_/a_193_47# _0218_ 0.026f
C53003 _0854_/a_510_47# clknet_1_0__leaf__0461_ 0
C53004 _1016_/a_1059_315# _1016_/a_891_413# 0.31086f
C53005 _1016_/a_193_47# _1016_/a_975_413# 0
C53006 _1016_/a_466_413# _1016_/a_381_47# 0.03733f
C53007 hold25/a_285_47# _1037_/a_634_159# 0
C53008 _0138_ _1061_/a_193_47# 0
C53009 _0331_ _0698_/a_199_47# 0
C53010 _0699_/a_150_297# _0330_ 0.0015f
C53011 VPWR _0726_/a_149_47# 0
C53012 hold54/a_391_47# _0178_ 0
C53013 net59 hold92/a_49_47# 0.34696f
C53014 _0378_ net177 0
C53015 net61 acc0.A\[8\] 0.02461f
C53016 comp0.B\[1\] _0956_/a_32_297# 0.08749f
C53017 _1028_/a_193_47# acc0.A\[28\] 0.00581f
C53018 control0.count\[2\] _1070_/a_27_47# 0
C53019 hold31/a_391_47# _0252_ 0.00603f
C53020 _0260_ _0465_ 0.01959f
C53021 hold87/a_391_47# _0982_/a_1059_315# 0
C53022 _0228_ _0486_ 0
C53023 _0432_ _0218_ 0.30011f
C53024 clknet_1_1__leaf__0459_ _0407_ 0
C53025 hold42/a_285_47# _0187_ 0
C53026 _1067_/a_381_47# control0.reset 0
C53027 _0213_ _0560_/a_68_297# 0.10609f
C53028 _1057_/a_1059_315# _0187_ 0.05792f
C53029 _0812_/a_215_47# _0422_ 0.00754f
C53030 _0812_/a_79_21# _0090_ 0.05046f
C53031 _0812_/a_510_47# net217 0
C53032 _0399_ acc0.A\[19\] 0.03062f
C53033 _0462_ clknet_0__0460_ 0.064f
C53034 _0385_ _0460_ 0.01513f
C53035 VPWR _0990_/a_561_413# 0.00262f
C53036 _0999_/a_381_47# _0096_ 0
C53037 VPWR _0793_/a_245_297# 0.00493f
C53038 hold44/a_285_47# hold50/a_49_47# 0
C53039 _0733_/a_79_199# _0345_ 0
C53040 _0397_ _0777_/a_47_47# 0.03108f
C53041 net39 _0994_/a_193_47# 0.16683f
C53042 pp[9] net37 0.0135f
C53043 acc0.A\[16\] hold19/a_391_47# 0.05073f
C53044 _0107_ _0780_/a_117_297# 0
C53045 _1059_/a_634_159# acc0.A\[14\] 0.04694f
C53046 _1041_/a_634_159# net7 0.01682f
C53047 _0554_/a_68_297# _1035_/a_27_47# 0
C53048 _0238_ _0104_ 0
C53049 _0313_ _0690_/a_68_297# 0
C53050 hold4/a_391_47# _1022_/a_193_47# 0.00283f
C53051 hold4/a_285_47# _1022_/a_634_159# 0.01163f
C53052 _0460_ _1006_/a_1017_47# 0
C53053 _0984_/a_27_47# _0294_ 0
C53054 _0742_/a_384_47# net52 0
C53055 _0143_ clknet_1_1__leaf__0464_ 0.19993f
C53056 _0198_ _1047_/a_634_159# 0
C53057 _0490_ _0169_ 0
C53058 _0170_ _0480_ 0.0023f
C53059 _1056_/a_193_47# input16/a_75_212# 0
C53060 _0764_/a_384_47# _0346_ 0
C53061 _0170_ _1072_/a_891_413# 0
C53062 _0753_/a_79_21# _0754_/a_240_47# 0
C53063 hold27/a_285_47# hold27/a_391_47# 0.41909f
C53064 A[11] _0512_/a_109_47# 0
C53065 _0562_/a_68_297# _0208_ 0
C53066 _0089_ _0267_ 0
C53067 net244 _0345_ 0.05819f
C53068 _0464_ _1049_/a_27_47# 0.00164f
C53069 hold18/a_285_47# _0635_/a_27_47# 0
C53070 hold23/a_49_47# hold23/a_391_47# 0.00188f
C53071 _1054_/a_634_159# VPWR 0.18423f
C53072 _0791_/a_113_297# net42 0
C53073 clknet_1_0__leaf__0462_ _1025_/a_891_413# 0
C53074 net137 _0987_/a_466_413# 0
C53075 _1051_/a_634_159# _0085_ 0
C53076 net231 hold84/a_49_47# 0
C53077 _1056_/a_561_413# VPWR 0.00292f
C53078 _0379_ net52 0
C53079 VPWR _0303_ 0.34647f
C53080 net53 _0345_ 0.08694f
C53081 _0770_/a_297_47# _0389_ 0.05126f
C53082 _0770_/a_79_21# _0390_ 0.12893f
C53083 _0770_/a_382_297# _0243_ 0
C53084 _0283_ acc0.A\[11\] 0.00238f
C53085 _0216_ hold92/a_391_47# 0.01375f
C53086 _1038_/a_193_47# VPWR 0.29315f
C53087 _0287_ clknet_1_1__leaf__0465_ 0.02454f
C53088 net154 _0524_/a_27_297# 0.01598f
C53089 _1041_/a_193_47# A[15] 0.00145f
C53090 _0372_ net52 0
C53091 hold77/a_285_47# _0317_ 0
C53092 _0713_/a_27_47# net1 0.0016f
C53093 _0268_ _0347_ 0
C53094 _0312_ _0368_ 0.01982f
C53095 _0767_/a_145_75# _0347_ 0
C53096 _1018_/a_466_413# acc0.A\[18\] 0.02895f
C53097 _0217_ _0576_/a_373_47# 0
C53098 _0183_ _0576_/a_109_297# 0.00919f
C53099 _0292_ _0088_ 0
C53100 hold74/a_49_47# _0219_ 0.0333f
C53101 _0996_/a_1017_47# net5 0
C53102 clknet_0_clk _1068_/a_975_413# 0
C53103 net120 _1065_/a_193_47# 0
C53104 pp[6] pp[2] 0.18013f
C53105 pp[19] VPWR 0.22041f
C53106 net207 clkbuf_0__0457_/a_110_47# 0.0247f
C53107 _0998_/a_1017_47# net84 0
C53108 hold1/a_391_47# net148 0.13588f
C53109 acc0.A\[12\] _0156_ 0.00208f
C53110 _0092_ net80 0.12107f
C53111 _1021_/a_1059_315# net220 0
C53112 _0552_/a_68_297# _0137_ 0
C53113 net206 _0773_/a_35_297# 0
C53114 _0479_ _0168_ 0
C53115 _0122_ acc0.A\[23\] 0
C53116 VPWR _0281_ 1.6476f
C53117 VPWR _0785_/a_81_21# 0.21985f
C53118 _1001_/a_466_413# _0195_ 0
C53119 _1001_/a_193_47# _0216_ 0
C53120 net64 net61 0.01866f
C53121 _0714_/a_51_297# net225 0.15209f
C53122 _0817_/a_81_21# _0346_ 0.21441f
C53123 _0857_/a_27_47# _1067_/a_27_47# 0.01123f
C53124 net35 _1071_/a_466_413# 0.00133f
C53125 net51 _1005_/a_561_413# 0
C53126 net189 _0188_ 0.02428f
C53127 net40 _0297_ 0.37493f
C53128 comp0.B\[13\] _1042_/a_193_47# 0
C53129 net174 _0540_/a_51_297# 0
C53130 _0216_ hold8/a_285_47# 0.01647f
C53131 net155 hold8/a_391_47# 0.1306f
C53132 _0789_/a_75_199# net5 0
C53133 _0172_ net198 0.04648f
C53134 _0353_ _0333_ 0.5067f
C53135 clknet_1_1__leaf__0460_ _0695_/a_80_21# 0.00224f
C53136 clknet_1_0__leaf__0458_ net149 0.03955f
C53137 _1038_/a_27_47# _0550_/a_51_297# 0
C53138 _0782_/a_27_47# _1014_/a_193_47# 0.00184f
C53139 _0082_ _0158_ 0
C53140 _0231_ net50 0
C53141 _0343_ _0995_/a_466_413# 0.00655f
C53142 _1014_/a_1059_315# clknet_1_0__leaf__0461_ 0.00577f
C53143 _0180_ _0177_ 0
C53144 _0575_/a_109_47# net50 0
C53145 _0726_/a_240_47# net227 0.05778f
C53146 _0259_ _0369_ 0
C53147 clknet_0__0461_ _0581_/a_27_297# 0.00128f
C53148 _0654_/a_27_413# _0281_ 0
C53149 _0269_ _0823_/a_109_297# 0
C53150 comp0.B\[1\] _1032_/a_193_47# 0.00114f
C53151 net199 net176 0.00188f
C53152 _0182_ _0178_ 0.55174f
C53153 _0781_/a_150_297# _0459_ 0
C53154 _0161_ _0468_ 0
C53155 net45 _0783_/a_510_47# 0
C53156 net34 _1064_/a_1059_315# 0.08373f
C53157 control0.state\[0\] _1064_/a_381_47# 0
C53158 control0.state\[1\] _1064_/a_891_413# 0
C53159 control0.state\[2\] net33 0
C53160 clknet_1_0__leaf__0465_ A[4] 0
C53161 _0402_ net37 0.00772f
C53162 _0996_/a_891_413# clkbuf_1_1__f__0459_/a_110_47# 0
C53163 _1033_/a_1059_315# clknet_1_1__leaf__0463_ 0
C53164 _0983_/a_27_47# _0266_ 0
C53165 _0130_ _1032_/a_381_47# 0
C53166 _1015_/a_193_47# net157 0
C53167 _0348_ hold61/a_285_47# 0
C53168 hold18/a_285_47# _0850_/a_68_297# 0
C53169 net214 _0179_ 0
C53170 _0237_ _0487_ 0
C53171 _0283_ hold81/a_391_47# 0.02899f
C53172 _0286_ hold81/a_285_47# 0
C53173 _1050_/a_466_413# _0148_ 0.00632f
C53174 hold46/a_391_47# net10 0.04079f
C53175 _1001_/a_891_413# _0247_ 0
C53176 _0430_ net63 0
C53177 _0716_/a_27_47# _0295_ 0
C53178 hold58/a_391_47# net23 0
C53179 _1059_/a_27_47# net228 0
C53180 _0180_ _0112_ 0.00192f
C53181 _0179_ _0515_/a_384_47# 0
C53182 _1001_/a_634_159# _0369_ 0.00667f
C53183 net58 _0447_ 0.17267f
C53184 _0739_/a_79_21# _0365_ 0.14327f
C53185 VPWR net84 0.34573f
C53186 clknet_0__0457_ _1001_/a_634_159# 0
C53187 net71 _0530_/a_384_47# 0
C53188 _0467_ _1065_/a_634_159# 0.01628f
C53189 clknet_1_0__leaf__0465_ _0085_ 0.00787f
C53190 _0195_ _1047_/a_1059_315# 0.03561f
C53191 _0216_ _1047_/a_634_159# 0
C53192 _0346_ _0084_ 0
C53193 _0450_ _0847_/a_109_297# 0.01181f
C53194 hold12/a_285_47# _0486_ 0
C53195 _0732_/a_80_21# _0743_/a_51_297# 0.0132f
C53196 _0179_ _0813_/a_109_297# 0.00106f
C53197 _0465_ _1048_/a_975_413# 0
C53198 pp[28] hold80/a_285_47# 0.00874f
C53199 _0996_/a_27_47# _0996_/a_193_47# 0.97021f
C53200 _0965_/a_129_47# control0.count\[1\] 0
C53201 control0.count\[3\] VPWR 1.5227f
C53202 _1048_/a_193_47# net147 0
C53203 net63 acc0.A\[5\] 0.70162f
C53204 _1054_/a_561_413# net9 0
C53205 _0552_/a_68_297# comp0.B\[6\] 0.17771f
C53206 _0990_/a_975_413# _0088_ 0
C53207 _0514_/a_109_297# net66 0.00396f
C53208 _0386_ _0245_ 0.17132f
C53209 net32 net153 0
C53210 _0205_ comp0.B\[9\] 0.02588f
C53211 comp0.B\[5\] _1066_/a_634_159# 0
C53212 _0174_ B[8] 0
C53213 _0982_/a_1059_315# _0264_ 0
C53214 _0100_ _0460_ 0.03596f
C53215 _0999_/a_193_47# _0219_ 0
C53216 _0999_/a_891_413# _0345_ 0.00133f
C53217 _0644_/a_285_47# acc0.A\[14\] 0
C53218 _0793_/a_512_297# _0407_ 0.00221f
C53219 hold63/a_391_47# _1025_/a_27_47# 0
C53220 _0949_/a_59_75# _0477_ 0
C53221 net178 net142 0.00757f
C53222 hold83/a_391_47# _0150_ 0
C53223 acc0.A\[16\] _1017_/a_466_413# 0
C53224 _0234_ _0754_/a_245_297# 0.00196f
C53225 _1060_/a_193_47# _0505_/a_27_297# 0.00538f
C53226 _1060_/a_27_47# _0505_/a_109_297# 0
C53227 _0229_ _0382_ 0
C53228 _0211_ _1035_/a_1059_315# 0
C53229 _0226_ _0237_ 0.11234f
C53230 hold56/a_285_47# hold56/a_391_47# 0.41909f
C53231 hold57/a_285_47# _0957_/a_32_297# 0.00192f
C53232 _0314_ _0359_ 0
C53233 _0175_ _0215_ 0
C53234 _0539_/a_68_297# net20 0
C53235 VPWR _0996_/a_634_159# 0.18921f
C53236 net66 _0512_/a_109_47# 0
C53237 _0995_/a_634_159# net60 0
C53238 _1065_/a_634_159# comp0.B\[0\] 0.00457f
C53239 comp0.B\[7\] _1039_/a_975_413# 0.00101f
C53240 hold53/a_285_47# acc0.A\[25\] 0
C53241 _0965_/a_285_47# clkbuf_1_0__f_clk/a_110_47# 0.00274f
C53242 _0965_/a_47_47# clknet_0_clk 0
C53243 hold68/a_49_47# net199 0
C53244 net215 _0575_/a_109_297# 0.02639f
C53245 clknet_1_1__leaf__0460_ hold77/a_391_47# 0.01911f
C53246 _0682_/a_68_297# _0219_ 0
C53247 _1037_/a_1059_315# net28 0.07587f
C53248 _1034_/a_975_413# comp0.B\[6\] 0
C53249 comp0.B\[2\] _0955_/a_32_297# 0
C53250 net56 clkbuf_1_1__f__0462_/a_110_47# 0.01038f
C53251 _1051_/a_891_413# _1051_/a_975_413# 0.00851f
C53252 _1051_/a_27_47# net137 0.22925f
C53253 _1051_/a_381_47# _1051_/a_561_413# 0.00123f
C53254 _1045_/a_634_159# _1044_/a_466_413# 0
C53255 _1045_/a_466_413# _1044_/a_634_159# 0.0036f
C53256 _1045_/a_1059_315# _1044_/a_193_47# 0.00562f
C53257 _1045_/a_27_47# _1044_/a_891_413# 0
C53258 _1045_/a_891_413# _1044_/a_27_47# 0
C53259 _0743_/a_51_297# _0250_ 0
C53260 _0336_ _0704_/a_68_297# 0.10679f
C53261 _0705_/a_59_75# acc0.A\[30\] 0
C53262 _0227_ _1005_/a_1059_315# 0
C53263 acc0.A\[21\] _1005_/a_891_413# 0
C53264 _1051_/a_634_159# net131 0
C53265 acc0.A\[14\] _0082_ 0.03143f
C53266 pp[27] _0336_ 0.01245f
C53267 net62 _0986_/a_634_159# 0.03587f
C53268 _0369_ net221 0.01892f
C53269 _1070_/a_1017_47# control0.count\[1\] 0
C53270 net106 net119 0
C53271 _1045_/a_1059_315# net131 0
C53272 _1045_/a_466_413# net184 0
C53273 hold56/a_391_47# _1032_/a_193_47# 0
C53274 _0979_/a_27_297# control0.count\[0\] 0
C53275 _0195_ _0186_ 0.02502f
C53276 net23 _1067_/a_1059_315# 0.01461f
C53277 _1003_/a_466_413# net213 0
C53278 _1072_/a_634_159# clknet_1_0__leaf_clk 0.00147f
C53279 VPWR _1043_/a_1017_47# 0
C53280 _0618_/a_510_47# _0219_ 0
C53281 _0218_ _0986_/a_381_47# 0
C53282 _0643_/a_103_199# _0465_ 0.00654f
C53283 clknet_1_0__leaf__0458_ hold100/a_391_47# 0.00228f
C53284 _0361_ _0697_/a_300_47# 0
C53285 _0733_/a_544_297# _0322_ 0
C53286 _0984_/a_193_47# _0158_ 0
C53287 _1018_/a_975_413# _0399_ 0
C53288 _1043_/a_1059_315# net129 0
C53289 _1043_/a_466_413# net196 0.00113f
C53290 _0451_ _0264_ 0.00288f
C53291 hold32/a_391_47# net16 0.00297f
C53292 _1060_/a_193_47# _0506_/a_81_21# 0
C53293 VPWR _0568_/a_109_297# 0.20366f
C53294 VPWR _1015_/a_381_47# 0.07715f
C53295 acc0.A\[21\] _0765_/a_297_297# 0.00356f
C53296 net125 _1048_/a_193_47# 0
C53297 clknet_1_0__leaf__0458_ _0982_/a_466_413# 0
C53298 _0195_ hold19/a_49_47# 0
C53299 clknet_0__0464_ _0540_/a_51_297# 0.0015f
C53300 _1016_/a_193_47# hold72/a_285_47# 0
C53301 net160 B[1] 0.00189f
C53302 _0176_ _1046_/a_891_413# 0
C53303 net103 clkbuf_0__0459_/a_110_47# 0
C53304 _1072_/a_27_47# _0974_/a_79_199# 0
C53305 _0286_ _0282_ 0
C53306 control0.state\[1\] hold84/a_49_47# 0
C53307 control0.state\[0\] hold84/a_285_47# 0.00138f
C53308 _1030_/a_891_413# _0128_ 0
C53309 clknet_1_1__leaf__0460_ _0395_ 0
C53310 clkbuf_0__0464_/a_110_47# _0138_ 0
C53311 _1021_/a_466_413# _0100_ 0
C53312 _0119_ _1002_/a_466_413# 0.00148f
C53313 net53 net52 0.02218f
C53314 _1032_/a_27_47# _1032_/a_466_413# 0.27314f
C53315 _1032_/a_193_47# _1032_/a_634_159# 0.12729f
C53316 net15 _0180_ 0.11575f
C53317 _0343_ _0601_/a_68_297# 0
C53318 _1054_/a_466_413# _1054_/a_592_47# 0.00553f
C53319 _1054_/a_634_159# _1054_/a_1017_47# 0
C53320 hold11/a_285_47# clknet_0__0464_ 0.00186f
C53321 _1071_/a_561_413# control0.count\[0\] 0
C53322 _1015_/a_1059_315# _1015_/a_891_413# 0.31086f
C53323 _1015_/a_193_47# _1015_/a_975_413# 0
C53324 _1015_/a_466_413# _1015_/a_381_47# 0.03733f
C53325 net1 _0399_ 0.00433f
C53326 _0983_/a_592_47# VPWR 0
C53327 clkbuf_1_0__f__0457_/a_110_47# _0586_/a_27_47# 0.01363f
C53328 _0307_ _0308_ 0.05856f
C53329 _0991_/a_466_413# _0347_ 0
C53330 _0357_ _1010_/a_466_413# 0.00132f
C53331 _0108_ _1010_/a_27_47# 0.0989f
C53332 _0557_/a_512_297# _0173_ 0
C53333 _0358_ _1010_/a_634_159# 0.00171f
C53334 _0751_/a_183_297# _0227_ 0
C53335 net113 _1027_/a_891_413# 0
C53336 clknet_1_1__leaf__0462_ _1027_/a_561_413# 0
C53337 _0352_ _0773_/a_285_297# 0.00548f
C53338 _0335_ hold80/a_49_47# 0
C53339 acc0.A\[7\] output63/a_27_47# 0.00852f
C53340 clkbuf_1_0__f__0463_/a_110_47# comp0.B\[8\] 0.00256f
C53341 _0792_/a_209_47# _0408_ 0
C53342 _0343_ _1031_/a_466_413# 0.01029f
C53343 net46 net87 0
C53344 _0399_ clkbuf_1_1__f__0461_/a_110_47# 0.03683f
C53345 VPWR _0550_/a_512_297# 0.00648f
C53346 net10 net153 0.08338f
C53347 pp[16] _0339_ 0
C53348 net247 _1047_/a_634_159# 0
C53349 _1038_/a_193_47# _1038_/a_592_47# 0
C53350 _1038_/a_466_413# _1038_/a_561_413# 0.00772f
C53351 _1038_/a_634_159# _1038_/a_975_413# 0
C53352 _1053_/a_1059_315# _0180_ 0
C53353 _0211_ _1037_/a_193_47# 0.00231f
C53354 _0689_/a_68_297# _0318_ 0
C53355 _0319_ _0686_/a_301_297# 0
C53356 _0203_ _0541_/a_68_297# 0.10751f
C53357 _0283_ _0303_ 0
C53358 _0105_ _0360_ 0.23136f
C53359 _0654_/a_207_413# _0654_/a_297_47# 0.00476f
C53360 _0319_ _1008_/a_381_47# 0
C53361 _1067_/a_27_47# net107 0.00183f
C53362 _1067_/a_634_159# clknet_1_0__leaf__0461_ 0.01286f
C53363 _0924_/a_27_47# _0171_ 0
C53364 _1041_/a_1059_315# _0138_ 0
C53365 clknet_0__0457_ _0782_/a_27_47# 0.01104f
C53366 _0290_ _0812_/a_297_297# 0.00179f
C53367 net231 _0471_ 0
C53368 net40 _0646_/a_377_297# 0.00334f
C53369 VPWR A[12] 0.26253f
C53370 _0647_/a_47_47# _0277_ 0
C53371 clknet_1_0__leaf__0465_ _1044_/a_193_47# 0.00462f
C53372 net145 _0158_ 0.00104f
C53373 hold24/a_49_47# _0473_ 0
C53374 _0983_/a_891_413# _0983_/a_1017_47# 0.00617f
C53375 output47/a_27_47# net141 0.04285f
C53376 _0983_/a_634_159# net69 0
C53377 hold86/a_49_47# clkbuf_0__0458_/a_110_47# 0
C53378 clkbuf_1_0__f__0461_/a_110_47# _0347_ 0
C53379 clknet_1_0__leaf__0465_ net131 0.01024f
C53380 _0352_ _0350_ 0.40788f
C53381 _0262_ _0447_ 0
C53382 _0627_/a_215_53# _0258_ 0.00205f
C53383 net245 _0995_/a_891_413# 0
C53384 net40 _0995_/a_561_413# 0
C53385 _0965_/a_285_47# control0.count\[2\] 0.00113f
C53386 net176 VPWR 0.45443f
C53387 net72 _0841_/a_79_21# 0
C53388 _0283_ _0281_ 0.15225f
C53389 _0659_/a_68_297# acc0.A\[8\] 0.17118f
C53390 _0659_/a_150_297# net66 0
C53391 _0399_ _0185_ 0.00127f
C53392 pp[28] _0220_ 0
C53393 net188 hold45/a_391_47# 0
C53394 _0984_/a_193_47# acc0.A\[14\] 0
C53395 _0294_ clkbuf_0__0460_/a_110_47# 0
C53396 hold69/a_285_47# VPWR 0.32058f
C53397 _0997_/a_193_47# net42 0.47162f
C53398 _0550_/a_51_297# _0550_/a_245_297# 0.01218f
C53399 _0230_ _0600_/a_103_199# 0.09306f
C53400 _0747_/a_79_21# _1006_/a_1059_315# 0.00163f
C53401 _0747_/a_215_47# _1006_/a_634_159# 0
C53402 _0726_/a_51_297# _0725_/a_209_297# 0
C53403 _1056_/a_1059_315# _0154_ 0.00147f
C53404 net1 _0466_ 0
C53405 _0466_ _1068_/a_381_47# 0.01718f
C53406 net90 _1007_/a_561_413# 0
C53407 clknet_1_0__leaf__0459_ net84 0.09983f
C53408 hold21/a_285_47# clknet_1_0__leaf__0465_ 0
C53409 net45 acc0.A\[18\] 0.48531f
C53410 _0835_/a_78_199# acc0.A\[3\] 0
C53411 _1048_/a_1059_315# _1047_/a_193_47# 0
C53412 _1048_/a_634_159# _1047_/a_466_413# 0
C53413 _0253_ _0369_ 0.61646f
C53414 _0278_ _0276_ 0.0353f
C53415 _1054_/a_27_47# acc0.A\[6\] 0.00471f
C53416 clkbuf_1_1__f__0462_/a_110_47# _0345_ 0
C53417 input16/a_75_212# clknet_1_1__leaf__0465_ 0
C53418 hold18/a_49_47# net149 0
C53419 _0317_ _0322_ 0.0944f
C53420 _0244_ net219 0.22863f
C53421 clknet_1_0__leaf__0462_ _1005_/a_634_159# 0
C53422 _1016_/a_381_47# net166 0.12256f
C53423 _1061_/a_634_159# acc0.A\[15\] 0
C53424 hold31/a_49_47# _0254_ 0.00229f
C53425 _0317_ _0327_ 0.1202f
C53426 clknet_1_1__leaf__0462_ _1026_/a_1017_47# 0
C53427 _0629_/a_145_75# acc0.A\[15\] 0
C53428 _0216_ _0336_ 0.00219f
C53429 net84 _0783_/a_79_21# 0
C53430 _0998_/a_1059_315# _0399_ 0
C53431 _0998_/a_466_413# _0096_ 0.04223f
C53432 _0802_/a_59_75# _0414_ 0.15802f
C53433 _0401_ _0347_ 0.00216f
C53434 VPWR _0617_/a_68_297# 0.1781f
C53435 input4/a_75_212# A[12] 0.20577f
C53436 hold17/a_391_47# _0168_ 0
C53437 _0263_ _0841_/a_215_47# 0
C53438 hold11/a_49_47# clknet_1_0__leaf__0464_ 0
C53439 clknet_0__0464_ _0524_/a_27_297# 0
C53440 control0.add control0.reset 0
C53441 _0780_/a_285_297# _0308_ 0.06887f
C53442 _0535_/a_68_297# _0548_/a_149_47# 0
C53443 _0535_/a_68_297# clknet_1_1__leaf__0464_ 0
C53444 hold68/a_49_47# VPWR 0.30013f
C53445 _0559_/a_240_47# VPWR 0.00649f
C53446 _0326_ _0370_ 0.15003f
C53447 _1008_/a_193_47# hold50/a_285_47# 0.01349f
C53448 _1008_/a_27_47# hold50/a_391_47# 0.00132f
C53449 net115 _0350_ 0
C53450 net222 _0347_ 0.0016f
C53451 _0216_ _0585_/a_109_47# 0.00519f
C53452 _1052_/a_466_413# net154 0
C53453 _1052_/a_27_47# net11 0.00203f
C53454 _0961_/a_113_297# _0466_ 0
C53455 _0645_/a_47_47# _0301_ 0
C53456 _1032_/a_592_47# _0352_ 0
C53457 hold62/a_391_47# net209 0.13094f
C53458 _0982_/a_27_47# _1014_/a_193_47# 0
C53459 _0982_/a_193_47# _1014_/a_27_47# 0.00169f
C53460 net145 acc0.A\[14\] 0
C53461 _0459_ net229 0
C53462 _0985_/a_466_413# _0219_ 0
C53463 hold54/a_391_47# comp0.B\[1\] 0.061f
C53464 net183 net20 0.03029f
C53465 _0195_ _1017_/a_193_47# 0.04563f
C53466 net160 _1035_/a_891_413# 0
C53467 _0210_ _1035_/a_1059_315# 0
C53468 clknet_1_1__leaf__0459_ _1057_/a_975_413# 0
C53469 hold64/a_285_47# _1001_/a_193_47# 0
C53470 hold64/a_391_47# _1001_/a_27_47# 0
C53471 _1057_/a_592_47# acc0.A\[11\] 0
C53472 _0179_ _0527_/a_109_47# 0.00208f
C53473 hold4/a_49_47# net151 0
C53474 hold48/a_49_47# net21 0
C53475 _0225_ net50 0.17564f
C53476 _1054_/a_193_47# _0523_/a_299_297# 0
C53477 acc0.A\[0\] _0262_ 0
C53478 hold39/a_49_47# _0213_ 0.03427f
C53479 _0552_/a_68_297# net26 0
C53480 hold17/a_49_47# clkbuf_1_0__f_clk/a_110_47# 0
C53481 _0752_/a_27_413# clknet_1_0__leaf__0460_ 0.01345f
C53482 _1057_/a_193_47# VPWR 0.29352f
C53483 comp0.B\[4\] _1034_/a_891_413# 0.00287f
C53484 _1048_/a_193_47# _0186_ 0
C53485 hold33/a_391_47# net174 0.02828f
C53486 net158 _0143_ 0
C53487 _0663_/a_27_413# net217 0
C53488 VPWR net29 1.3986f
C53489 _1056_/a_561_413# net182 0
C53490 _0647_/a_377_297# _0404_ 0
C53491 _0241_ _0195_ 0
C53492 _0179_ acc0.A\[7\] 0.22322f
C53493 _0241_ net92 0
C53494 net140 VPWR 0.44133f
C53495 _0272_ _0257_ 0.0161f
C53496 _0153_ net16 0.48125f
C53497 clknet_1_1__leaf__0459_ _0096_ 0
C53498 acc0.A\[5\] _0987_/a_1017_47# 0
C53499 _0149_ net73 0.00362f
C53500 net137 _0085_ 0
C53501 _0399_ _0832_/a_113_47# 0
C53502 clknet_1_0__leaf__0459_ _1015_/a_381_47# 0
C53503 _0366_ _1007_/a_27_47# 0.06808f
C53504 _0174_ _0548_/a_149_47# 0.01702f
C53505 _0174_ clknet_1_1__leaf__0464_ 0.02128f
C53506 _0513_/a_299_297# net192 0
C53507 _0992_/a_27_47# _0181_ 0
C53508 _0469_ _0487_ 0
C53509 net154 _0194_ 0.10169f
C53510 net45 hold59/a_49_47# 0
C53511 net186 _0133_ 0
C53512 _0257_ _0837_/a_368_297# 0
C53513 net65 net75 0
C53514 _1050_/a_27_47# clknet_1_1__leaf__0464_ 0
C53515 _0989_/a_466_413# net75 0
C53516 _0312_ clknet_0__0460_ 0.06337f
C53517 _1017_/a_27_47# _0240_ 0
C53518 net35 _1072_/a_891_413# 0.01594f
C53519 _1067_/a_381_47# _0460_ 0
C53520 _1067_/a_975_413# clknet_1_0__leaf__0457_ 0
C53521 _0967_/a_215_297# _0468_ 0.00272f
C53522 _0690_/a_68_297# _0321_ 0.10505f
C53523 _0411_ net42 0
C53524 _1017_/a_27_47# _0369_ 0.02583f
C53525 _0294_ _1009_/a_27_47# 0
C53526 net203 comp0.B\[15\] 0
C53527 _0981_/a_27_297# _1068_/a_27_47# 0
C53528 _0473_ _0954_/a_304_297# 0
C53529 hold101/a_285_47# net62 0
C53530 net185 hold39/a_285_47# 0
C53531 _0607_/a_27_297# _0347_ 0.00968f
C53532 _1059_/a_466_413# net41 0
C53533 hold100/a_285_47# hold18/a_285_47# 0.02819f
C53534 clknet_0__0463_ _0214_ 0.00136f
C53535 _1020_/a_1059_315# net118 0
C53536 _0760_/a_47_47# _0237_ 0.04044f
C53537 _0760_/a_377_297# _0381_ 0.00557f
C53538 _0757_/a_150_297# _0380_ 0
C53539 net178 _0988_/a_27_47# 0.16146f
C53540 _0369_ net74 0.00464f
C53541 _0982_/a_466_413# hold18/a_49_47# 0
C53542 net207 _0350_ 0
C53543 _0286_ _0654_/a_297_47# 0.00132f
C53544 _0343_ hold16/a_285_47# 0.01792f
C53545 _1031_/a_1059_315# _1030_/a_891_413# 0.00126f
C53546 _1031_/a_891_413# _1030_/a_1059_315# 0
C53547 _0983_/a_27_47# _0399_ 0.04907f
C53548 clknet_1_0__leaf__0464_ _0159_ 0
C53549 _0457_ _1067_/a_381_47# 0
C53550 net60 _0345_ 0
C53551 _0181_ hold60/a_49_47# 0
C53552 hold58/a_285_47# _0173_ 0.00517f
C53553 clknet_1_0__leaf__0463_ _1061_/a_193_47# 0.05351f
C53554 clknet_1_1__leaf__0460_ _0329_ 0.0693f
C53555 _0822_/a_109_297# clknet_0__0465_ 0
C53556 net211 net45 0
C53557 _0349_ clknet_1_1__leaf__0462_ 0.02582f
C53558 control0.state\[1\] _0471_ 0.68663f
C53559 net5 _0345_ 0.02001f
C53560 _0498_/a_51_297# _0177_ 0.11636f
C53561 _1038_/a_27_47# _0172_ 0
C53562 _1038_/a_634_159# net180 0
C53563 _1038_/a_193_47# net30 0
C53564 clknet_1_1__leaf__0460_ clknet_1_0__leaf__0460_ 0.00333f
C53565 net160 _1037_/a_634_159# 0
C53566 hold7/a_285_47# net12 0
C53567 _0218_ output40/a_27_47# 0
C53568 _0324_ _1006_/a_891_413# 0
C53569 _1025_/a_466_413# _1025_/a_561_413# 0.00772f
C53570 _1025_/a_634_159# _1025_/a_975_413# 0
C53571 _0289_ _0399_ 0
C53572 acc0.A\[13\] _0669_/a_29_53# 0.06953f
C53573 hold64/a_391_47# _0459_ 0.00533f
C53574 _0389_ _0462_ 0.0024f
C53575 clknet_0__0461_ _0116_ 0
C53576 _0154_ VPWR 0.24584f
C53577 _0369_ output61/a_27_47# 0.00182f
C53578 clkbuf_0__0465_/a_110_47# _0401_ 0
C53579 _0093_ clknet_1_1__leaf__0459_ 0.00602f
C53580 _0114_ _0219_ 0
C53581 net59 _0218_ 0
C53582 hold5/a_391_47# _1042_/a_27_47# 0
C53583 hold5/a_285_47# _1042_/a_193_47# 0
C53584 _0369_ _0973_/a_27_297# 0.06641f
C53585 _0216_ _0208_ 0.22198f
C53586 _0982_/a_193_47# _0195_ 0
C53587 output42/a_27_47# acc0.A\[13\] 0
C53588 acc0.A\[4\] _0196_ 0
C53589 _0168_ _0976_/a_218_47# 0
C53590 control0.count\[1\] _0976_/a_505_21# 0.07195f
C53591 _1070_/a_381_47# _0466_ 0
C53592 hold38/a_285_47# control0.reset 0
C53593 net248 _0625_/a_145_75# 0.00173f
C53594 _0369_ _0772_/a_215_47# 0.05066f
C53595 hold54/a_285_47# _1032_/a_466_413# 0
C53596 hold54/a_391_47# _1032_/a_634_159# 0
C53597 clknet_1_1__leaf__0460_ _0221_ 0.02984f
C53598 clknet_1_1__leaf__0459_ _0808_/a_368_297# 0.00164f
C53599 comp0.B\[5\] _0564_/a_68_297# 0
C53600 net123 input24/a_75_212# 0.01082f
C53601 _0972_/a_250_297# _1063_/a_27_47# 0.02019f
C53602 net38 net79 0
C53603 acc0.A\[11\] _0808_/a_266_47# 0
C53604 _0982_/a_1059_315# _0856_/a_79_21# 0.00135f
C53605 _0982_/a_634_159# _0856_/a_215_47# 0.00117f
C53606 _0403_ _0994_/a_466_413# 0
C53607 hold17/a_49_47# control0.count\[2\] 0.32345f
C53608 clknet_0__0463_ _1061_/a_1059_315# 0
C53609 _0255_ _0438_ 0
C53610 _0473_ _0540_/a_240_47# 0.00131f
C53611 control0.reset clknet_1_1__leaf__0457_ 0
C53612 hold58/a_391_47# _0212_ 0.03469f
C53613 _0996_/a_466_413# _0996_/a_592_47# 0.00553f
C53614 _0996_/a_634_159# _0996_/a_1017_47# 0
C53615 hold59/a_285_47# net104 0.03658f
C53616 _0244_ _0352_ 0.29993f
C53617 hold57/a_49_47# _0173_ 0.03378f
C53618 net45 _1031_/a_891_413# 0
C53619 net204 net8 0
C53620 clknet_0__0463_ _0207_ 0.00142f
C53621 _0174_ net247 0.15691f
C53622 _0753_/a_381_47# acc0.A\[23\] 0
C53623 _0129_ _0708_/a_68_297# 0
C53624 _0849_/a_79_21# _0350_ 0.01207f
C53625 comp0.B\[1\] _0182_ 0
C53626 _0255_ _0636_/a_59_75# 0
C53627 hold53/a_285_47# net210 0.00125f
C53628 net200 _0572_/a_27_297# 0
C53629 _0407_ _0095_ 0.0379f
C53630 clknet_1_1__leaf__0457_ _1061_/a_891_413# 0
C53631 pp[19] pp[22] 0.17884f
C53632 _0730_/a_79_21# _0685_/a_68_297# 0
C53633 _0375_ net241 0.00623f
C53634 _1060_/a_193_47# _0184_ 0
C53635 _1060_/a_466_413# net6 0
C53636 _1052_/a_27_47# clknet_1_1__leaf__0458_ 0
C53637 _0607_/a_27_297# _1016_/a_891_413# 0
C53638 _0714_/a_245_297# _0341_ 0.0024f
C53639 _0714_/a_51_297# _0340_ 0
C53640 _0559_/a_245_297# _0559_/a_240_47# 0
C53641 _0698_/a_113_297# _0318_ 0
C53642 hold42/a_285_47# clknet_1_1__leaf__0465_ 0.03099f
C53643 hold70/a_285_47# net228 0.08056f
C53644 clknet_1_0__leaf__0463_ _1039_/a_193_47# 0.00333f
C53645 _0701_/a_209_297# clknet_1_1__leaf__0462_ 0
C53646 VPWR _1036_/a_466_413# 0.25507f
C53647 _1057_/a_1059_315# clknet_1_1__leaf__0465_ 0.02461f
C53648 clknet_0__0458_ _0265_ 0
C53649 hold24/a_391_47# _0174_ 0.00601f
C53650 net98 _0776_/a_27_47# 0
C53651 clknet_0__0457_ _0982_/a_27_47# 0.00221f
C53652 _1044_/a_27_47# _1044_/a_1059_315# 0.04875f
C53653 _1044_/a_193_47# _1044_/a_466_413# 0.07402f
C53654 _0354_ acc0.A\[29\] 0.04181f
C53655 _0274_ _0640_/a_297_297# 0
C53656 _0643_/a_103_199# _0254_ 0
C53657 _0275_ _0640_/a_109_53# 0
C53658 hold11/a_285_47# _0536_/a_51_297# 0
C53659 VPWR _0725_/a_209_297# 0.19638f
C53660 comp0.B\[2\] _0474_ 0.02349f
C53661 _0149_ _1044_/a_27_47# 0
C53662 hold52/a_285_47# _0575_/a_27_297# 0
C53663 _0966_/a_109_297# VPWR 0.00385f
C53664 _1056_/a_27_47# net16 0.00347f
C53665 hold65/a_285_47# _0087_ 0
C53666 net131 _1044_/a_466_413# 0
C53667 clknet_1_1__leaf__0459_ _0395_ 0
C53668 _0383_ net51 0.09194f
C53669 _1021_/a_193_47# _0764_/a_81_21# 0
C53670 _0349_ net242 0.03149f
C53671 _0992_/a_1017_47# acc0.A\[10\] 0.00125f
C53672 net137 net131 0
C53673 _0442_ _0346_ 0.09742f
C53674 _0548_/a_51_297# _0206_ 0.11448f
C53675 _0430_ _0824_/a_59_75# 0.00112f
C53676 clkload3/a_268_47# _0306_ 0
C53677 _0803_/a_68_297# VPWR 0.20453f
C53678 net98 _0219_ 0
C53679 hold56/a_49_47# net202 0
C53680 _0802_/a_59_75# _0404_ 0.13068f
C53681 _0169_ control0.count\[0\] 0
C53682 acc0.A\[11\] _0345_ 0
C53683 _0101_ net213 0.30985f
C53684 net46 _1023_/a_634_159# 0.00549f
C53685 output46/a_27_47# _1023_/a_891_413# 0.01437f
C53686 control0.state\[1\] hold93/a_391_47# 0
C53687 clknet_1_0__leaf__0458_ net206 0
C53688 hold56/a_49_47# clknet_1_1__leaf__0463_ 0.01118f
C53689 _0399_ _0793_/a_149_47# 0
C53690 _0789_/a_208_47# VPWR 0.00212f
C53691 _0369_ net17 0
C53692 clknet_0__0459_ _0399_ 0.0268f
C53693 clknet_1_1__leaf__0459_ _0304_ 0
C53694 _0369_ net238 0.09786f
C53695 _0359_ _0360_ 0.11003f
C53696 _0346_ _0374_ 0
C53697 _0714_/a_240_47# _1013_/a_634_159# 0
C53698 _0443_ clkbuf_0__0465_/a_110_47# 0.04442f
C53699 clknet_1_0__leaf__0458_ _0080_ 0
C53700 _0575_/a_27_297# net52 0.01022f
C53701 VPWR _0673_/a_337_297# 0.00291f
C53702 _0458_ net10 0.00307f
C53703 clkload3/Y _0219_ 0.01279f
C53704 _0343_ _0819_/a_299_297# 0
C53705 hold101/a_49_47# _0270_ 0
C53706 net58 _0275_ 0.02406f
C53707 VPWR _0672_/a_215_47# 0.00454f
C53708 _0627_/a_297_297# clknet_1_1__leaf__0458_ 0
C53709 _0627_/a_215_53# net72 0
C53710 _0972_/a_250_297# _1062_/a_1059_315# 0
C53711 _0259_ _0817_/a_81_21# 0.01022f
C53712 _0858_/a_27_47# _0532_/a_384_47# 0
C53713 clknet_1_0__leaf__0463_ _1040_/a_592_47# 0
C53714 _0119_ _0100_ 0
C53715 A[9] pp[4] 0
C53716 _1032_/a_27_47# net202 0.12587f
C53717 _1032_/a_1059_315# _1032_/a_1017_47# 0
C53718 _1054_/a_592_47# net169 0
C53719 _1015_/a_381_47# _0113_ 0.13122f
C53720 output42/a_27_47# net245 0.00561f
C53721 pp[15] hold98/a_391_47# 0.02195f
C53722 _0288_ _0508_/a_299_297# 0
C53723 _1057_/a_193_47# _0283_ 0
C53724 net113 _0319_ 0
C53725 _1032_/a_27_47# clknet_1_1__leaf__0463_ 0
C53726 _0089_ _0347_ 0.02054f
C53727 _0374_ hold94/a_49_47# 0.04492f
C53728 VPWR input14/a_75_212# 0.24709f
C53729 _0134_ _0173_ 0.00119f
C53730 _0578_/a_27_297# _0721_/a_27_47# 0
C53731 _0343_ _0437_ 0.07189f
C53732 _0226_ _0222_ 0
C53733 _0233_ clknet_1_0__leaf__0460_ 0.06396f
C53734 VPWR acc0.A\[18\] 0.73921f
C53735 _1051_/a_381_47# _0180_ 0.00634f
C53736 hold46/a_49_47# _0540_/a_51_297# 0
C53737 _0820_/a_79_21# _0990_/a_1059_315# 0.01742f
C53738 VPWR _0137_ 1.61868f
C53739 _1014_/a_592_47# net149 0.00285f
C53740 _1014_/a_1059_315# _0112_ 0
C53741 _0310_ _0614_/a_29_53# 0
C53742 _0783_/a_79_21# _0783_/a_510_47# 0.00844f
C53743 _0783_/a_297_297# _0783_/a_215_47# 0
C53744 _0716_/a_27_47# _0346_ 0.24882f
C53745 _0385_ _0373_ 0.00632f
C53746 _0346_ net165 0.21417f
C53747 net242 _0701_/a_209_297# 0
C53748 comp0.B\[13\] clknet_1_1__leaf__0464_ 0.11096f
C53749 comp0.B\[7\] _0173_ 0
C53750 hold44/a_49_47# VPWR 0.31572f
C53751 _0765_/a_79_21# _0352_ 0.1511f
C53752 acc0.A\[27\] _1028_/a_27_47# 0.03749f
C53753 _0315_ _0460_ 0
C53754 _0343_ _1055_/a_193_47# 0.002f
C53755 hold25/a_285_47# comp0.B\[8\] 0
C53756 _0343_ _0791_/a_199_47# 0
C53757 control0.state\[1\] control0.reset 0
C53758 _0259_ _0084_ 0
C53759 net81 _0218_ 0.18246f
C53760 hold81/a_391_47# _0345_ 0.00563f
C53761 hold27/a_49_47# net10 0
C53762 net163 _1030_/a_27_47# 0
C53763 _1020_/a_891_413# net1 0.00245f
C53764 clkbuf_1_1__f__0465_/a_110_47# _0088_ 0.00206f
C53765 _0289_ _0295_ 0.38254f
C53766 net168 _1052_/a_634_159# 0
C53767 net108 _0222_ 0
C53768 _0997_/a_381_47# net43 0.02548f
C53769 acc0.A\[21\] _0369_ 0.26911f
C53770 net9 _0150_ 0.09085f
C53771 _0352_ _1006_/a_634_159# 0.01551f
C53772 pp[1] _0988_/a_193_47# 0
C53773 _0454_ _0451_ 0
C53774 _0287_ _0296_ 0
C53775 VPWR _0995_/a_891_413# 0.19937f
C53776 _0284_ _0993_/a_634_159# 0.0011f
C53777 clknet_0__0457_ acc0.A\[21\] 0
C53778 clknet_1_0__leaf__0458_ _0637_/a_139_47# 0
C53779 _0346_ acc0.A\[19\] 0
C53780 hold87/a_285_47# _0350_ 0
C53781 VPWR _0605_/a_109_297# 0.00447f
C53782 output42/a_27_47# net45 0
C53783 _0280_ _0670_/a_510_47# 0
C53784 hold28/a_391_47# _1048_/a_891_413# 0.00406f
C53785 net150 _0460_ 0.0361f
C53786 _0216_ _0747_/a_79_21# 0.00998f
C53787 _0550_/a_149_47# net180 0.00683f
C53788 hold23/a_391_47# net170 0.18044f
C53789 _0550_/a_512_297# net30 0.00101f
C53790 net216 _1006_/a_975_413# 0
C53791 _0662_/a_299_297# _0275_ 0.05387f
C53792 _1013_/a_1059_315# net41 0
C53793 _0247_ _0393_ 0.11832f
C53794 _0104_ _1006_/a_891_413# 0
C53795 _0126_ _1008_/a_634_159# 0
C53796 net190 _1008_/a_891_413# 0
C53797 _0443_ _0824_/a_59_75# 0
C53798 _0355_ _0725_/a_303_47# 0
C53799 _0968_/a_109_297# clknet_1_0__leaf_clk 0
C53800 _0226_ net220 0
C53801 acc0.A\[12\] _1058_/a_1017_47# 0.00174f
C53802 _0282_ net79 0
C53803 _0180_ _0268_ 0
C53804 clkbuf_0__0464_/a_110_47# net22 0
C53805 acc0.A\[24\] _1007_/a_27_47# 0.01478f
C53806 hold71/a_49_47# hold71/a_391_47# 0.00188f
C53807 hold14/a_285_47# _0211_ 0.06808f
C53808 pp[9] output47/a_27_47# 0
C53809 _1000_/a_381_47# _0461_ 0.002f
C53810 output66/a_27_47# hold34/a_285_47# 0.00143f
C53811 VPWR comp0.B\[6\] 1.81598f
C53812 _0272_ clknet_1_1__leaf__0458_ 0.17314f
C53813 comp0.B\[12\] comp0.B\[10\] 0
C53814 net147 acc0.A\[15\] 0
C53815 hold45/a_49_47# acc0.A\[11\] 0.33674f
C53816 _0216_ hold9/a_49_47# 0
C53817 _0195_ hold9/a_391_47# 0.02869f
C53818 clkbuf_1_1__f__0463_/a_110_47# net23 0
C53819 VPWR _1023_/a_466_413# 0.25139f
C53820 net157 _0545_/a_68_297# 0
C53821 _1047_/a_193_47# clkbuf_1_1__f__0457_/a_110_47# 0.02077f
C53822 _1036_/a_975_413# _0175_ 0
C53823 _0240_ _0245_ 0.41391f
C53824 _0534_/a_299_297# _0199_ 0.00863f
C53825 _0446_ _0844_/a_79_21# 0.12245f
C53826 hold59/a_49_47# VPWR 0.31166f
C53827 _0369_ _0245_ 0
C53828 _0313_ _0365_ 0
C53829 comp0.B\[14\] _0540_/a_51_297# 0.02404f
C53830 comp0.B\[15\] _0176_ 0
C53831 _0991_/a_193_47# _0991_/a_381_47# 0.09799f
C53832 _0991_/a_634_159# _0991_/a_891_413# 0.03684f
C53833 _0991_/a_27_47# _0991_/a_561_413# 0.0027f
C53834 _0726_/a_149_47# _0345_ 0.00154f
C53835 _0236_ _0763_/a_109_47# 0
C53836 clknet_0__0464_ _0194_ 0
C53837 net21 _0203_ 0.02888f
C53838 _0346_ _0249_ 0.0323f
C53839 clknet_0__0458_ _0267_ 0.04693f
C53840 _0794_/a_27_47# _0794_/a_326_47# 0.0034f
C53841 _0432_ _0268_ 0
C53842 clknet_1_0__leaf__0463_ clkbuf_0__0464_/a_110_47# 0
C53843 _1041_/a_1059_315# net22 0
C53844 _0747_/a_297_297# _0369_ 0.00328f
C53845 _0461_ _0565_/a_51_297# 0
C53846 _0773_/a_285_297# _0392_ 0.07632f
C53847 _0216_ _1029_/a_27_47# 0.04627f
C53848 hold26/a_49_47# net157 0
C53849 net160 _0473_ 0
C53850 net233 hold18/a_285_47# 0
C53851 net94 hold50/a_49_47# 0.0012f
C53852 _0183_ _0635_/a_109_297# 0
C53853 net48 _0605_/a_109_297# 0
C53854 _0799_/a_80_21# acc0.A\[13\] 0.00114f
C53855 net100 _0208_ 0.01165f
C53856 _0793_/a_245_297# _0345_ 0.00285f
C53857 _0083_ _0219_ 0.01564f
C53858 clknet_1_1__leaf__0459_ _0811_/a_384_47# 0
C53859 net55 _0360_ 0
C53860 net7 _1046_/a_27_47# 0
C53861 _1001_/a_466_413# _0183_ 0.00375f
C53862 _1001_/a_891_413# _0217_ 0
C53863 clknet_1_0__leaf__0463_ _1037_/a_193_47# 0.001f
C53864 net186 _0208_ 0
C53865 control0.state\[0\] _0948_/a_109_297# 0
C53866 _0399_ _0996_/a_1059_315# 0.02376f
C53867 _0520_/a_27_297# net138 0
C53868 net45 _0611_/a_150_297# 0
C53869 acc0.A\[17\] _0394_ 0
C53870 net176 pp[22] 0
C53871 _0598_/a_297_47# _0369_ 0
C53872 _0230_ _0762_/a_79_21# 0.00508f
C53873 _0598_/a_79_21# _0383_ 0.01963f
C53874 net211 VPWR 0.25107f
C53875 _0808_/a_266_47# _0281_ 0.04973f
C53876 _0808_/a_266_297# _0418_ 0
C53877 _0543_/a_68_297# _0540_/a_51_297# 0.00163f
C53878 _1021_/a_634_159# _0217_ 0.01716f
C53879 _1021_/a_27_47# _0183_ 0.00656f
C53880 hold35/a_391_47# _0154_ 0
C53881 _0548_/a_149_47# comp0.B\[9\] 0.02894f
C53882 _0854_/a_215_47# _0347_ 0.05706f
C53883 clkbuf_1_1__f__0461_/a_110_47# _0306_ 0.00578f
C53884 _0731_/a_384_47# _0326_ 0.00121f
C53885 clknet_0__0458_ _0642_/a_215_297# 0
C53886 _0665_/a_109_297# _0299_ 0.00178f
C53887 _1058_/a_1059_315# acc0.A\[10\] 0.06211f
C53888 _0218_ _0797_/a_207_413# 0.00248f
C53889 _0391_ _0771_/a_215_297# 0.11562f
C53890 clknet_1_0__leaf__0465_ _0525_/a_81_21# 0.0148f
C53891 _0446_ _0846_/a_240_47# 0.00267f
C53892 net125 acc0.A\[15\] 0.08226f
C53893 _0195_ net136 0
C53894 _0600_/a_103_199# _0380_ 0
C53895 _0234_ _1003_/a_1059_315# 0
C53896 _0218_ _0841_/a_215_47# 0.00104f
C53897 _0546_/a_51_297# _1042_/a_27_47# 0
C53898 net158 _0174_ 0
C53899 _0305_ clkload4/Y 0.00889f
C53900 _0361_ _0318_ 0.28443f
C53901 _0619_/a_68_297# _0436_ 0
C53902 _0719_/a_27_47# control0.add 0.2039f
C53903 _0522_/a_27_297# _0193_ 0.16788f
C53904 _0303_ _0345_ 0.00766f
C53905 _0722_/a_510_47# _0352_ 0.00381f
C53906 _0800_/a_51_297# _0413_ 0.11253f
C53907 _0800_/a_245_297# _0412_ 0.00176f
C53908 control0.add _0460_ 0.00167f
C53909 _0461_ _1018_/a_466_413# 0
C53910 _0371_ clkbuf_0__0460_/a_110_47# 0
C53911 net201 _0563_/a_51_297# 0
C53912 _0170_ _1068_/a_27_47# 0
C53913 net167 _1068_/a_466_413# 0
C53914 _0996_/a_891_413# _0277_ 0
C53915 net168 A[8] 0.21217f
C53916 _0483_ _0466_ 0.09185f
C53917 VPWR _1031_/a_891_413# 0.19427f
C53918 clknet_1_0__leaf__0459_ acc0.A\[18\] 0.05595f
C53919 clkbuf_0__0465_/a_110_47# _0986_/a_891_413# 0.01365f
C53920 clknet_0__0465_ _0986_/a_27_47# 0.00955f
C53921 _0295_ _0655_/a_109_93# 0
C53922 _0216_ _1019_/a_193_47# 0
C53923 net88 _0487_ 0.00189f
C53924 acc0.A\[12\] _0648_/a_27_297# 0.00628f
C53925 net203 _0176_ 0
C53926 _0287_ _0811_/a_81_21# 0
C53927 _0290_ _0991_/a_891_413# 0
C53928 _0891_/a_27_47# net1 0
C53929 output44/a_27_47# _0221_ 0
C53930 net56 _0568_/a_109_297# 0
C53931 _1043_/a_27_47# hold51/a_391_47# 0.0042f
C53932 _1043_/a_193_47# hold51/a_285_47# 0.0148f
C53933 hold68/a_391_47# net50 0.06882f
C53934 _0457_ control0.add 0
C53935 _0372_ clknet_1_0__leaf__0457_ 0
C53936 net51 _1022_/a_1017_47# 0
C53937 net61 _0369_ 0.04172f
C53938 _0345_ _0281_ 0.02408f
C53939 net205 _0132_ 0
C53940 _0820_/a_79_21# VPWR 0.45499f
C53941 _0596_/a_59_75# net49 0.19594f
C53942 _0971_/a_81_21# _1063_/a_27_47# 0
C53943 hold41/a_285_47# output67/a_27_47# 0.00293f
C53944 clkbuf_1_0__f__0458_/a_110_47# _0450_ 0.01561f
C53945 _0486_ clknet_1_0__leaf_clk 0.05969f
C53946 _0399_ pp[4] 0
C53947 hold15/a_391_47# _0336_ 0
C53948 _0154_ net182 0
C53949 hold44/a_391_47# _0569_/a_27_297# 0.01653f
C53950 hold44/a_285_47# _0569_/a_109_297# 0
C53951 _1004_/a_891_413# clknet_1_0__leaf__0460_ 0.00242f
C53952 _0523_/a_299_297# acc0.A\[6\] 0
C53953 _0251_ hold65/a_49_47# 0.03522f
C53954 _0195_ net219 0.02161f
C53955 _1025_/a_1059_315# acc0.A\[25\] 0.12819f
C53956 _1020_/a_193_47# _1015_/a_193_47# 0
C53957 _1020_/a_634_159# _1015_/a_27_47# 0
C53958 _1020_/a_27_47# _1015_/a_634_159# 0
C53959 _1030_/a_975_413# _0221_ 0
C53960 _0971_/a_299_297# clknet_1_0__leaf__0457_ 0
C53961 hold5/a_49_47# net128 0.01387f
C53962 _0369_ _0165_ 0
C53963 clknet_1_0__leaf__0457_ hold40/a_49_47# 0.00152f
C53964 net54 _1008_/a_634_159# 0.00411f
C53965 _0217_ _0586_/a_27_47# 0.00562f
C53966 acc0.A\[12\] output39/a_27_47# 0
C53967 control0.count\[1\] _0466_ 0.23617f
C53968 _0962_/a_109_297# _0479_ 0
C53969 hold20/a_391_47# _1072_/a_634_159# 0
C53970 hold20/a_49_47# _1072_/a_1059_315# 0.0037f
C53971 clknet_0__0457_ _1019_/a_634_159# 0.00301f
C53972 clkbuf_1_0__f__0457_/a_110_47# _1019_/a_891_413# 0
C53973 net236 _0483_ 0.10128f
C53974 _0244_ hold72/a_285_47# 0
C53975 _0164_ _1063_/a_27_47# 0
C53976 _1021_/a_466_413# control0.add 0
C53977 hold63/a_285_47# _0572_/a_109_297# 0.00197f
C53978 hold63/a_391_47# _0572_/a_27_297# 0
C53979 acc0.A\[14\] _0302_ 0.03985f
C53980 _1036_/a_27_47# _1036_/a_466_413# 0.27314f
C53981 _1036_/a_193_47# _1036_/a_634_159# 0.12729f
C53982 _0090_ hold70/a_285_47# 0
C53983 net84 _0345_ 0
C53984 _1047_/a_1059_315# acc0.A\[15\] 0
C53985 _0769_/a_299_297# _0244_ 0.01645f
C53986 _0769_/a_81_21# _0386_ 0.05911f
C53987 net36 _0175_ 0
C53988 net206 _0247_ 0.00141f
C53989 _0183_ hold19/a_49_47# 0
C53990 _0217_ hold19/a_391_47# 0
C53991 net231 _0460_ 0
C53992 _0993_/a_466_413# _0218_ 0
C53993 _0644_/a_47_47# _0644_/a_377_297# 0.00899f
C53994 clknet_1_0__leaf__0458_ clknet_0__0465_ 0
C53995 _0994_/a_466_413# acc0.A\[13\] 0
C53996 net200 _0124_ 0.00525f
C53997 _1049_/a_193_47# net154 0
C53998 _0108_ _0685_/a_150_297# 0
C53999 hold68/a_285_47# net215 0.01024f
C54000 _0523_/a_299_297# _0523_/a_384_47# 0
C54001 net214 _0292_ 0
C54002 _0158_ net6 0.03069f
C54003 hold27/a_285_47# _0498_/a_51_297# 0
C54004 net226 _0978_/a_109_297# 0.01144f
C54005 acc0.A\[16\] _1016_/a_1017_47# 0.0016f
C54006 hold59/a_49_47# clknet_1_0__leaf__0459_ 0
C54007 net225 _0340_ 0
C54008 hold31/a_49_47# _0273_ 0
C54009 _0176_ _0546_/a_149_47# 0
C54010 _0422_ net67 0.45115f
C54011 _1041_/a_891_413# _0544_/a_51_297# 0
C54012 _1041_/a_193_47# _0544_/a_240_47# 0
C54013 clkload1/Y _0433_ 0
C54014 VPWR net161 0.39119f
C54015 hold54/a_391_47# _0180_ 0
C54016 _1050_/a_27_47# net148 0
C54017 _1059_/a_1059_315# clkbuf_0__0459_/a_110_47# 0.0152f
C54018 comp0.B\[2\] _0563_/a_51_297# 0
C54019 _0403_ _0787_/a_209_297# 0.00283f
C54020 clknet_1_0__leaf__0463_ _0953_/a_114_297# 0.0016f
C54021 _1044_/a_891_413# _1044_/a_1017_47# 0.00617f
C54022 _1044_/a_634_159# net130 0
C54023 _1065_/a_193_47# _0175_ 0.00254f
C54024 _0292_ _0813_/a_109_297# 0.00114f
C54025 _0181_ clknet_1_1__leaf__0458_ 0
C54026 hold33/a_391_47# hold46/a_49_47# 0.00142f
C54027 _0606_/a_297_297# _0383_ 0
C54028 _0343_ _0252_ 0
C54029 hold49/a_391_47# _0542_/a_51_297# 0.01217f
C54030 VPWR _0776_/a_109_297# 0.00404f
C54031 _0401_ _0425_ 0.01974f
C54032 _0985_/a_1059_315# _0465_ 0.00236f
C54033 _0971_/a_81_21# _1062_/a_1059_315# 0.01733f
C54034 net184 net130 0
C54035 _0682_/a_150_297# _1007_/a_27_47# 0
C54036 _0682_/a_68_297# _1007_/a_193_47# 0
C54037 _1058_/a_1059_315# _0510_/a_109_297# 0
C54038 _0995_/a_27_47# _0297_ 0
C54039 _0804_/a_79_21# acc0.A\[12\] 0
C54040 net36 _1038_/a_1059_315# 0
C54041 pp[0] _1038_/a_634_159# 0
C54042 clknet_1_1__leaf_clk _1065_/a_381_47# 0.01419f
C54043 _0777_/a_47_47# _0777_/a_377_297# 0.00899f
C54044 net238 _0409_ 0
C54045 _1049_/a_193_47# _0465_ 0
C54046 net55 net59 0
C54047 _0368_ _1007_/a_634_159# 0
C54048 _0218_ _0790_/a_35_297# 0
C54049 _0624_/a_59_75# _0835_/a_215_47# 0
C54050 _0985_/a_1059_315# acc0.A\[2\] 0
C54051 _0467_ _0974_/a_79_199# 0.00414f
C54052 _0427_ _0990_/a_27_47# 0
C54053 hold86/a_49_47# _0447_ 0.00397f
C54054 net61 _0844_/a_79_21# 0.07636f
C54055 _0237_ _1005_/a_1059_315# 0
C54056 _0585_/a_109_297# clkbuf_1_1__f__0457_/a_110_47# 0.0023f
C54057 VPWR net26 1.60571f
C54058 _0675_/a_68_297# _0459_ 0.00208f
C54059 _0670_/a_79_21# net41 0.09143f
C54060 net46 net109 0
C54061 _0195_ _1028_/a_561_413# 0.00203f
C54062 _0216_ _1028_/a_891_413# 0
C54063 net57 _0723_/a_207_413# 0.00768f
C54064 _1057_/a_466_413# _1057_/a_561_413# 0.00772f
C54065 _1057_/a_634_159# _1057_/a_975_413# 0
C54066 _0258_ _0838_/a_109_297# 0.00232f
C54067 VPWR net241 0.15219f
C54068 _0426_ _0346_ 0.0688f
C54069 acc0.A\[2\] _1049_/a_193_47# 0
C54070 B[13] _1042_/a_466_413# 0
C54071 _0269_ _0986_/a_466_413# 0
C54072 _0984_/a_193_47# _0991_/a_193_47# 0
C54073 net211 clknet_1_0__leaf__0459_ 0.0293f
C54074 pp[17] hold78/a_49_47# 0.00176f
C54075 _0111_ _1013_/a_1059_315# 0.00226f
C54076 _0455_ net206 0
C54077 VPWR _1064_/a_381_47# 0.07375f
C54078 _0789_/a_75_199# _0789_/a_208_47# 0.0159f
C54079 _0789_/a_201_297# _0789_/a_544_297# 0.00702f
C54080 _0412_ _0995_/a_27_47# 0
C54081 _1059_/a_634_159# _1059_/a_975_413# 0
C54082 _1059_/a_466_413# _1059_/a_561_413# 0.00772f
C54083 VPWR _0669_/a_29_53# 0.15013f
C54084 A[11] acc0.A\[9\] 0
C54085 hold59/a_391_47# _0266_ 0
C54086 net231 _1062_/a_891_413# 0.02063f
C54087 hold13/a_285_47# net160 0.00997f
C54088 hold13/a_49_47# _0210_ 0
C54089 hold19/a_49_47# acc0.A\[15\] 0
C54090 _0458_ _0146_ 0.00229f
C54091 _0528_/a_299_297# _0528_/a_384_47# 0
C54092 _1015_/a_381_47# _0345_ 0
C54093 _0568_/a_109_297# _0345_ 0.00663f
C54094 _0153_ net142 0.031f
C54095 clkload4/Y _0181_ 0.02822f
C54096 output42/a_27_47# VPWR 0.2784f
C54097 net33 _0175_ 0
C54098 hold101/a_391_47# _0431_ 0
C54099 _0181_ _1047_/a_27_47# 0.00637f
C54100 _0682_/a_68_297# _0328_ 0
C54101 _0982_/a_1017_47# net247 0
C54102 _0820_/a_510_47# clknet_1_1__leaf__0465_ 0.00167f
C54103 _0673_/a_103_199# _0673_/a_253_297# 0.01483f
C54104 clknet_1_0__leaf__0458_ _0849_/a_215_47# 0.004f
C54105 _0924_/a_27_47# _0464_ 0.10939f
C54106 _0520_/a_27_297# hold83/a_285_47# 0.0015f
C54107 _0181_ _0582_/a_373_47# 0
C54108 _0679_/a_68_297# _0347_ 0
C54109 acc0.A\[5\] _0180_ 0
C54110 net193 _0540_/a_240_47# 0.04825f
C54111 acc0.A\[14\] net6 1.57338f
C54112 _0672_/a_79_21# _0672_/a_297_297# 0.01735f
C54113 _0244_ _0392_ 0.03521f
C54114 _1058_/a_891_413# _0181_ 0.00101f
C54115 net23 _0163_ 0.00568f
C54116 _0369_ _0812_/a_215_47# 0.0548f
C54117 _1030_/a_193_47# clknet_1_1__leaf__0462_ 0
C54118 pp[17] _0129_ 0
C54119 net44 net163 0
C54120 _0984_/a_634_159# _0350_ 0
C54121 _0337_ _0336_ 0.2201f
C54122 _0179_ clkbuf_1_1__f__0464_/a_110_47# 0
C54123 net158 comp0.B\[13\] 0.00185f
C54124 net61 _0846_/a_240_47# 0.00136f
C54125 _0372_ _0748_/a_299_297# 0.00103f
C54126 _0430_ _0432_ 0
C54127 net40 _0994_/a_891_413# 0
C54128 VPWR _1008_/a_193_47# 0.31117f
C54129 _0960_/a_109_47# control0.count\[0\] 0
C54130 net120 _0133_ 0
C54131 _0180_ _0528_/a_299_297# 0
C54132 hold100/a_391_47# _0448_ 0
C54133 net158 _1046_/a_193_47# 0.24269f
C54134 _0467_ _1062_/a_193_47# 0
C54135 _0216_ _0739_/a_79_21# 0.00132f
C54136 _0949_/a_59_75# _0469_ 0.13282f
C54137 _0195_ _0352_ 0
C54138 _0432_ acc0.A\[5\] 0.00159f
C54139 _1003_/a_27_47# _0166_ 0
C54140 _0352_ net92 0
C54141 _0785_/a_81_21# _0819_/a_81_21# 0.00117f
C54142 hold39/a_285_47# net119 0
C54143 clknet_1_0__leaf__0458_ hold71/a_285_47# 0.01f
C54144 _0386_ clknet_0__0461_ 0
C54145 rst B[0] 0.00942f
C54146 _0179_ _0186_ 1.46958f
C54147 _0949_/a_145_75# _0468_ 0
C54148 VPWR _0826_/a_27_53# 0.08302f
C54149 clkbuf_1_1__f__0463_/a_110_47# _0213_ 0.0171f
C54150 _0972_/a_584_47# net17 0.00294f
C54151 _0217_ net149 0.71814f
C54152 _1036_/a_193_47# comp0.B\[5\] 0
C54153 _0399_ _0297_ 0.02495f
C54154 pp[18] _0219_ 0
C54155 _1056_/a_1059_315# net181 0.0082f
C54156 _0183_ _1017_/a_193_47# 0
C54157 VPWR _0611_/a_150_297# 0.00115f
C54158 _1030_/a_27_47# _0720_/a_68_297# 0
C54159 net30 _0137_ 0.25111f
C54160 acc0.A\[1\] net8 0
C54161 _0182_ _0180_ 0.6454f
C54162 _1000_/a_634_159# _0459_ 0
C54163 _0968_/a_193_297# clk 0
C54164 control0.state\[0\] clkbuf_0_clk/a_110_47# 0.018f
C54165 comp0.B\[0\] _1062_/a_193_47# 0
C54166 pp[27] hold95/a_285_47# 0.00187f
C54167 _0152_ acc0.A\[8\] 0
C54168 _0182_ net218 0.02196f
C54169 clknet_0__0463_ _0472_ 0.17994f
C54170 _0181_ clknet_1_0__leaf__0461_ 0.17119f
C54171 hold76/a_49_47# net104 0
C54172 B[12] net19 0
C54173 net105 _1014_/a_193_47# 0
C54174 net207 _1014_/a_27_47# 0.002f
C54175 control0.state\[1\] _1063_/a_193_47# 0.04989f
C54176 net45 _0461_ 0.08747f
C54177 _0183_ _0241_ 0.02998f
C54178 VPWR hold84/a_285_47# 0.30178f
C54179 _0156_ acc0.A\[11\] 0.35786f
C54180 clknet_1_0__leaf__0462_ _1022_/a_891_413# 0.0069f
C54181 _0123_ _1024_/a_891_413# 0
C54182 _1005_/a_193_47# _1005_/a_466_413# 0.07855f
C54183 _1005_/a_27_47# _1005_/a_1059_315# 0.04875f
C54184 _0978_/a_373_47# _0485_ 0
C54185 _0383_ hold3/a_391_47# 0
C54186 net55 _0335_ 0
C54187 _0334_ net209 0
C54188 VPWR _0511_/a_81_21# 0.21069f
C54189 _0546_/a_240_47# _0139_ 0
C54190 VPWR net177 0.3736f
C54191 _0984_/a_1059_315# _0849_/a_215_47# 0
C54192 acc0.A\[20\] net118 0
C54193 _0222_ _0350_ 0
C54194 _1013_/a_27_47# _1013_/a_193_47# 0.97064f
C54195 acc0.A\[16\] _0387_ 0
C54196 control0.state\[1\] _0460_ 0.09189f
C54197 _0991_/a_193_47# net67 0
C54198 _0991_/a_1059_315# _0089_ 0
C54199 _0991_/a_891_413# net77 0
C54200 _1067_/a_891_413# _0487_ 0
C54201 net227 _0219_ 0.131f
C54202 net226 _0480_ 0.01276f
C54203 net205 net25 0
C54204 _1043_/a_891_413# _0541_/a_68_297# 0
C54205 net53 hold90/a_391_47# 0.00695f
C54206 _0497_/a_68_297# acc0.A\[15\] 0.17101f
C54207 hold96/a_49_47# _0352_ 0
C54208 _0366_ _0740_/a_113_47# 0.00938f
C54209 _0985_/a_634_159# _0261_ 0.00555f
C54210 _0607_/a_27_297# _0607_/a_109_297# 0.17136f
C54211 clknet_1_1__leaf__0459_ _0997_/a_27_47# 0.03162f
C54212 _0195_ net115 0
C54213 _0414_ _0404_ 0.16957f
C54214 clknet_0__0458_ net63 0
C54215 clknet_1_1__leaf__0459_ _0992_/a_1059_315# 0.0204f
C54216 net66 acc0.A\[9\] 0.23187f
C54217 _0559_/a_245_297# net26 0
C54218 _0411_ net5 0.29127f
C54219 hold31/a_49_47# _0086_ 0
C54220 _0407_ _0219_ 0.06436f
C54221 _0982_/a_381_47# acc0.A\[0\] 0.01346f
C54222 net245 _0997_/a_1059_315# 0
C54223 _0174_ _0542_/a_240_47# 0.01387f
C54224 VPWR _1065_/a_561_413# 0.00233f
C54225 _1012_/a_27_47# hold92/a_285_47# 0
C54226 _1012_/a_193_47# hold92/a_49_47# 0
C54227 _0107_ _0462_ 0.00132f
C54228 _0247_ _0774_/a_150_297# 0.00151f
C54229 _0343_ clkload4/a_268_47# 0
C54230 net123 _1037_/a_1017_47# 0
C54231 _1056_/a_27_47# net142 0.22482f
C54232 clknet_1_1__leaf_clk _0471_ 0.03234f
C54233 _0353_ acc0.A\[29\] 0.06031f
C54234 _0995_/a_193_47# _0995_/a_381_47# 0.09972f
C54235 _0995_/a_634_159# _0995_/a_891_413# 0.03684f
C54236 _0995_/a_27_47# _0995_/a_561_413# 0.0027f
C54237 _0529_/a_373_47# net170 0.00245f
C54238 _0413_ _0277_ 0
C54239 _0443_ _0432_ 0.19228f
C54240 _0365_ _0321_ 0
C54241 _0091_ _0418_ 0
C54242 _0119_ net150 0.00115f
C54243 _1002_/a_1059_315# _0382_ 0
C54244 _1060_/a_592_47# acc0.A\[15\] 0
C54245 _0983_/a_27_47# _0346_ 0.01665f
C54246 net158 comp0.B\[9\] 0
C54247 _0750_/a_27_47# net213 0
C54248 _0435_ _0434_ 0.13226f
C54249 hold87/a_49_47# _0854_/a_79_21# 0.05861f
C54250 net48 net177 0
C54251 net23 _1066_/a_27_47# 0
C54252 clknet_0_clk _1065_/a_27_47# 0.01237f
C54253 net32 _1042_/a_193_47# 0.05082f
C54254 _0205_ _1042_/a_1059_315# 0
C54255 net152 _1042_/a_634_159# 0
C54256 input4/a_75_212# _0511_/a_81_21# 0
C54257 hold57/a_49_47# net204 0
C54258 net53 _1007_/a_975_413# 0.00141f
C54259 _0227_ hold66/a_285_47# 0
C54260 acc0.A\[21\] hold66/a_391_47# 0.00202f
C54261 _1070_/a_891_413# _1069_/a_891_413# 0.00175f
C54262 _0289_ _0346_ 0.18597f
C54263 control0.state\[0\] _1062_/a_381_47# 0.00123f
C54264 control0.state\[1\] _1062_/a_891_413# 0.00283f
C54265 _0982_/a_193_47# _0183_ 0.02496f
C54266 _0982_/a_466_413# _0217_ 0
C54267 _1034_/a_193_47# _0473_ 0
C54268 _0954_/a_32_297# _1045_/a_1059_315# 0.00659f
C54269 hold74/a_285_47# _0115_ 0
C54270 pp[28] hold95/a_49_47# 0
C54271 clknet_1_1__leaf__0463_ _0562_/a_68_297# 0
C54272 hold25/a_49_47# A[1] 0
C54273 clkbuf_1_0__f__0465_/a_110_47# _0825_/a_68_297# 0.00186f
C54274 acc0.A\[30\] hold62/a_49_47# 0
C54275 net167 _0166_ 0
C54276 _1011_/a_466_413# _1011_/a_561_413# 0.00772f
C54277 _1011_/a_634_159# _1011_/a_975_413# 0
C54278 _0608_/a_27_47# _0347_ 0.0034f
C54279 net50 _1023_/a_891_413# 0
C54280 VPWR _0087_ 0.35779f
C54281 _0133_ _1034_/a_466_413# 0.00902f
C54282 hold29/a_285_47# acc0.A\[23\] 0.02033f
C54283 net133 _0181_ 0.18198f
C54284 clkload2/a_110_47# net170 0
C54285 acc0.A\[9\] _0350_ 0.02188f
C54286 _0205_ net10 0
C54287 _0247_ _0773_/a_35_297# 0
C54288 _0350_ _1006_/a_592_47# 0.00282f
C54289 _0195_ net207 0.02248f
C54290 net45 _0997_/a_1059_315# 0.00203f
C54291 _0272_ _0218_ 0
C54292 acc0.A\[12\] _0280_ 0.28746f
C54293 _0425_ _0089_ 0.21708f
C54294 _0423_ net67 0.0215f
C54295 hold14/a_285_47# clknet_1_0__leaf__0463_ 0
C54296 _0216_ _1025_/a_193_47# 0
C54297 _1030_/a_27_47# net116 0.22113f
C54298 _1055_/a_466_413# VPWR 0.26559f
C54299 _1018_/a_27_47# clknet_1_0__leaf__0461_ 0.04762f
C54300 _0352_ net90 0.30286f
C54301 _1020_/a_1017_47# VPWR 0
C54302 _1001_/a_27_47# _0242_ 0
C54303 _1001_/a_634_159# acc0.A\[19\] 0
C54304 _0577_/a_27_297# net49 0.00223f
C54305 _1003_/a_634_159# VPWR 0.19682f
C54306 _0251_ _0828_/a_199_47# 0
C54307 _0857_/a_27_47# net118 0
C54308 _0181_ _1063_/a_891_413# 0
C54309 _0837_/a_368_297# _0218_ 0.00126f
C54310 net9 _0527_/a_27_297# 0.00893f
C54311 clknet_0__0464_ _1049_/a_193_47# 0.01473f
C54312 net35 _1068_/a_27_47# 0
C54313 comp0.B\[3\] comp0.B\[6\] 0.28011f
C54314 VPWR net181 0.13112f
C54315 output67/a_27_47# net4 0
C54316 _0216_ hold95/a_285_47# 0.00167f
C54317 hold44/a_391_47# _0127_ 0.05487f
C54318 _0404_ _0300_ 0.30428f
C54319 _0585_/a_27_297# _0181_ 0.11053f
C54320 _0299_ _0297_ 0.77062f
C54321 net148 _0987_/a_27_47# 0.1188f
C54322 _0305_ _0218_ 0.03852f
C54323 _0225_ hold94/a_49_47# 0
C54324 _0349_ _0218_ 0
C54325 _0733_/a_222_93# clknet_0__0462_ 0.00572f
C54326 _0293_ _0427_ 0
C54327 acc0.A\[7\] _0435_ 0.00515f
C54328 net65 _0436_ 0.00136f
C54329 _0435_ _0989_/a_1059_315# 0.00107f
C54330 clkbuf_1_0__f__0458_/a_110_47# _0637_/a_56_297# 0
C54331 _1023_/a_193_47# _1023_/a_634_159# 0.12729f
C54332 _1023_/a_27_47# _1023_/a_466_413# 0.27314f
C54333 _0343_ net239 0
C54334 _0183_ _0450_ 0
C54335 VPWR _0799_/a_80_21# 0.14755f
C54336 net9 hold1/a_391_47# 0
C54337 _1042_/a_634_159# _1042_/a_466_413# 0.23992f
C54338 _1042_/a_193_47# _1042_/a_1059_315# 0.03405f
C54339 _1042_/a_27_47# _1042_/a_891_413# 0.03089f
C54340 hold100/a_49_47# acc0.A\[15\] 0.01459f
C54341 _0181_ _1060_/a_891_413# 0.05475f
C54342 net165 net221 0
C54343 net54 net94 0
C54344 hold85/a_49_47# _0467_ 0
C54345 hold12/a_285_47# clknet_0_clk 0.00216f
C54346 _0255_ _0150_ 0.00179f
C54347 clknet_0__0457_ net105 0.07073f
C54348 _1010_/a_891_413# _0352_ 0.01137f
C54349 _0982_/a_193_47# acc0.A\[15\] 0
C54350 _0734_/a_47_47# _0317_ 0
C54351 _1045_/a_891_413# _0540_/a_51_297# 0
C54352 _0459_ _0507_/a_109_47# 0
C54353 _0531_/a_373_47# _0465_ 0
C54354 acc0.A\[27\] _0350_ 0.00105f
C54355 net176 net52 0
C54356 _0119_ control0.add 0.1941f
C54357 _0179_ _1050_/a_634_159# 0.01758f
C54358 hold63/a_391_47# _0124_ 0.01517f
C54359 _0413_ _0298_ 0.06226f
C54360 _0412_ _0299_ 0
C54361 _0800_/a_512_297# _0219_ 0.00229f
C54362 _0347_ _0841_/a_297_297# 0
C54363 _0470_ net231 0.28603f
C54364 _1036_/a_27_47# net161 0.10478f
C54365 _1036_/a_1059_315# _1036_/a_1017_47# 0
C54366 clknet_1_1__leaf__0459_ _0421_ 0.0031f
C54367 _0714_/a_149_47# _0339_ 0.0014f
C54368 _0346_ _0990_/a_592_47# 0
C54369 hold69/a_285_47# net52 0.0598f
C54370 control0.sh _0563_/a_240_47# 0
C54371 output59/a_27_47# net209 0
C54372 pp[30] hold62/a_391_47# 0.00561f
C54373 net10 _1042_/a_193_47# 0.03404f
C54374 _0153_ _0988_/a_27_47# 0
C54375 clknet_0__0459_ _0346_ 0
C54376 _0644_/a_285_47# _0276_ 0.04395f
C54377 _0693_/a_68_297# acc0.A\[23\] 0
C54378 VPWR _1040_/a_466_413# 0.24826f
C54379 _0992_/a_27_47# clknet_1_1__leaf__0465_ 0.011f
C54380 _0891_/a_27_47# net157 0
C54381 _0129_ _0567_/a_109_297# 0.00417f
C54382 hold27/a_391_47# net7 0.06703f
C54383 comp0.B\[7\] net204 0
C54384 _0449_ _0350_ 0.39374f
C54385 _0227_ _0183_ 0.01978f
C54386 _0410_ acc0.A\[15\] 0.02537f
C54387 _0366_ _0758_/a_215_47# 0
C54388 control0.reset _0564_/a_68_297# 0.00199f
C54389 pp[10] _0188_ 0
C54390 _1036_/a_27_47# net26 0
C54391 hold88/a_49_47# output47/a_27_47# 0
C54392 _1011_/a_634_159# _0334_ 0
C54393 control0.count\[3\] _0490_ 0.00263f
C54394 hold49/a_49_47# _0141_ 0.31275f
C54395 clknet_1_0__leaf__0458_ _0986_/a_27_47# 0
C54396 _1002_/a_27_47# _0765_/a_215_47# 0
C54397 clkload4/Y clknet_1_1__leaf__0461_ 0.00161f
C54398 _0305_ _0775_/a_215_47# 0
C54399 _0617_/a_68_297# net52 0
C54400 _0256_ _0444_ 0
C54401 clknet_1_0__leaf__0462_ _1024_/a_975_413# 0
C54402 _0467_ _1063_/a_975_413# 0
C54403 _1058_/a_891_413# _0187_ 0
C54404 _0450_ acc0.A\[15\] 0.03499f
C54405 _0178_ clkbuf_1_1__f__0457_/a_110_47# 0.02417f
C54406 hold59/a_391_47# _0399_ 0.02067f
C54407 _0459_ _0242_ 0.0592f
C54408 clknet_1_1__leaf__0460_ hold90/a_285_47# 0
C54409 _1021_/a_561_413# _0181_ 0
C54410 _1032_/a_466_413# _1067_/a_27_47# 0
C54411 _1032_/a_634_159# _1067_/a_193_47# 0
C54412 _1032_/a_27_47# _1067_/a_466_413# 0
C54413 _1052_/a_27_47# net15 0
C54414 pp[0] net124 0.00247f
C54415 _0777_/a_285_47# _0395_ 0.0478f
C54416 clknet_1_1__leaf_clk control0.reset 0.21915f
C54417 _0368_ net93 0
C54418 _0646_/a_47_47# _0093_ 0
C54419 _0083_ net58 0
C54420 _1012_/a_381_47# net239 0
C54421 _0428_ _0990_/a_1017_47# 0
C54422 clknet_0__0458_ _0347_ 0.0037f
C54423 _0382_ net91 0.0023f
C54424 _0110_ _0350_ 0
C54425 _0217_ _0393_ 0
C54426 _1054_/a_1059_315# net65 0
C54427 _1054_/a_466_413# acc0.A\[7\] 0
C54428 _0257_ _0438_ 0
C54429 _0346_ _0655_/a_109_93# 0.00446f
C54430 _0618_/a_79_21# net51 0.04618f
C54431 net197 hold8/a_391_47# 0
C54432 net190 hold8/a_49_47# 0
C54433 clkbuf_1_1__f__0463_/a_110_47# _1033_/a_466_413# 0
C54434 clknet_0__0463_ _1033_/a_27_47# 0
C54435 _0680_/a_217_297# _0246_ 0
C54436 _0803_/a_68_297# _0345_ 0
C54437 clknet_1_0__leaf__0464_ _1049_/a_27_47# 0.07905f
C54438 hold41/a_49_47# input2/a_75_212# 0.00138f
C54439 _0984_/a_27_47# net77 0
C54440 net70 _0991_/a_27_47# 0
C54441 _0736_/a_56_297# _0219_ 0.07679f
C54442 _0675_/a_150_297# _0218_ 0.00145f
C54443 _0457_ _0565_/a_245_297# 0
C54444 _0279_ _0788_/a_68_297# 0.18343f
C54445 _1053_/a_634_159# _1052_/a_634_159# 0
C54446 _1053_/a_193_47# _1052_/a_466_413# 0
C54447 _1053_/a_466_413# _1052_/a_193_47# 0
C54448 clknet_1_1__leaf__0459_ _0809_/a_81_21# 0
C54449 _0156_ _0281_ 0.00231f
C54450 _0217_ _0758_/a_79_21# 0
C54451 _0257_ _0636_/a_59_75# 0
C54452 _0550_/a_51_297# _1040_/a_634_159# 0
C54453 _0093_ _0995_/a_381_47# 0.11464f
C54454 _0643_/a_337_297# _0256_ 0
C54455 _0643_/a_253_47# _0270_ 0
C54456 VPWR A[3] 0.32313f
C54457 net170 _0148_ 0
C54458 net208 _0219_ 0.00178f
C54459 _0992_/a_1059_315# _0655_/a_215_53# 0
C54460 _0322_ _0462_ 0
C54461 _0346_ _0418_ 0
C54462 _0673_/a_337_297# _0345_ 0
C54463 _1055_/a_381_47# clknet_1_1__leaf__0465_ 0.01255f
C54464 _0672_/a_215_47# _0345_ 0.00156f
C54465 hold11/a_391_47# clknet_1_0__leaf__0465_ 0.01183f
C54466 _0191_ net148 0
C54467 net120 _0208_ 0
C54468 _0779_/a_510_47# _0352_ 0.00295f
C54469 _0327_ _0462_ 0.09988f
C54470 net160 net25 0
C54471 clkbuf_0_clk/a_110_47# _1068_/a_193_47# 0.00231f
C54472 net170 _0845_/a_109_47# 0
C54473 _0673_/a_253_47# _0304_ 0.01528f
C54474 _0728_/a_59_75# net208 0
C54475 _0186_ hold83/a_49_47# 0
C54476 _1038_/a_27_47# _0207_ 0
C54477 _1038_/a_193_47# net171 0
C54478 _0304_ _0672_/a_510_47# 0
C54479 _1051_/a_634_159# _0524_/a_109_297# 0
C54480 _1051_/a_466_413# _0524_/a_27_297# 0
C54481 _0461_ VPWR 1.27948f
C54482 net248 acc0.A\[8\] 0
C54483 VPWR _0703_/a_109_297# 0.00653f
C54484 _0081_ _0849_/a_79_21# 0
C54485 _0854_/a_79_21# _0082_ 0
C54486 _0455_ _0849_/a_215_47# 0
C54487 _0992_/a_891_413# _0281_ 0
C54488 _1046_/a_891_413# _0142_ 0
C54489 _0845_/a_109_297# _0845_/a_109_47# 0
C54490 _1053_/a_466_413# net12 0.01045f
C54491 _0243_ hold76/a_49_47# 0
C54492 _0389_ hold76/a_285_47# 0.00366f
C54493 _0734_/a_377_297# clknet_1_1__leaf__0460_ 0
C54494 net70 _0350_ 0.00281f
C54495 acc0.A\[18\] _0345_ 0
C54496 _0189_ _0369_ 0
C54497 VPWR _0318_ 0.70121f
C54498 net224 _0219_ 0.03667f
C54499 _0530_/a_384_47# _0186_ 0
C54500 VPWR _0994_/a_466_413# 0.26198f
C54501 _0343_ _1060_/a_27_47# 0.00171f
C54502 _1039_/a_27_47# _0175_ 0
C54503 net118 net107 0
C54504 _0179_ net62 0
C54505 _0981_/a_373_47# clknet_0_clk 0
C54506 clknet_1_0__leaf__0462_ _0367_ 0.08811f
C54507 output60/a_27_47# net41 0
C54508 _0195_ hold72/a_285_47# 0
C54509 _0229_ _0217_ 0
C54510 _0179_ _0450_ 0.02125f
C54511 _0461_ _1015_/a_466_413# 0.00857f
C54512 hold75/a_49_47# _0219_ 0.05011f
C54513 _1010_/a_193_47# _0350_ 0.46865f
C54514 pp[27] _1011_/a_193_47# 0
C54515 _0601_/a_68_297# _0601_/a_150_297# 0.00477f
C54516 _0399_ _0830_/a_297_297# 0
C54517 _0576_/a_109_47# net176 0.00201f
C54518 _0662_/a_81_21# _0990_/a_1059_315# 0
C54519 net45 _0582_/a_27_297# 0.00402f
C54520 _0222_ _1005_/a_1059_315# 0
C54521 _0339_ hold62/a_391_47# 0.02422f
C54522 hold74/a_391_47# _1017_/a_1059_315# 0
C54523 _0280_ net42 0.26563f
C54524 _0697_/a_217_297# _0697_/a_472_297# 0.00517f
C54525 _0697_/a_80_21# _0697_/a_300_47# 0.00997f
C54526 clknet_1_1__leaf__0460_ _0748_/a_81_21# 0
C54527 _0218_ _0181_ 0.06374f
C54528 net157 _0935_/a_27_47# 0.00629f
C54529 _0305_ _1017_/a_975_413# 0
C54530 hold87/a_285_47# _0195_ 0
C54531 net157 _1061_/a_193_47# 0.01126f
C54532 net14 A[6] 0.11417f
C54533 _0702_/a_113_47# _0334_ 0.00937f
C54534 hold70/a_49_47# hold70/a_285_47# 0.22264f
C54535 hold63/a_49_47# _1026_/a_193_47# 0
C54536 hold63/a_285_47# _1026_/a_27_47# 0.00319f
C54537 _0990_/a_193_47# clknet_1_1__leaf__0458_ 0
C54538 _1056_/a_27_47# _0988_/a_27_47# 0
C54539 _0369_ _0381_ 0.0314f
C54540 _0995_/a_193_47# _0219_ 0.00471f
C54541 comp0.B\[4\] _0955_/a_304_297# 0
C54542 _0521_/a_384_47# _0179_ 0
C54543 _0174_ _0544_/a_512_297# 0
C54544 _1009_/a_634_159# _0350_ 0
C54545 clknet_1_0__leaf__0462_ _0217_ 0.30925f
C54546 _0531_/a_27_297# _1047_/a_27_47# 0
C54547 _1031_/a_193_47# _1031_/a_381_47# 0.09972f
C54548 _1031_/a_634_159# _1031_/a_891_413# 0.03684f
C54549 _1031_/a_27_47# _1031_/a_561_413# 0.0027f
C54550 net86 _0459_ 0.0206f
C54551 net63 input15/a_75_212# 0
C54552 _0369_ hold72/a_49_47# 0.00992f
C54553 net31 net152 0
C54554 input31/a_75_212# _0139_ 0
C54555 B[8] net32 0
C54556 _0996_/a_1059_315# _0346_ 0
C54557 _0804_/a_510_47# _0403_ 0
C54558 _0416_ _0788_/a_68_297# 0
C54559 control0.add _0373_ 0.001f
C54560 _1000_/a_466_413# _0218_ 0
C54561 net108 net151 0
C54562 _0722_/a_79_21# _0722_/a_215_47# 0.04584f
C54563 _1005_/a_634_159# net91 0
C54564 _1005_/a_193_47# _0103_ 0.41139f
C54565 _1005_/a_891_413# _1005_/a_1017_47# 0.00617f
C54566 _0336_ _0333_ 0
C54567 _0769_/a_81_21# _0240_ 0
C54568 control0.state\[1\] _0470_ 0
C54569 acc0.A\[12\] net143 0.00898f
C54570 hold55/a_391_47# _0183_ 0
C54571 clknet_0__0458_ clkbuf_0__0465_/a_110_47# 0.02354f
C54572 comp0.B\[3\] net26 0
C54573 _0984_/a_561_413# _0082_ 0
C54574 _0151_ net12 0.10048f
C54575 _1013_/a_466_413# _1013_/a_592_47# 0.00553f
C54576 _1013_/a_634_159# _1013_/a_1017_47# 0
C54577 _0976_/a_505_21# _1069_/a_27_47# 0
C54578 _0976_/a_76_199# _1069_/a_193_47# 0
C54579 net1 _1062_/a_193_47# 0
C54580 VPWR net154 0.56208f
C54581 _1002_/a_634_159# _1002_/a_381_47# 0
C54582 _0792_/a_80_21# _0790_/a_35_297# 0.0163f
C54583 _0985_/a_193_47# hold28/a_391_47# 0
C54584 clknet_1_0__leaf__0465_ _0524_/a_109_297# 0.0055f
C54585 clknet_1_1__leaf__0460_ clknet_0__0462_ 0.00924f
C54586 _0467_ net17 0.06369f
C54587 _0640_/a_215_297# VPWR 0.13269f
C54588 _0984_/a_1059_315# clknet_1_0__leaf__0458_ 0.00909f
C54589 _0437_ acc0.A\[6\] 0.0051f
C54590 net22 _1046_/a_634_159# 0.00101f
C54591 _0310_ _0773_/a_117_297# 0
C54592 _0083_ _0262_ 0
C54593 _0583_/a_27_297# _0158_ 0.0012f
C54594 _0390_ _0461_ 0.00212f
C54595 hold28/a_49_47# _1049_/a_27_47# 0
C54596 _0965_/a_47_47# clknet_1_0__leaf_clk 0.11441f
C54597 _0154_ _1055_/a_27_47# 0
C54598 hold35/a_285_47# _1055_/a_1059_315# 0.0054f
C54599 hold87/a_285_47# _0852_/a_35_297# 0.01561f
C54600 _0372_ _0246_ 0
C54601 VPWR _0989_/a_975_413# 0.00417f
C54602 VPWR _0997_/a_1059_315# 0.41732f
C54603 _0678_/a_68_297# _0347_ 0.00343f
C54604 _0421_ _0655_/a_215_53# 0.00976f
C54605 _1059_/a_634_159# _0369_ 0.01084f
C54606 _0217_ _1019_/a_891_413# 0
C54607 _0183_ _1019_/a_466_413# 0.0065f
C54608 VPWR _0992_/a_975_413# 0.00489f
C54609 _0223_ _0232_ 0.26771f
C54610 output54/a_27_47# hold8/a_49_47# 0.00529f
C54611 hold35/a_391_47# net181 0
C54612 control0.state\[1\] _0958_/a_303_47# 0
C54613 _0354_ clknet_1_1__leaf__0462_ 0
C54614 _1035_/a_466_413# _0175_ 0.01858f
C54615 _0305_ _0359_ 0
C54616 _0765_/a_79_21# net220 0.05418f
C54617 VPWR _0465_ 1.88943f
C54618 _0170_ hold17/a_49_47# 0
C54619 VPWR _1061_/a_381_47# 0.07852f
C54620 net17 comp0.B\[0\] 0.00766f
C54621 net214 clkbuf_1_1__f__0465_/a_110_47# 0.00503f
C54622 _1015_/a_1059_315# control0.reset 0
C54623 clknet_1_0__leaf__0463_ _1046_/a_634_159# 0
C54624 _0195_ _0392_ 0
C54625 net82 acc0.A\[13\] 0.00427f
C54626 _1034_/a_561_413# _0213_ 0.00114f
C54627 _1034_/a_381_47# _0173_ 0.00334f
C54628 _1034_/a_193_47# _0132_ 0.01286f
C54629 acc0.A\[2\] VPWR 1.47918f
C54630 clkbuf_1_0__f__0465_/a_110_47# net148 0
C54631 net211 _0345_ 0.45818f
C54632 hold87/a_285_47# _0081_ 0
C54633 _0217_ net206 0.70361f
C54634 _0183_ net219 0.51956f
C54635 _1035_/a_1059_315# control0.sh 0.01185f
C54636 hold9/a_391_47# net156 0.1415f
C54637 A[12] _0156_ 0
C54638 _1018_/a_1017_47# _0459_ 0
C54639 _1070_/a_1059_315# control0.count\[0\] 0.00116f
C54640 control0.count\[1\] _1069_/a_1059_315# 0.07147f
C54641 VPWR _1069_/a_592_47# 0
C54642 _0327_ _0725_/a_303_47# 0
C54643 _0985_/a_193_47# _0218_ 0
C54644 net53 hold53/a_285_47# 0.03949f
C54645 _0080_ _0217_ 0
C54646 hold18/a_285_47# _0264_ 0.00212f
C54647 _0096_ _0219_ 0
C54648 _1018_/a_27_47# _0218_ 0
C54649 _1030_/a_891_413# _0705_/a_59_75# 0
C54650 _1030_/a_27_47# _0220_ 0
C54651 _1018_/a_193_47# _0294_ 0
C54652 clkbuf_1_0__f__0458_/a_110_47# _0849_/a_79_21# 0.00102f
C54653 net44 net116 0.16328f
C54654 _0762_/a_79_21# _1005_/a_891_413# 0
C54655 _0216_ _1011_/a_193_47# 0.00532f
C54656 _1011_/a_1059_315# net57 0.10543f
C54657 _0985_/a_975_413# _0186_ 0
C54658 _1000_/a_27_47# _0245_ 0.03038f
C54659 _0525_/a_81_21# _0525_/a_384_47# 0.00138f
C54660 _0399_ _0669_/a_183_297# 0
C54661 _1055_/a_891_413# A[9] 0
C54662 clknet_0__0458_ _0824_/a_59_75# 0.00553f
C54663 _1006_/a_634_159# _1006_/a_592_47# 0
C54664 _0993_/a_193_47# net246 0
C54665 _0107_ _0312_ 0
C54666 acc0.A\[1\] _1014_/a_891_413# 0
C54667 input33/a_75_212# input26/a_75_212# 0.01252f
C54668 _0461_ clknet_1_0__leaf__0459_ 2.24592f
C54669 _0655_/a_215_53# _0809_/a_81_21# 0.01091f
C54670 _0116_ _0580_/a_109_297# 0
C54671 clknet_1_0__leaf__0460_ _0754_/a_51_297# 0.00152f
C54672 _0695_/a_80_21# _0219_ 0.02679f
C54673 _0984_/a_634_159# _0984_/a_381_47# 0
C54674 _0441_ net62 0
C54675 net21 _1043_/a_891_413# 0
C54676 _0181_ _0177_ 0
C54677 _0692_/a_113_47# _0324_ 0.00937f
C54678 _1031_/a_193_47# _0219_ 0
C54679 acc0.A\[14\] _0583_/a_27_297# 0
C54680 _0808_/a_266_297# _0417_ 0.01101f
C54681 net179 VPWR 0.32141f
C54682 net182 net181 0
C54683 _0610_/a_59_75# net223 0
C54684 acc0.A\[19\] _0772_/a_215_47# 0
C54685 acc0.A\[26\] _0687_/a_59_75# 0.13166f
C54686 net89 VPWR 0.46788f
C54687 _0550_/a_245_297# _0207_ 0
C54688 _0163_ _0161_ 0.26428f
C54689 hold66/a_285_47# _0352_ 0
C54690 output37/a_27_47# acc0.A\[11\] 0
C54691 comp0.B\[3\] hold84/a_285_47# 0
C54692 _0260_ _0350_ 0.09706f
C54693 _1039_/a_381_47# VPWR 0.07135f
C54694 net44 hold92/a_285_47# 0.00468f
C54695 _0343_ hold19/a_391_47# 0.01668f
C54696 _0986_/a_634_159# _0986_/a_592_47# 0
C54697 _0112_ _0181_ 0.01055f
C54698 _1056_/a_975_413# _0153_ 0
C54699 net242 _0354_ 0
C54700 _0856_/a_215_47# _0264_ 0.04611f
C54701 _1017_/a_975_413# _0181_ 0
C54702 _1023_/a_1059_315# _1023_/a_1017_47# 0
C54703 _1023_/a_193_47# net109 0.00707f
C54704 _1023_/a_27_47# net177 0.09799f
C54705 net1 _0782_/a_27_47# 0.00983f
C54706 net46 _0869_/a_27_47# 0.00101f
C54707 _0247_ _1006_/a_27_47# 0
C54708 clknet_0__0461_ _0240_ 0.00244f
C54709 _0294_ _0816_/a_68_297# 0.00157f
C54710 _1037_/a_27_47# _0175_ 0
C54711 _0948_/a_109_297# VPWR 0.0044f
C54712 hold49/a_285_47# net18 0
C54713 _0369_ clknet_0__0461_ 0.20447f
C54714 hold38/a_49_47# _0487_ 0
C54715 net54 _0328_ 0
C54716 _0495_/a_68_297# _0495_/a_150_297# 0.00477f
C54717 clknet_1_0__leaf__0458_ hold18/a_49_47# 0.01268f
C54718 _0313_ _0216_ 0
C54719 _0662_/a_81_21# VPWR 0.21727f
C54720 net23 _0584_/a_27_297# 0.18103f
C54721 control0.state\[0\] _0946_/a_30_53# 0.13649f
C54722 clknet_1_1__leaf__0464_ _1044_/a_592_47# 0.00114f
C54723 VPWR hold4/a_49_47# 0.2676f
C54724 hold9/a_391_47# acc0.A\[26\] 0.002f
C54725 _1037_/a_193_47# control0.sh 0.00228f
C54726 _0438_ clknet_1_1__leaf__0458_ 0.75614f
C54727 _0718_/a_47_47# hold62/a_391_47# 0
C54728 _0093_ _0219_ 0.00866f
C54729 net150 _0761_/a_113_47# 0
C54730 net125 _0171_ 0.00206f
C54731 net243 _0350_ 0.36446f
C54732 _0592_/a_68_297# _0222_ 0.01782f
C54733 _0195_ _0196_ 0.00938f
C54734 net71 _0219_ 0.00123f
C54735 net133 _0531_/a_27_297# 0.00114f
C54736 _0129_ _1031_/a_27_47# 0.00639f
C54737 hold16/a_391_47# _1031_/a_466_413# 0
C54738 hold16/a_49_47# _1031_/a_891_413# 0
C54739 _0305_ net228 0.02711f
C54740 _0216_ net202 0.00292f
C54741 _0230_ net213 0.00526f
C54742 _0710_/a_381_47# _0216_ 0
C54743 _0616_/a_78_199# _0616_/a_292_297# 0.01295f
C54744 net208 hold61/a_49_47# 0
C54745 _0404_ _0419_ 0
C54746 _1059_/a_27_47# net229 0.04216f
C54747 hold22/a_49_47# acc0.A\[7\] 0.06804f
C54748 hold31/a_49_47# _0621_/a_35_297# 0.00533f
C54749 net165 _0446_ 0.11078f
C54750 net61 net75 0
C54751 net123 _0555_/a_51_297# 0
C54752 _1057_/a_193_47# _0156_ 0
C54753 _1038_/a_27_47# _1037_/a_1059_315# 0
C54754 _1038_/a_466_413# _1037_/a_193_47# 0
C54755 _1038_/a_634_159# _1037_/a_634_159# 0
C54756 _1038_/a_193_47# _1037_/a_466_413# 0
C54757 hold77/a_391_47# _0219_ 0.00542f
C54758 _0346_ _0462_ 0.13706f
C54759 _0732_/a_209_297# net51 0
C54760 VPWR net174 1.17714f
C54761 net193 _0544_/a_51_297# 0
C54762 _0981_/a_109_47# _0488_ 0
C54763 _0981_/a_109_297# _0466_ 0.01982f
C54764 _0997_/a_27_47# _0095_ 0.09664f
C54765 _0997_/a_891_413# _0407_ 0
C54766 net118 _0208_ 0
C54767 _0324_ _0618_/a_79_21# 0
C54768 _0855_/a_81_21# _0265_ 0.00155f
C54769 net234 _0633_/a_109_297# 0.00324f
C54770 net240 _0181_ 0.04138f
C54771 acc0.A\[4\] _0194_ 0
C54772 clknet_1_0__leaf__0458_ _0856_/a_297_297# 0
C54773 _0837_/a_81_21# clkbuf_1_0__f__0465_/a_110_47# 0
C54774 net97 _0334_ 0
C54775 net42 output41/a_27_47# 0
C54776 _0770_/a_79_21# clknet_1_0__leaf__0457_ 0.00103f
C54777 net88 _0765_/a_79_21# 0
C54778 _0777_/a_129_47# _0394_ 0.00125f
C54779 _1002_/a_381_47# net220 0
C54780 net55 _0349_ 0
C54781 _0143_ net9 0
C54782 hold30/a_391_47# _0217_ 0.05866f
C54783 hold30/a_49_47# _0183_ 0.04331f
C54784 hold30/a_285_47# acc0.A\[22\] 0.02208f
C54785 _0363_ _0308_ 0
C54786 _0571_/a_109_297# acc0.A\[27\] 0.01055f
C54787 clkbuf_0__0464_/a_110_47# net157 0.00119f
C54788 _0532_/a_81_21# _0532_/a_384_47# 0.00138f
C54789 hold85/a_49_47# net1 0
C54790 net58 _0088_ 0
C54791 _0743_/a_512_297# _0219_ 0.00125f
C54792 _0999_/a_1017_47# _0218_ 0.00125f
C54793 clknet_1_1__leaf__0463_ _1067_/a_27_47# 0.00865f
C54794 clknet_0__0460_ net93 0
C54795 _0637_/a_56_297# acc0.A\[15\] 0.00509f
C54796 net169 acc0.A\[7\] 0.23957f
C54797 _0664_/a_79_21# _0282_ 0
C54798 _0627_/a_109_93# clkbuf_0__0465_/a_110_47# 0
C54799 _0359_ _0181_ 0
C54800 _0238_ _0749_/a_299_297# 0
C54801 clkbuf_1_1__f__0463_/a_110_47# _0131_ 0.03347f
C54802 net133 _1049_/a_592_47# 0
C54803 net32 clknet_1_1__leaf__0464_ 0
C54804 VPWR _0582_/a_27_297# 0.27447f
C54805 hold38/a_49_47# net119 0.00209f
C54806 VPWR _1007_/a_27_47# 0.72847f
C54807 VPWR _1035_/a_592_47# 0
C54808 _0137_ _1040_/a_27_47# 0
C54809 net180 _1040_/a_1059_315# 0.00132f
C54810 _0172_ _1040_/a_634_159# 0.00313f
C54811 _0183_ _0352_ 0.08989f
C54812 _1058_/a_634_159# VPWR 0.18357f
C54813 net236 _0981_/a_109_297# 0
C54814 _0345_ net241 0.24954f
C54815 VPWR B[15] 0.22275f
C54816 _0982_/a_975_413# _0181_ 0
C54817 net171 net29 0.28594f
C54818 _0669_/a_29_53# _0345_ 0.00952f
C54819 _1055_/a_891_413# _0516_/a_27_297# 0
C54820 _1055_/a_1059_315# _0516_/a_109_297# 0
C54821 _1064_/a_1059_315# _1064_/a_891_413# 0.31086f
C54822 _1064_/a_193_47# _1064_/a_975_413# 0
C54823 _1064_/a_466_413# _1064_/a_381_47# 0.03733f
C54824 _0234_ _0750_/a_109_47# 0
C54825 _0294_ clknet_0__0460_ 0
C54826 _0218_ clknet_1_1__leaf__0461_ 0.78958f
C54827 clknet_1_1__leaf_clk _1063_/a_193_47# 0.0137f
C54828 _0707_/a_201_297# _0334_ 0.01241f
C54829 _0346_ _0297_ 0.00136f
C54830 _0672_/a_297_297# _0301_ 0
C54831 hold97/a_285_47# _0350_ 0
C54832 _0473_ _0171_ 0
C54833 _0386_ _0771_/a_215_297# 0
C54834 _0388_ _0771_/a_27_413# 0
C54835 _0786_/a_80_21# VPWR 0.2207f
C54836 _0694_/a_113_47# acc0.A\[24\] 0
C54837 _0770_/a_79_21# _1001_/a_1059_315# 0.00105f
C54838 _0100_ net187 0
C54839 clkbuf_1_0__f__0459_/a_110_47# _1060_/a_27_47# 0.01237f
C54840 _0166_ _1063_/a_27_47# 0
C54841 _0149_ _0524_/a_27_297# 0.02142f
C54842 _1051_/a_466_413# _0194_ 0
C54843 _0316_ _0701_/a_80_21# 0
C54844 _0983_/a_891_413# _0582_/a_109_297# 0
C54845 _0343_ _1017_/a_466_413# 0
C54846 _1002_/a_193_47# _0369_ 0
C54847 _0752_/a_27_413# _0227_ 0.05607f
C54848 _0521_/a_299_297# hold83/a_285_47# 0
C54849 net24 net29 0
C54850 _0626_/a_68_297# _0624_/a_59_75# 0.00101f
C54851 net1 _0585_/a_373_47# 0.00271f
C54852 comp0.B\[14\] hold6/a_391_47# 0
C54853 _0467_ _0165_ 0
C54854 hold41/a_49_47# _0512_/a_109_297# 0
C54855 hold41/a_285_47# _0512_/a_27_297# 0.00129f
C54856 clknet_1_1__leaf_clk _0460_ 0.01108f
C54857 control0.state\[0\] _0967_/a_109_93# 0.02375f
C54858 _0598_/a_297_47# _0374_ 0
C54859 net34 _0484_ 0.03407f
C54860 control0.state\[0\] _0487_ 0.62154f
C54861 control0.state\[1\] _0485_ 0
C54862 _0701_/a_80_21# _0347_ 0.00526f
C54863 clknet_1_0__leaf__0458_ _0455_ 0.0045f
C54864 clknet_0__0465_ _0444_ 0.00231f
C54865 _1017_/a_634_159# acc0.A\[17\] 0.00229f
C54866 _0461_ _0113_ 0.00901f
C54867 _0457_ _0564_/a_68_297# 0
C54868 output39/a_27_47# net5 0
C54869 output55/a_27_47# net57 0.02879f
C54870 _0412_ _0346_ 0
C54871 _1008_/a_193_47# _0345_ 0
C54872 comp0.B\[2\] _0959_/a_80_21# 0
C54873 _0737_/a_285_297# _0364_ 0.07187f
C54874 net45 _0115_ 0.00626f
C54875 _0854_/a_215_47# _0854_/a_510_47# 0.00529f
C54876 clknet_1_1__leaf__0464_ _1042_/a_1059_315# 0
C54877 hold2/a_285_47# hold2/a_391_47# 0.41909f
C54878 VPWR clknet_0__0464_ 2.0632f
C54879 _0763_/a_193_47# net92 0
C54880 net201 _0173_ 0.14642f
C54881 hold74/a_391_47# _1016_/a_27_47# 0
C54882 hold74/a_285_47# _1016_/a_193_47# 0
C54883 _0252_ acc0.A\[6\] 0.06276f
C54884 _0305_ _1016_/a_1059_315# 0.00364f
C54885 _0217_ _0574_/a_373_47# 0
C54886 _0229_ _0235_ 0
C54887 clkbuf_1_1__f_clk/a_110_47# _1063_/a_634_159# 0
C54888 _0457_ clknet_1_1__leaf_clk 0.00609f
C54889 _0204_ _0543_/a_68_297# 0.12411f
C54890 _0800_/a_240_47# _0997_/a_466_413# 0
C54891 _0712_/a_79_21# _0129_ 0.04524f
C54892 hold36/a_391_47# net183 0.13562f
C54893 hold36/a_285_47# net21 0
C54894 _0165_ comp0.B\[0\] 0
C54895 _0627_/a_109_93# _0824_/a_59_75# 0
C54896 hold6/a_49_47# net153 0
C54897 _0787_/a_209_297# VPWR 0.22159f
C54898 _0179_ _0812_/a_510_47# 0.00217f
C54899 _0174_ _0140_ 0
C54900 _1015_/a_27_47# clknet_1_0__leaf__0461_ 0.00747f
C54901 _0719_/a_27_47# net46 0.0015f
C54902 _0312_ _0327_ 0.00481f
C54903 _0429_ _0829_/a_27_47# 0.03802f
C54904 _0180_ net7 0
C54905 net8 net247 0
C54906 _0179_ _0514_/a_109_297# 0.01072f
C54907 clknet_1_0__leaf__0465_ _1052_/a_1059_315# 0.00459f
C54908 _0643_/a_337_297# clknet_0__0465_ 0
C54909 _1038_/a_193_47# _0553_/a_51_297# 0
C54910 _0675_/a_68_297# _0347_ 0
C54911 _1037_/a_381_47# VPWR 0.07618f
C54912 net46 _0460_ 0.04018f
C54913 _0557_/a_51_297# _0557_/a_245_297# 0.01218f
C54914 net61 _0442_ 0
C54915 net10 clknet_1_1__leaf__0464_ 0.02899f
C54916 net7 net152 0
C54917 _0255_ hold1/a_391_47# 0.04096f
C54918 net40 input5/a_75_212# 0.01791f
C54919 _1041_/a_592_47# VPWR 0
C54920 _0402_ hold81/a_49_47# 0.00332f
C54921 _0366_ _0350_ 0
C54922 _0489_ _0976_/a_505_21# 0
C54923 _0098_ _0218_ 0.00336f
C54924 pp[15] _0995_/a_975_413# 0
C54925 _0217_ _0773_/a_35_297# 0
C54926 _0722_/a_510_47# _0110_ 0
C54927 _0226_ _0603_/a_150_297# 0
C54928 net28 _0176_ 0.01994f
C54929 hold24/a_391_47# net8 0.04913f
C54930 _1048_/a_193_47# _0196_ 0
C54931 hold43/a_49_47# hold44/a_285_47# 0.03151f
C54932 _0835_/a_493_297# _0465_ 0
C54933 control0.sh _1062_/a_193_47# 0
C54934 clknet_1_1__leaf_clk _1062_/a_891_413# 0.01031f
C54935 _1056_/a_891_413# pp[9] 0
C54936 _1018_/a_634_159# _0581_/a_27_297# 0
C54937 net146 acc0.A\[13\] 0
C54938 VPWR _0831_/a_117_297# 0.00563f
C54939 _0488_ _1069_/a_193_47# 0
C54940 _0466_ _1069_/a_27_47# 0
C54941 _0401_ _0841_/a_215_47# 0
C54942 _1021_/a_466_413# clknet_1_1__leaf_clk 0
C54943 hold16/a_285_47# hold16/a_391_47# 0.41909f
C54944 pp[27] _0707_/a_75_199# 0.00858f
C54945 hold91/a_49_47# hold91/a_391_47# 0.00188f
C54946 _1002_/a_891_413# _0100_ 0.05367f
C54947 _1002_/a_381_47# net88 0.02207f
C54948 _1020_/a_193_47# _1020_/a_891_413# 0.19489f
C54949 _1020_/a_27_47# _1020_/a_381_47# 0.06222f
C54950 _1020_/a_634_159# _1020_/a_1059_315# 0
C54951 acc0.A\[23\] _0754_/a_240_47# 0
C54952 _0408_ _0790_/a_117_297# 0
C54953 _0792_/a_209_47# _0406_ 0.00108f
C54954 pp[16] pp[18] 0.00103f
C54955 net156 _0739_/a_215_47# 0.00104f
C54956 hold12/a_49_47# hold12/a_391_47# 0.00188f
C54957 _0083_ hold28/a_49_47# 0
C54958 _1021_/a_1017_47# net1 0
C54959 _0102_ _0379_ 0
C54960 _0254_ VPWR 0.80116f
C54961 clkbuf_1_0__f__0464_/a_110_47# _1049_/a_27_47# 0.01273f
C54962 _0747_/a_79_21# clkbuf_1_0__f__0460_/a_110_47# 0.00537f
C54963 _0983_/a_1059_315# net47 0.13535f
C54964 control0.count\[3\] control0.count\[0\] 0.00466f
C54965 _0589_/a_113_47# _0221_ 0.00963f
C54966 _0984_/a_1059_315# _0455_ 0
C54967 _0984_/a_891_413# _0454_ 0
C54968 _1028_/a_27_47# hold50/a_285_47# 0.01524f
C54969 _1028_/a_193_47# hold50/a_49_47# 0.00269f
C54970 hold35/a_391_47# net179 0
C54971 _1058_/a_891_413# clknet_1_1__leaf__0465_ 0.00181f
C54972 net117 net99 0
C54973 _0559_/a_51_297# _0957_/a_32_297# 0.00473f
C54974 net145 _0369_ 0
C54975 _0259_ _0785_/a_384_47# 0.01022f
C54976 _0183_ net207 0.00114f
C54977 _0747_/a_79_21# _0250_ 0.04949f
C54978 _0182_ _1048_/a_891_413# 0
C54979 _0180_ _1048_/a_1059_315# 0.00342f
C54980 _0998_/a_27_47# _1017_/a_1059_315# 0
C54981 _1001_/a_381_47# net46 0
C54982 _0457_ _0584_/a_109_47# 0
C54983 _0274_ clkbuf_1_1__f__0458_/a_110_47# 0.02412f
C54984 _0217_ _1025_/a_891_413# 0
C54985 _0133_ _0175_ 0.41265f
C54986 _0337_ hold95/a_285_47# 0
C54987 _0483_ _0974_/a_79_199# 0
C54988 _0846_/a_51_297# _0845_/a_109_47# 0
C54989 _0664_/a_297_47# VPWR 0.00702f
C54990 net40 pp[12] 0.00396f
C54991 hold94/a_285_47# _0754_/a_51_297# 0
C54992 _0545_/a_68_297# _1040_/a_891_413# 0
C54993 _0352_ hold40/a_285_47# 0.05243f
C54994 net44 _0220_ 0.08424f
C54995 comp0.B\[2\] _0173_ 0.24504f
C54996 _0622_/a_109_47# _0253_ 0
C54997 _0558_/a_68_297# _0175_ 0.1031f
C54998 _1036_/a_466_413# net24 0
C54999 _0216_ _0232_ 0
C55000 _0856_/a_79_21# hold18/a_285_47# 0
C55001 _1072_/a_27_47# _0468_ 0
C55002 _1016_/a_891_413# _0675_/a_68_297# 0
C55003 _0098_ _0775_/a_215_47# 0.00305f
C55004 _1000_/a_975_413# _0393_ 0
C55005 _1058_/a_27_47# _1057_/a_27_47# 0.02074f
C55006 VPWR _0705_/a_145_75# 0
C55007 clknet_1_0__leaf__0463_ hold5/a_391_47# 0
C55008 _0343_ _0094_ 0.00454f
C55009 comp0.B\[4\] net33 0
C55010 _0305_ _0238_ 0
C55011 comp0.B\[12\] _1044_/a_561_413# 0
C55012 _0403_ _0807_/a_68_297# 0.00183f
C55013 _0269_ _0084_ 0
C55014 _0534_/a_81_21# clknet_1_1__leaf__0457_ 0.04846f
C55015 clkbuf_0_clk/a_110_47# VPWR 1.25225f
C55016 clkbuf_0__0459_/a_110_47# _0184_ 0
C55017 net186 clknet_1_1__leaf__0463_ 0.2254f
C55018 net1 net17 0
C55019 net35 hold17/a_49_47# 0.00187f
C55020 clknet_1_0__leaf__0465_ clknet_1_1__leaf__0457_ 0.00138f
C55021 _1000_/a_634_159# _0347_ 0.0032f
C55022 _0558_/a_150_297# control0.sh 0
C55023 _1030_/a_1017_47# _0336_ 0
C55024 _0414_ _0994_/a_561_413# 0
C55025 VPWR _1063_/a_634_159# 0.18958f
C55026 _0323_ net237 0
C55027 hold66/a_285_47# _0237_ 0.01585f
C55028 _0572_/a_109_47# net155 0
C55029 _0572_/a_109_297# _0216_ 0.0068f
C55030 hold23/a_391_47# clknet_1_1__leaf__0457_ 0
C55031 _0216_ _1006_/a_561_413# 0.00132f
C55032 clknet_1_1__leaf__0458_ _0522_/a_109_297# 0
C55033 _0179_ net73 0.16345f
C55034 _0369_ net67 0.02951f
C55035 _0329_ _0219_ 0
C55036 _0330_ _0324_ 0
C55037 net182 net179 0
C55038 _0266_ _0261_ 0
C55039 _0452_ _0263_ 0
C55040 acc0.A\[26\] _0739_/a_215_47# 0.00273f
C55041 net197 hold9/a_285_47# 0.0716f
C55042 _0655_/a_369_297# _0420_ 0
C55043 clknet_1_0__leaf__0460_ _0219_ 0.22663f
C55044 pp[30] _0342_ 0
C55045 _0272_ _0268_ 0.00192f
C55046 _0984_/a_381_47# net70 0
C55047 _0352_ acc0.A\[26\] 0.10837f
C55048 _0573_/a_27_47# _0199_ 0.00157f
C55049 _0579_/a_373_47# _0461_ 0
C55050 _0236_ _0604_/a_113_47# 0.00954f
C55051 hold55/a_49_47# net118 0
C55052 clkbuf_1_0__f__0459_/a_110_47# hold19/a_391_47# 0.01183f
C55053 VPWR _1060_/a_634_159# 0.18218f
C55054 clknet_0_clk clknet_1_0__leaf_clk 0.11973f
C55055 _1019_/a_27_47# _0242_ 0
C55056 _0215_ clknet_1_0__leaf__0461_ 0
C55057 _0417_ _0091_ 0
C55058 _0714_/a_51_297# _0999_/a_1059_315# 0
C55059 _0714_/a_240_47# _0999_/a_27_47# 0
C55060 _0329_ _0728_/a_59_75# 0
C55061 net114 _0738_/a_68_297# 0
C55062 hold75/a_285_47# _0465_ 0.00383f
C55063 _0856_/a_79_21# _0856_/a_215_47# 0.04584f
C55064 _0497_/a_68_297# _0171_ 0
C55065 _0137_ net171 0
C55066 comp0.B\[5\] _0214_ 0
C55067 _0474_ _0563_/a_240_47# 0
C55068 VPWR _0988_/a_561_413# 0.00306f
C55069 VPWR _0553_/a_149_47# 0.00428f
C55070 _1044_/a_27_47# _0542_/a_512_297# 0
C55071 _0327_ _0728_/a_145_75# 0
C55072 _1015_/a_381_47# clknet_1_0__leaf__0457_ 0
C55073 _0504_/a_27_47# _0186_ 0
C55074 _1054_/a_466_413# _0186_ 0
C55075 _0174_ _1043_/a_634_159# 0
C55076 _0786_/a_80_21# _0283_ 0.16732f
C55077 hold75/a_49_47# net58 0.34718f
C55078 net157 _1047_/a_466_413# 0.0239f
C55079 _0216_ _0616_/a_493_297# 0
C55080 pp[30] _0334_ 0
C55081 _0221_ _0219_ 0.25106f
C55082 _0305_ _0767_/a_145_75# 0.0025f
C55083 hold21/a_49_47# output63/a_27_47# 0
C55084 _1016_/a_1059_315# _0181_ 0.02085f
C55085 _0581_/a_373_47# _0242_ 0
C55086 _0236_ _0603_/a_68_297# 0.00143f
C55087 _0233_ _0227_ 0.00978f
C55088 hold45/a_285_47# hold45/a_391_47# 0.41909f
C55089 _1044_/a_891_413# net20 0.0422f
C55090 hold18/a_391_47# _0449_ 0
C55091 _0732_/a_209_297# _0324_ 0.04288f
C55092 _0697_/a_80_21# _0318_ 0.00228f
C55093 _0728_/a_59_75# _0221_ 0.02012f
C55094 _0298_ _0799_/a_303_47# 0
C55095 net66 _0658_/a_113_47# 0
C55096 _0217_ hold71/a_285_47# 0
C55097 _0195_ acc0.A\[27\] 0.10581f
C55098 _0457_ _1015_/a_1059_315# 0.00575f
C55099 _0195_ _0707_/a_544_297# 0
C55100 net184 _0142_ 0
C55101 _0201_ _0172_ 0
C55102 _0329_ _1008_/a_634_159# 0
C55103 net56 _0318_ 0
C55104 acc0.A\[21\] net1 0.00374f
C55105 _0350_ _0378_ 0
C55106 _0276_ _0302_ 0
C55107 _1037_/a_466_413# net29 0
C55108 net82 VPWR 0.45693f
C55109 clknet_0__0458_ _0432_ 0.20778f
C55110 _0234_ _0606_/a_215_297# 0.17624f
C55111 _1001_/a_561_413# VPWR 0.00292f
C55112 net45 _1017_/a_891_413# 0.00599f
C55113 _0551_/a_27_47# acc0.A\[15\] 0
C55114 _0343_ _0393_ 0.13924f
C55115 VPWR _1062_/a_381_47# 0.0758f
C55116 _0616_/a_215_47# _0240_ 0.05427f
C55117 _0780_/a_285_47# _0347_ 0
C55118 _0780_/a_35_297# _0352_ 0
C55119 _0849_/a_79_21# acc0.A\[15\] 0.01969f
C55120 _1021_/a_1059_315# VPWR 0.41569f
C55121 _1039_/a_891_413# _0172_ 0
C55122 _1039_/a_466_413# _0137_ 0.03205f
C55123 _0787_/a_80_21# _0286_ 0
C55124 hold57/a_391_47# clkbuf_1_0__f__0463_/a_110_47# 0
C55125 net172 _1037_/a_193_47# 0
C55126 _1038_/a_193_47# _0135_ 0
C55127 net43 pp[14] 0
C55128 hold58/a_49_47# _0557_/a_51_297# 0
C55129 comp0.B\[13\] _0140_ 0
C55130 _0258_ _0255_ 0.46163f
C55131 _0762_/a_79_21# _0369_ 0.09711f
C55132 acc0.A\[1\] _0580_/a_27_297# 0
C55133 net101 _0118_ 0
C55134 _0279_ _0647_/a_47_47# 0.15521f
C55135 _0343_ _0758_/a_79_21# 0.00149f
C55136 _0998_/a_466_413# _0410_ 0
C55137 _0365_ _0738_/a_68_297# 0.10761f
C55138 _0183_ net106 0
C55139 _0452_ clknet_1_0__leaf__0461_ 0
C55140 comp0.B\[6\] net171 0.06186f
C55141 _0984_/a_634_159# clkbuf_1_0__f__0458_/a_110_47# 0
C55142 _0776_/a_109_297# _0394_ 0
C55143 _0846_/a_240_47# clkbuf_0__0458_/a_110_47# 0
C55144 _0195_ _0364_ 0
C55145 hold10/a_285_47# net36 0.07266f
C55146 output37/a_27_47# A[12] 0.06727f
C55147 hold14/a_49_47# _0175_ 0.01412f
C55148 net53 _0102_ 0
C55149 _1065_/a_634_159# _1065_/a_592_47# 0
C55150 _0677_/a_47_47# _0347_ 0.01798f
C55151 _0183_ _0237_ 0.03074f
C55152 _0217_ _0382_ 0
C55153 _0967_/a_215_297# _1066_/a_27_47# 0.00144f
C55154 _0485_ _1066_/a_634_159# 0
C55155 hold66/a_285_47# _1005_/a_27_47# 0
C55156 hold66/a_49_47# _1005_/a_193_47# 0
C55157 clknet_0__0463_ comp0.B\[15\] 0
C55158 _0198_ _0146_ 0.0184f
C55159 _0520_/a_27_297# net13 0.01725f
C55160 _1036_/a_27_47# B[15] 0
C55161 _1068_/a_193_47# _0487_ 0.00331f
C55162 _0992_/a_27_47# _0811_/a_81_21# 0
C55163 _0216_ _0351_ 0
C55164 _0985_/a_891_413# _0271_ 0
C55165 _0571_/a_27_297# _1027_/a_27_47# 0
C55166 _0658_/a_113_47# _0350_ 0
C55167 net24 comp0.B\[6\] 0.03871f
C55168 _1033_/a_1059_315# net201 0.00467f
C55169 hold79/a_285_47# _1070_/a_381_47# 0
C55170 net226 _1070_/a_27_47# 0
C55171 comp0.B\[12\] _1042_/a_634_159# 0
C55172 comp0.B\[11\] _1042_/a_466_413# 0.02636f
C55173 _0389_ _0609_/a_109_297# 0
C55174 _0266_ net47 0.09615f
C55175 _1014_/a_193_47# _1014_/a_381_47# 0.09503f
C55176 _1014_/a_634_159# _1014_/a_891_413# 0.03684f
C55177 _1014_/a_27_47# _1014_/a_561_413# 0.0027f
C55178 _1071_/a_27_47# _1071_/a_193_47# 0.97386f
C55179 net228 hold82/a_391_47# 0.0681f
C55180 net152 _0202_ 0
C55181 VPWR _1047_/a_975_413# 0.00506f
C55182 _0996_/a_27_47# _0796_/a_79_21# 0.00139f
C55183 net59 _0704_/a_150_297# 0
C55184 _0218_ clkbuf_1_1__f__0459_/a_110_47# 0
C55185 net36 hold60/a_49_47# 0
C55186 _0183_ hold72/a_285_47# 0
C55187 _0130_ _0565_/a_245_297# 0
C55188 _1015_/a_193_47# _0173_ 0
C55189 hold101/a_391_47# net248 0.13057f
C55190 _0985_/a_634_159# _0458_ 0.01206f
C55191 VPWR _0115_ 0.34501f
C55192 _0476_ _1034_/a_27_47# 0
C55193 net45 net223 0
C55194 net30 net174 0.00434f
C55195 _0342_ _0339_ 0.14065f
C55196 _1050_/a_27_47# net9 0.03672f
C55197 net144 VPWR 0.46621f
C55198 _0478_ _0487_ 0.00215f
C55199 clknet_1_1__leaf__0459_ _0410_ 0
C55200 _0183_ _0769_/a_299_297# 0
C55201 _0312_ _0346_ 0.02695f
C55202 _1021_/a_1059_315# net48 0.00284f
C55203 hold87/a_285_47# _0183_ 0
C55204 VPWR _0536_/a_51_297# 0.4802f
C55205 _0541_/a_68_297# hold51/a_285_47# 0.00112f
C55206 VPWR _0796_/a_297_297# 0.01144f
C55207 acc0.A\[8\] A[8] 0
C55208 _1039_/a_466_413# comp0.B\[6\] 0
C55209 _1039_/a_1059_315# comp0.B\[5\] 0
C55210 _0280_ net5 0
C55211 _0717_/a_80_21# _0334_ 0.16097f
C55212 _1055_/a_561_413# net16 0
C55213 _1055_/a_891_413# _0190_ 0
C55214 _0316_ _0330_ 0.13789f
C55215 net185 VPWR 0.38686f
C55216 _0436_ output61/a_27_47# 0.01297f
C55217 clknet_1_1__leaf__0465_ _1060_/a_891_413# 0
C55218 _0344_ _0219_ 0.16865f
C55219 acc0.A\[7\] _0830_/a_79_21# 0
C55220 hold41/a_391_47# net2 0
C55221 net72 _0840_/a_68_297# 0.04611f
C55222 _0179_ _0849_/a_79_21# 0
C55223 _0956_/a_304_297# comp0.B\[0\] 0
C55224 _1000_/a_975_413# net206 0
C55225 _0802_/a_145_75# _0218_ 0.00325f
C55226 _0664_/a_382_297# _0286_ 0
C55227 _0339_ _0334_ 0.10781f
C55228 _0440_ _0085_ 0.26274f
C55229 _1026_/a_466_413# acc0.A\[25\] 0.01582f
C55230 _0276_ net6 0
C55231 _1032_/a_193_47# _0181_ 0.01432f
C55232 _1012_/a_27_47# _0347_ 0.04247f
C55233 _0819_/a_299_297# _0819_/a_384_47# 0
C55234 hold67/a_49_47# net66 0.31263f
C55235 _0149_ _0194_ 0.03982f
C55236 _0330_ _0347_ 0.02301f
C55237 _0470_ clknet_1_1__leaf_clk 0
C55238 hold13/a_49_47# control0.sh 0
C55239 hold21/a_49_47# _0179_ 0
C55240 _0183_ _1059_/a_466_413# 0
C55241 clknet_1_0__leaf__0462_ _0343_ 0
C55242 _1033_/a_193_47# _0564_/a_68_297# 0
C55243 hold47/a_285_47# VPWR 0.28512f
C55244 _0174_ _0175_ 0
C55245 _0311_ _0370_ 0
C55246 _0461_ _0345_ 0.0722f
C55247 _0555_/a_51_297# _0209_ 0
C55248 _0512_/a_27_297# net4 0
C55249 _1013_/a_592_47# _0339_ 0
C55250 hold4/a_49_47# _1023_/a_27_47# 0
C55251 hold46/a_285_47# _0537_/a_68_297# 0
C55252 _0416_ _0647_/a_47_47# 0.00168f
C55253 _0275_ _0991_/a_193_47# 0
C55254 clknet_1_0__leaf__0459_ _1060_/a_634_159# 0
C55255 net103 acc0.A\[17\] 0
C55256 net57 acc0.A\[30\] 0
C55257 _0318_ _0345_ 0
C55258 _1042_/a_27_47# net20 0
C55259 _1050_/a_891_413# net135 0
C55260 _1033_/a_193_47# clknet_1_1__leaf_clk 0
C55261 _0208_ _0526_/a_27_47# 0.06129f
C55262 _0402_ _0654_/a_207_413# 0
C55263 _0481_ _1070_/a_891_413# 0
C55264 _0963_/a_35_297# _0168_ 0
C55265 _0963_/a_285_297# VPWR 0.25621f
C55266 _1037_/a_27_47# _1036_/a_381_47# 0
C55267 _1037_/a_634_159# _1036_/a_1059_315# 0
C55268 _1037_/a_193_47# _1036_/a_891_413# 0
C55269 _1037_/a_466_413# _1036_/a_466_413# 0
C55270 _0955_/a_32_297# _1062_/a_193_47# 0
C55271 output59/a_27_47# pp[30] 0.1618f
C55272 _0518_/a_27_297# net9 0
C55273 _0553_/a_51_297# net29 0.17718f
C55274 _0836_/a_68_297# _0087_ 0.00119f
C55275 _0817_/a_368_297# _0425_ 0.01897f
C55276 _0424_ _0815_/a_199_47# 0
C55277 net203 clknet_0__0463_ 0.02751f
C55278 _0347_ _0242_ 0.01543f
C55279 net144 input4/a_75_212# 0.00562f
C55280 hold67/a_285_47# net76 0
C55281 _0277_ _0668_/a_382_297# 0
C55282 hold55/a_285_47# net1 0
C55283 _0346_ _0417_ 0.10527f
C55284 _0999_/a_381_47# _0352_ 0.01677f
C55285 _0093_ _0997_/a_891_413# 0
C55286 _0983_/a_1059_315# _0294_ 0
C55287 _1013_/a_466_413# pp[31] 0
C55288 _0498_/a_245_297# net247 0.00169f
C55289 _0498_/a_51_297# net7 0.09305f
C55290 net212 _0087_ 0
C55291 A[9] net47 0
C55292 net22 _0546_/a_51_297# 0.11708f
C55293 _0181_ _0721_/a_27_47# 0
C55294 _0625_/a_59_75# VPWR 0.20512f
C55295 _0444_ _0986_/a_27_47# 0
C55296 hold87/a_285_47# acc0.A\[15\] 0
C55297 _0820_/a_510_47# _0428_ 0.00189f
C55298 _0730_/a_510_47# acc0.A\[29\] 0
C55299 comp0.B\[2\] _1033_/a_1059_315# 0
C55300 _1038_/a_1059_315# _0174_ 0
C55301 net150 _1005_/a_466_413# 0.00704f
C55302 acc0.A\[22\] _1005_/a_193_47# 0
C55303 _0183_ _1005_/a_27_47# 0
C55304 net190 _1028_/a_1059_315# 0.0701f
C55305 _0126_ _1028_/a_193_47# 0.27695f
C55306 hold46/a_49_47# VPWR 0.27513f
C55307 _0216_ _1014_/a_891_413# 0
C55308 net158 net10 0.02668f
C55309 net55 clknet_1_1__leaf__0461_ 0
C55310 _0343_ _0714_/a_51_297# 0.00146f
C55311 net16 net142 0.05351f
C55312 hold67/a_49_47# _0350_ 0.04666f
C55313 clknet_1_0__leaf__0458_ _0448_ 0
C55314 _0489_ _0466_ 0
C55315 net43 _0408_ 0.00239f
C55316 net151 _1005_/a_1059_315# 0
C55317 _1003_/a_466_413# clknet_1_0__leaf__0460_ 0.01821f
C55318 net82 clknet_1_0__leaf__0459_ 0.12688f
C55319 _0686_/a_219_297# _0686_/a_301_297# 0.00516f
C55320 net11 _0150_ 0.08037f
C55321 net1 _0165_ 0
C55322 net34 hold89/a_391_47# 0
C55323 _1059_/a_1059_315# net42 0
C55324 _1059_/a_466_413# acc0.A\[15\] 0.00328f
C55325 net3 _0181_ 0.08053f
C55326 _0643_/a_253_297# _0986_/a_193_47# 0
C55327 _0804_/a_79_21# _0281_ 0
C55328 net58 net71 0
C55329 _0663_/a_27_413# _0179_ 0.00936f
C55330 _1018_/a_634_159# _0116_ 0.04134f
C55331 _0315_ acc0.A\[25\] 0
C55332 _1055_/a_27_47# _1055_/a_466_413# 0.27314f
C55333 _1055_/a_193_47# _1055_/a_634_159# 0.12388f
C55334 net31 A[15] 0.00101f
C55335 _1008_/a_466_413# _1008_/a_561_413# 0.00772f
C55336 _1008_/a_634_159# _1008_/a_975_413# 0
C55337 _0119_ clknet_1_1__leaf_clk 0
C55338 _0648_/a_277_297# VPWR 0.00146f
C55339 _0505_/a_27_297# _0505_/a_109_47# 0.00393f
C55340 pp[27] _0338_ 0.04902f
C55341 pp[16] _0995_/a_193_47# 0
C55342 _1020_/a_466_413# _0118_ 0.03059f
C55343 net53 _1025_/a_1059_315# 0.01627f
C55344 _1035_/a_1059_315# _0474_ 0
C55345 _0343_ net206 0
C55346 _1003_/a_27_47# _1003_/a_193_47# 0.96639f
C55347 _0175_ _0208_ 0.84794f
C55348 _1055_/a_27_47# net181 0
C55349 _0229_ _0376_ 0
C55350 VPWR _0614_/a_111_297# 0
C55351 _0679_/a_68_297# _0679_/a_150_297# 0.00477f
C55352 _0430_ _0272_ 0.00192f
C55353 _0371_ clknet_0__0460_ 0.00673f
C55354 net69 _0265_ 0
C55355 clknet_0__0458_ _0986_/a_381_47# 0.00161f
C55356 clknet_0__0457_ _1014_/a_381_47# 0.00304f
C55357 net248 _0369_ 0
C55358 _0176_ _0542_/a_51_297# 0.01322f
C55359 _0627_/a_109_93# _0432_ 0
C55360 _1054_/a_891_413# _0518_/a_27_297# 0
C55361 _1054_/a_1059_315# _0518_/a_109_297# 0
C55362 net84 _1017_/a_634_159# 0
C55363 _0275_ _0423_ 0.00244f
C55364 _1032_/a_1059_315# comp0.B\[0\] 0.08444f
C55365 _1041_/a_975_413# _0172_ 0
C55366 _0997_/a_27_47# _0219_ 0.01661f
C55367 clknet_1_1__leaf__0460_ _0352_ 0.03494f
C55368 _0846_/a_149_47# _0449_ 0.00653f
C55369 _0180_ clkbuf_1_1__f__0457_/a_110_47# 0.00168f
C55370 clkbuf_1_1__f__0457_/a_110_47# net218 0
C55371 clknet_1_1__leaf__0457_ hold71/a_391_47# 0
C55372 hold94/a_285_47# _0219_ 0.03809f
C55373 hold94/a_391_47# net241 0.15575f
C55374 net190 _0347_ 0
C55375 _0991_/a_561_413# acc0.A\[15\] 0
C55376 clknet_0__0459_ net238 0.01554f
C55377 clkbuf_1_0__f__0459_/a_110_47# _0094_ 0
C55378 clknet_1_0__leaf__0462_ _0376_ 0
C55379 _0826_/a_301_297# _0434_ 0
C55380 _0176_ _0142_ 0
C55381 _1038_/a_1059_315# _0208_ 0
C55382 _0734_/a_47_47# _0462_ 0.00144f
C55383 _0734_/a_285_47# clkbuf_0__0462_/a_110_47# 0
C55384 _1054_/a_27_47# _1053_/a_27_47# 0.0045f
C55385 _0465_ _0345_ 0.05553f
C55386 _0221_ hold61/a_49_47# 0
C55387 clknet_1_0__leaf__0459_ _0115_ 0.11942f
C55388 _0559_/a_51_297# _0212_ 0.11546f
C55389 _0982_/a_193_47# _0456_ 0.03286f
C55390 _0982_/a_1059_315# net234 0.00588f
C55391 net161 net24 0.00142f
C55392 _0218_ clknet_1_1__leaf__0465_ 0.00237f
C55393 _0305_ _0401_ 0
C55394 net26 net171 0
C55395 VPWR comp0.B\[14\] 0.81086f
C55396 _0578_/a_373_47# _0183_ 0.00241f
C55397 hold65/a_391_47# clknet_1_0__leaf__0465_ 0
C55398 net187 net150 0
C55399 _0403_ net80 0.09304f
C55400 _0298_ _0668_/a_382_297# 0.01543f
C55401 _0299_ _0668_/a_79_21# 0.19822f
C55402 _0404_ _0668_/a_297_47# 0
C55403 control0.sh net17 0
C55404 acc0.A\[2\] _0345_ 0
C55405 _0745_/a_193_47# _0250_ 0.00394f
C55406 _0464_ net147 0
C55407 _0661_/a_27_297# _0347_ 0
C55408 _0280_ hold81/a_391_47# 0
C55409 _0179_ _1059_/a_466_413# 0
C55410 acc0.A\[3\] _0446_ 0
C55411 hold26/a_391_47# net174 0
C55412 _0180_ input15/a_75_212# 0
C55413 net86 _0347_ 0.06309f
C55414 _1000_/a_1017_47# _0352_ 0.00205f
C55415 hold33/a_391_47# clkbuf_1_0__f__0463_/a_110_47# 0.00133f
C55416 output59/a_27_47# _0339_ 0
C55417 _0367_ _0737_/a_35_297# 0
C55418 hold2/a_49_47# _0465_ 0.01041f
C55419 _0902_/a_27_47# _0460_ 0
C55420 _1016_/a_1059_315# clknet_1_1__leaf__0461_ 0.05688f
C55421 _0459_ net102 0
C55422 _1014_/a_891_413# net247 0
C55423 net24 net26 0.00349f
C55424 _0369_ _0771_/a_215_297# 0
C55425 VPWR _1017_/a_891_413# 0.17297f
C55426 net247 _0492_/a_27_47# 0
C55427 clkbuf_1_0__f__0458_/a_110_47# _0449_ 0
C55428 net87 _0586_/a_27_47# 0.0123f
C55429 _1037_/a_1059_315# comp0.B\[5\] 0.08536f
C55430 acc0.A\[2\] hold2/a_49_47# 0
C55431 _0350_ _0610_/a_59_75# 0
C55432 _0415_ _0802_/a_59_75# 0.11041f
C55433 _0092_ clknet_1_1__leaf__0459_ 0.00302f
C55434 _0116_ _0615_/a_109_297# 0
C55435 _0378_ _1005_/a_1059_315# 0
C55436 VPWR net146 0.53205f
C55437 _0563_/a_51_297# _0563_/a_240_47# 0.03076f
C55438 _0548_/a_51_297# net173 0.07934f
C55439 net105 acc0.A\[19\] 0
C55440 _0506_/a_81_21# _0506_/a_384_47# 0.00138f
C55441 _0695_/a_80_21# _1007_/a_193_47# 0
C55442 VPWR _0543_/a_68_297# 0.16745f
C55443 _0333_ hold95/a_285_47# 0
C55444 pp[28] _0335_ 0.07025f
C55445 _0804_/a_510_47# VPWR 0.00396f
C55446 clkload1/Y _0346_ 0.08206f
C55447 acc0.A\[29\] hold80/a_391_47# 0.01406f
C55448 _1017_/a_466_413# clkbuf_0__0461_/a_110_47# 0.00208f
C55449 _0255_ net72 0
C55450 VPWR _1033_/a_634_159# 0.18459f
C55451 _0724_/a_113_297# _0339_ 0
C55452 clknet_1_1__leaf__0460_ net115 0
C55453 _1044_/a_27_47# _0141_ 0
C55454 _1044_/a_1059_315# net195 0
C55455 clknet_1_0__leaf__0458_ _0217_ 0
C55456 _0243_ _0614_/a_183_297# 0.00358f
C55457 clknet_1_0__leaf__0465_ _1049_/a_634_159# 0.00106f
C55458 _0770_/a_79_21# _0246_ 0
C55459 _0718_/a_47_47# _0334_ 0
C55460 _0251_ _0619_/a_150_297# 0.00193f
C55461 net169 _0186_ 0
C55462 _0174_ net129 0
C55463 _0402_ _0286_ 0.32023f
C55464 VPWR _1050_/a_381_47# 0.07595f
C55465 _0172_ B[12] 0
C55466 _0511_/a_81_21# _0156_ 0.11562f
C55467 _0511_/a_384_47# net192 0.0104f
C55468 net157 _0145_ 0.00576f
C55469 _0579_/a_27_297# clknet_1_0__leaf__0461_ 0
C55470 _0272_ _0443_ 0.10789f
C55471 _1010_/a_634_159# _1010_/a_1059_315# 0
C55472 _1010_/a_27_47# _1010_/a_381_47# 0.06222f
C55473 _1010_/a_193_47# _1010_/a_891_413# 0.19489f
C55474 clknet_1_0__leaf__0462_ _1004_/a_466_413# 0.00483f
C55475 _0717_/a_209_297# _0195_ 0
C55476 net130 _0142_ 0
C55477 net60 output41/a_27_47# 0.00176f
C55478 net54 _1028_/a_193_47# 0
C55479 _0991_/a_466_413# _0181_ 0.01583f
C55480 net125 _0464_ 0
C55481 _1040_/a_193_47# _1040_/a_634_159# 0.11072f
C55482 _1040_/a_27_47# _1040_/a_466_413# 0.26005f
C55483 clknet_1_1__leaf__0458_ _0150_ 0
C55484 _0183_ _0199_ 0
C55485 _0423_ _0657_/a_109_297# 0.00283f
C55486 _0266_ _0848_/a_109_297# 0
C55487 _0305_ _0607_/a_27_297# 0.01908f
C55488 VPWR pp[3] 0.50899f
C55489 _0473_ _0494_/a_27_47# 0.00737f
C55490 acc0.A\[13\] net41 0.09971f
C55491 clknet_1_0__leaf__0457_ acc0.A\[18\] 0.00158f
C55492 _0146_ _1048_/a_466_413# 0.03902f
C55493 _0216_ _0338_ 0
C55494 _0233_ hold30/a_49_47# 0
C55495 _0329_ net94 0.00888f
C55496 net71 _0262_ 0.00569f
C55497 _0452_ _0218_ 0
C55498 _0662_/a_81_21# _0345_ 0.00536f
C55499 _0662_/a_81_21# _0814_/a_27_47# 0.01737f
C55500 _1002_/a_634_159# _0183_ 0.01082f
C55501 _1002_/a_891_413# net150 0.00873f
C55502 _1002_/a_1059_315# _0217_ 0
C55503 _0328_ _0695_/a_80_21# 0.08456f
C55504 _0746_/a_299_297# _0346_ 0.00863f
C55505 _0385_ _0764_/a_81_21# 0.11414f
C55506 _0642_/a_27_413# _0829_/a_27_47# 0
C55507 _0135_ net29 0
C55508 control0.state\[0\] _0949_/a_59_75# 0.08673f
C55509 _0671_/a_199_47# net228 0
C55510 _0369_ _0302_ 0
C55511 VPWR net223 0.271f
C55512 _0248_ _1006_/a_27_47# 0.00626f
C55513 hold54/a_391_47# _0181_ 0
C55514 hold66/a_285_47# _0222_ 0
C55515 _0217_ acc0.A\[16\] 0.09089f
C55516 _0218_ _0567_/a_27_297# 0
C55517 _1020_/a_561_413# _0461_ 0
C55518 _0751_/a_29_53# _0248_ 0
C55519 net74 pp[4] 0.00151f
C55520 _0846_/a_51_297# _0846_/a_512_297# 0.0116f
C55521 output42/a_27_47# _0411_ 0
C55522 net45 _1016_/a_193_47# 0.00241f
C55523 _1067_/a_27_47# _1067_/a_466_413# 0.27314f
C55524 _1067_/a_193_47# _1067_/a_634_159# 0.12497f
C55525 net9 _0987_/a_27_47# 0.03366f
C55526 _1018_/a_1017_47# _0347_ 0
C55527 _0553_/a_51_297# _0137_ 0
C55528 _0136_ _0550_/a_51_297# 0.00136f
C55529 net187 control0.add 0.00512f
C55530 net224 _0108_ 0
C55531 _0178_ _0566_/a_27_47# 0.11533f
C55532 _0369_ _1067_/a_1059_315# 0
C55533 _0210_ _0560_/a_68_297# 0
C55534 _0195_ output60/a_27_47# 0
C55535 acc0.A\[12\] net37 0.57902f
C55536 _0233_ _0352_ 0.355f
C55537 net194 net157 0
C55538 _0399_ net47 0.12062f
C55539 _1072_/a_193_47# _1071_/a_634_159# 0
C55540 _1072_/a_27_47# _1071_/a_466_413# 0
C55541 _0269_ net165 0
C55542 _0575_/a_27_297# _0102_ 0
C55543 VPWR _0740_/a_113_47# 0
C55544 clknet_1_0__leaf__0462_ _0224_ 0.03934f
C55545 net70 clkbuf_1_0__f__0458_/a_110_47# 0.00194f
C55546 _1009_/a_634_159# _1009_/a_381_47# 0
C55547 _0317_ acc0.A\[28\] 0
C55548 _0833_/a_215_47# clknet_1_1__leaf__0465_ 0
C55549 _0989_/a_27_47# _0989_/a_634_159# 0.14145f
C55550 hold1/a_49_47# hold1/a_391_47# 0.00188f
C55551 net69 _0267_ 0
C55552 _0273_ VPWR 0.57001f
C55553 hold65/a_49_47# acc0.A\[8\] 0
C55554 _0800_/a_51_297# _0218_ 0.00243f
C55555 _1065_/a_891_413# control0.reset 0.00905f
C55556 hold5/a_285_47# _0140_ 0.01119f
C55557 hold18/a_49_47# _0448_ 0
C55558 _0313_ _0319_ 0.2638f
C55559 _0982_/a_891_413# VPWR 0.18398f
C55560 clknet_0_clk _1062_/a_1017_47# 0
C55561 _0476_ _1066_/a_1059_315# 0.00106f
C55562 _0280_ _0303_ 0.06044f
C55563 net213 _1005_/a_891_413# 0
C55564 _0992_/a_27_47# _0992_/a_634_159# 0.14145f
C55565 _0817_/a_266_47# _0089_ 0
C55566 _0817_/a_81_21# net67 0
C55567 _1036_/a_561_413# net121 0.00165f
C55568 comp0.B\[4\] _1035_/a_466_413# 0
C55569 clkbuf_1_1__f__0465_/a_110_47# _0186_ 0
C55570 VPWR _1053_/a_193_47# 0.30542f
C55571 _0125_ _1027_/a_27_47# 0.0187f
C55572 acc0.A\[27\] _1027_/a_466_413# 0
C55573 _0199_ acc0.A\[15\] 0.08409f
C55574 _1032_/a_466_413# net118 0
C55575 _0557_/a_149_47# _0211_ 0.00544f
C55576 hold79/a_285_47# control0.count\[1\] 0.00332f
C55577 _1014_/a_193_47# acc0.A\[0\] 0
C55578 _1014_/a_891_413# net100 0
C55579 _1071_/a_466_413# _1071_/a_592_47# 0.00553f
C55580 _1071_/a_634_159# _1071_/a_1017_47# 0
C55581 _0996_/a_193_47# _0094_ 0.26987f
C55582 _0996_/a_466_413# _0410_ 0
C55583 _0996_/a_1059_315# net238 0.06086f
C55584 _1045_/a_27_47# _1043_/a_193_47# 0
C55585 _1045_/a_193_47# _1043_/a_27_47# 0
C55586 _1015_/a_592_47# _0208_ 0
C55587 _1000_/a_27_47# clknet_0__0461_ 0.00494f
C55588 _1000_/a_466_413# clkbuf_1_0__f__0461_/a_110_47# 0.00166f
C55589 hold96/a_49_47# net243 0
C55590 clknet_0__0463_ _0176_ 0.01645f
C55591 net61 _0436_ 0.02763f
C55592 _0343_ _0774_/a_150_297# 0
C55593 net45 _0714_/a_512_297# 0
C55594 net46 _0373_ 0
C55595 _0343_ _0405_ 0.2773f
C55596 _0626_/a_68_297# _0626_/a_150_297# 0.00477f
C55597 _0401_ _0181_ 0.3195f
C55598 _0946_/a_30_53# VPWR 0.18214f
C55599 net64 _0517_/a_81_21# 0
C55600 _0216_ _1026_/a_27_47# 0.00987f
C55601 net155 _1026_/a_193_47# 0
C55602 acc0.A\[11\] net143 0
C55603 net157 _1046_/a_634_159# 0
C55604 _0464_ _0473_ 0
C55605 _0553_/a_51_297# comp0.B\[6\] 0.17687f
C55606 _0350_ hold50/a_285_47# 0
C55607 _0343_ _0356_ 0
C55608 hold79/a_391_47# clkbuf_1_0__f_clk/a_110_47# 0.00974f
C55609 _0216_ _1024_/a_1059_315# 0
C55610 _0487_ clkbuf_1_1__f_clk/a_110_47# 0.00608f
C55611 _0437_ _0989_/a_561_413# 0.00118f
C55612 _0087_ _0989_/a_891_413# 0
C55613 _0216_ net99 0
C55614 _0179_ _0196_ 0.02662f
C55615 net245 net41 0
C55616 net16 _0988_/a_27_47# 0
C55617 net40 pp[14] 0.29779f
C55618 _0650_/a_68_297# net37 0.13685f
C55619 _0181_ net222 0
C55620 _1020_/a_634_159# acc0.A\[20\] 0
C55621 _0330_ _0106_ 0
C55622 clkbuf_1_1__f__0459_/a_110_47# net228 0.00154f
C55623 acc0.A\[29\] _0336_ 0.0025f
C55624 _0243_ _0391_ 0.16237f
C55625 _0787_/a_80_21# net79 0
C55626 _0390_ net223 0.01283f
C55627 _1002_/a_891_413# control0.add 0
C55628 _1042_/a_1059_315# _0542_/a_240_47# 0
C55629 _1042_/a_193_47# _0203_ 0
C55630 _1012_/a_975_413# _0352_ 0
C55631 _0369_ net6 0.01986f
C55632 _0183_ _0157_ 0
C55633 _0530_/a_81_21# hold71/a_285_47# 0
C55634 input10/a_75_212# A[3] 0.19906f
C55635 _0343_ _1016_/a_1017_47# 0
C55636 _1054_/a_27_47# A[5] 0
C55637 _1033_/a_891_413# _0215_ 0.02325f
C55638 _0786_/a_80_21# _0345_ 0.00786f
C55639 _0780_/a_35_297# _0392_ 0
C55640 _0984_/a_634_159# acc0.A\[15\] 0.00465f
C55641 clknet_1_0__leaf__0459_ _1017_/a_891_413# 0.00134f
C55642 _0752_/a_27_413# _0237_ 0.01667f
C55643 hold87/a_49_47# net165 0
C55644 _0183_ _0222_ 0.02066f
C55645 B[2] control0.sh 0
C55646 hold30/a_391_47# _0376_ 0
C55647 _1069_/a_27_47# _1069_/a_1059_315# 0.04672f
C55648 _1069_/a_193_47# _1069_/a_466_413# 0.08301f
C55649 VPWR _1028_/a_27_47# 0.40311f
C55650 net3 _0187_ 0
C55651 net211 clknet_1_0__leaf__0457_ 0.11207f
C55652 _1052_/a_1017_47# _0180_ 0
C55653 _0786_/a_217_297# _0304_ 0
C55654 _0343_ _0773_/a_35_297# 0.00877f
C55655 net230 VPWR 0.15243f
C55656 net120 clknet_1_1__leaf__0463_ 0.23906f
C55657 hold60/a_49_47# hold60/a_391_47# 0.00188f
C55658 net61 acc0.A\[3\] 0.33878f
C55659 clkbuf_0__0465_/a_110_47# _0990_/a_27_47# 0.00126f
C55660 _0735_/a_109_297# _0362_ 0.00158f
C55661 _0954_/a_32_297# _0954_/a_220_297# 0.00132f
C55662 _0179_ _0199_ 0
C55663 _1037_/a_27_47# comp0.B\[4\] 0
C55664 _0225_ _0606_/a_465_297# 0.00163f
C55665 _0191_ net9 0.01264f
C55666 _0998_/a_381_47# _0347_ 0
C55667 input31/a_75_212# input22/a_75_212# 0.01223f
C55668 hold66/a_391_47# _0762_/a_79_21# 0.01558f
C55669 _0361_ _0350_ 0
C55670 hold10/a_285_47# _1039_/a_27_47# 0
C55671 _0182_ _0181_ 0.236f
C55672 _1059_/a_27_47# hold82/a_285_47# 0.00287f
C55673 hold37/a_49_47# VPWR 0.2857f
C55674 _1030_/a_891_413# hold62/a_49_47# 0
C55675 _1030_/a_466_413# hold62/a_391_47# 0
C55676 _0985_/a_1059_315# _0350_ 0
C55677 _0343_ clknet_0__0465_ 0.02485f
C55678 _1018_/a_27_47# clkbuf_1_0__f__0461_/a_110_47# 0
C55679 _0445_ _0986_/a_1017_47# 0
C55680 net243 net90 0
C55681 hold97/a_391_47# _0125_ 0
C55682 _0592_/a_68_297# _0378_ 0.00487f
C55683 net93 net50 0
C55684 _1038_/a_1017_47# _0136_ 0.00192f
C55685 _0577_/a_109_297# _1022_/a_27_47# 0
C55686 _0577_/a_27_297# _1022_/a_193_47# 0
C55687 net45 net41 0.00139f
C55688 _0217_ net91 0
C55689 net150 _0103_ 0.01541f
C55690 _0607_/a_27_297# _0181_ 0.00464f
C55691 _0538_/a_51_297# _0538_/a_512_297# 0.0116f
C55692 _0787_/a_209_297# _0345_ 0
C55693 _0260_ _0846_/a_149_47# 0
C55694 clknet_1_1__leaf__0462_ _1008_/a_381_47# 0
C55695 comp0.B\[6\] _0561_/a_149_47# 0
C55696 _0474_ _0561_/a_245_297# 0.00116f
C55697 comp0.B\[5\] _0561_/a_240_47# 0
C55698 _0481_ clkbuf_1_0__f_clk/a_110_47# 0
C55699 _1032_/a_27_47# net201 0
C55700 _0343_ net225 0.02223f
C55701 net21 hold51/a_285_47# 0
C55702 _0217_ hold18/a_49_47# 0
C55703 VPWR _1046_/a_561_413# 0.00213f
C55704 VPWR _0798_/a_113_297# 0.24689f
C55705 _1022_/a_634_159# _1022_/a_975_413# 0
C55706 _1022_/a_466_413# _1022_/a_561_413# 0.00772f
C55707 _1022_/a_193_47# _1022_/a_592_47# 0.00135f
C55708 comp0.B\[13\] net129 0
C55709 _0231_ _0326_ 0
C55710 hold22/a_391_47# _0518_/a_27_297# 0
C55711 _0313_ _0681_/a_113_47# 0.00961f
C55712 _0101_ clknet_1_0__leaf__0460_ 0.04288f
C55713 net119 clkbuf_1_1__f_clk/a_110_47# 0
C55714 clknet_1_0__leaf__0459_ net223 0
C55715 _1052_/a_381_47# _0525_/a_81_21# 0
C55716 _0157_ acc0.A\[15\] 0.00399f
C55717 _0348_ pp[27] 0.05252f
C55718 _0153_ net2 0
C55719 _0994_/a_27_47# _0994_/a_466_413# 0.27314f
C55720 _0994_/a_193_47# _0994_/a_634_159# 0.12497f
C55721 net105 net1 0.00499f
C55722 _0357_ _0331_ 0
C55723 A[15] net7 0.01221f
C55724 _0285_ _0808_/a_81_21# 0.07524f
C55725 _0275_ _0986_/a_466_413# 0.03043f
C55726 _0779_/a_79_21# _0779_/a_215_47# 0.04584f
C55727 net211 _1001_/a_1059_315# 0
C55728 _0292_ _0812_/a_510_47# 0.00273f
C55729 net104 _0116_ 0.01063f
C55730 _0472_ comp0.B\[5\] 0.00608f
C55731 net44 _0347_ 0.3978f
C55732 _0183_ net220 0
C55733 clknet_1_1__leaf__0459_ _0352_ 0
C55734 clk _0488_ 0.01877f
C55735 _1055_/a_27_47# net179 0.09498f
C55736 _1055_/a_193_47# net141 0.00707f
C55737 _1055_/a_1059_315# _1055_/a_1017_47# 0
C55738 hold88/a_285_47# _0439_ 0
C55739 _0313_ _0733_/a_448_47# 0
C55740 net36 _0263_ 0
C55741 _0718_/a_377_297# _0195_ 0
C55742 hold24/a_391_47# comp0.B\[7\] 0.00107f
C55743 _0305_ _0656_/a_145_75# 0
C55744 hold88/a_285_47# VPWR 0.27304f
C55745 _0984_/a_634_159# _0179_ 0
C55746 VPWR _0758_/a_215_47# 0.00761f
C55747 clkbuf_0__0461_/a_110_47# _0393_ 0.01485f
C55748 hold86/a_391_47# _0452_ 0
C55749 _1003_/a_634_159# _1003_/a_1017_47# 0
C55750 _1003_/a_466_413# _1003_/a_592_47# 0.00553f
C55751 net36 _1047_/a_27_47# 0.0926f
C55752 hold59/a_391_47# net221 0
C55753 _1036_/a_193_47# net27 0
C55754 _0954_/a_32_297# _0540_/a_149_47# 0
C55755 hold45/a_285_47# _1058_/a_193_47# 0
C55756 hold45/a_391_47# _1058_/a_27_47# 0
C55757 _0207_ _1040_/a_634_159# 0.00633f
C55758 _0967_/a_109_93# VPWR 0.13108f
C55759 _0168_ _0484_ 0
C55760 _0466_ net159 0.08348f
C55761 VPWR _0487_ 1.13249f
C55762 clknet_0__0457_ acc0.A\[0\] 0
C55763 clknet_1_0__leaf__0460_ hold4/a_285_47# 0
C55764 net185 comp0.B\[3\] 0.66952f
C55765 hold16/a_391_47# net239 0
C55766 hold20/a_391_47# clknet_0_clk 0.0127f
C55767 hold46/a_285_47# net180 0
C55768 net84 net103 0
C55769 _1054_/a_891_413# _0191_ 0.01713f
C55770 _0217_ _0856_/a_297_297# 0
C55771 _0467_ _0468_ 0.01829f
C55772 _0086_ _0439_ 0
C55773 _0195_ _0097_ 0
C55774 _0216_ _0396_ 0
C55775 _0844_/a_79_21# _0447_ 0.16653f
C55776 _1004_/a_891_413# _0352_ 0
C55777 VPWR _0086_ 0.29652f
C55778 net190 _0106_ 0
C55779 _0410_ _0095_ 0
C55780 _0983_/a_634_159# _0347_ 0.0019f
C55781 hold56/a_49_47# comp0.B\[2\] 0.30063f
C55782 _0603_/a_150_297# _0765_/a_79_21# 0
C55783 net23 _1065_/a_466_413# 0.02301f
C55784 _0330_ _1011_/a_27_47# 0
C55785 _1054_/a_381_47# _1053_/a_891_413# 0
C55786 _0765_/a_215_47# hold73/a_285_47# 0.00236f
C55787 _0799_/a_80_21# _0411_ 0.19186f
C55788 _1012_/a_1059_315# _0350_ 0.00778f
C55789 _0195_ _0580_/a_109_47# 0
C55790 _0216_ _0580_/a_27_297# 0
C55791 _0284_ _0404_ 0
C55792 _0664_/a_297_47# _0345_ 0.00426f
C55793 _0226_ VPWR 0.94704f
C55794 VPWR _0987_/a_381_47# 0.07795f
C55795 _1024_/a_634_159# _1024_/a_466_413# 0.23992f
C55796 _1024_/a_193_47# _1024_/a_1059_315# 0.03405f
C55797 _1024_/a_27_47# _1024_/a_891_413# 0.03224f
C55798 _0217_ _0247_ 0.09158f
C55799 hold93/a_285_47# hold93/a_391_47# 0.41909f
C55800 _0557_/a_240_47# net160 0.04547f
C55801 hold58/a_391_47# _0211_ 0
C55802 _0816_/a_68_297# _0290_ 0
C55803 hold41/a_49_47# net67 0
C55804 clkbuf_1_0__f__0457_/a_110_47# _0217_ 0.04156f
C55805 _0337_ _0707_/a_75_199# 0
C55806 _0293_ _0347_ 0
C55807 B[9] _1042_/a_27_47# 0.00311f
C55808 comp0.B\[0\] _0468_ 0
C55809 _1011_/a_193_47# _0333_ 0.003f
C55810 VPWR _0727_/a_193_47# 0
C55811 _0179_ _0157_ 0.08057f
C55812 _0985_/a_27_47# _0180_ 0
C55813 _0985_/a_193_47# _0182_ 0
C55814 _0458_ _0636_/a_145_75# 0
C55815 _1007_/a_27_47# net52 0
C55816 _0285_ _0296_ 0.00913f
C55817 _1000_/a_1059_315# _0388_ 0
C55818 _1000_/a_891_413# _0386_ 0.01242f
C55819 VPWR _1029_/a_381_47# 0.07897f
C55820 _0433_ clkbuf_1_1__f__0458_/a_110_47# 0.00168f
C55821 _0387_ _0397_ 0.0098f
C55822 net80 acc0.A\[13\] 0
C55823 comp0.B\[2\] _1032_/a_27_47# 0
C55824 _0343_ _0591_/a_109_297# 0.00376f
C55825 _0540_/a_51_297# _0540_/a_240_47# 0.03076f
C55826 _0982_/a_891_413# _0453_ 0
C55827 clk _1064_/a_27_47# 0.01094f
C55828 net48 _0487_ 0
C55829 clkbuf_1_1__f__0460_/a_110_47# _1010_/a_634_159# 0
C55830 _1048_/a_1059_315# _1048_/a_891_413# 0.31086f
C55831 _1048_/a_193_47# _1048_/a_975_413# 0
C55832 _1048_/a_466_413# _1048_/a_381_47# 0.03733f
C55833 net36 clknet_1_0__leaf__0461_ 0.0128f
C55834 _0481_ control0.count\[2\] 0
C55835 _1034_/a_466_413# clknet_1_1__leaf__0463_ 0.00627f
C55836 _0343_ _0387_ 0
C55837 net63 _0522_/a_27_297# 0
C55838 _0399_ _0796_/a_510_47# 0.00386f
C55839 _0086_ output62/a_27_47# 0
C55840 clknet_0__0461_ acc0.A\[19\] 0
C55841 hold48/a_49_47# clknet_1_1__leaf__0464_ 0.00134f
C55842 _0135_ comp0.B\[6\] 0
C55843 VPWR _1016_/a_193_47# 0.28074f
C55844 net108 VPWR 0.47562f
C55845 clknet_1_1__leaf__0465_ net228 0
C55846 _0223_ _0368_ 0
C55847 _0846_/a_240_47# _0447_ 0.00166f
C55848 _0846_/a_245_297# _0448_ 0
C55849 _0556_/a_150_297# _0211_ 0
C55850 _0251_ _0434_ 0.18742f
C55851 _0804_/a_79_21# _0803_/a_68_297# 0
C55852 VPWR net119 0.69062f
C55853 net23 clknet_1_0__leaf__0460_ 0.04107f
C55854 net124 comp0.B\[8\] 0
C55855 _0427_ _0818_/a_193_47# 0.01319f
C55856 clknet_1_0__leaf__0465_ net135 0.00655f
C55857 _0190_ net47 0
C55858 _0600_/a_103_199# _0249_ 0.00932f
C55859 _0223_ _0618_/a_215_47# 0.05376f
C55860 _0670_/a_79_21# acc0.A\[15\] 0.10578f
C55861 _0670_/a_297_297# net42 0
C55862 _0399_ _0294_ 0.0231f
C55863 _0398_ _0218_ 0.40199f
C55864 net55 _0354_ 0
C55865 _0810_/a_113_47# _0421_ 0.00937f
C55866 VPWR acc0.A\[4\] 1.29698f
C55867 _0226_ net48 0.34814f
C55868 _0217_ _0455_ 0
C55869 net152 _0544_/a_149_47# 0.03548f
C55870 _0546_/a_512_297# net18 0
C55871 _0981_/a_109_297# _0974_/a_79_199# 0
C55872 _0981_/a_27_297# _0974_/a_222_93# 0
C55873 acc0.A\[21\] _0462_ 0
C55874 _0729_/a_68_297# _0729_/a_150_297# 0.00477f
C55875 pp[30] hold15/a_285_47# 0.01308f
C55876 _0348_ _0216_ 0
C55877 VPWR clkbuf_0__0457_/a_110_47# 1.22661f
C55878 _1056_/a_27_47# net2 0
C55879 _0130_ _1015_/a_1059_315# 0.01116f
C55880 net165 _0082_ 0
C55881 _0089_ _0181_ 0.41762f
C55882 _0366_ net90 0
C55883 _0797_/a_27_413# _0797_/a_207_413# 0.18542f
C55884 _1040_/a_1059_315# _1040_/a_1017_47# 0
C55885 _1040_/a_27_47# net174 0.08739f
C55886 _0302_ _0409_ 0
C55887 _0195_ _0689_/a_68_297# 0
C55888 clknet_1_0__leaf__0465_ _1054_/a_27_47# 0
C55889 hold28/a_49_47# net71 0.00212f
C55890 _0795_/a_299_297# _0409_ 0.06696f
C55891 clknet_1_1__leaf__0460_ _0392_ 0
C55892 _0979_/a_109_47# _0480_ 0.00219f
C55893 _0979_/a_109_297# net164 0.01201f
C55894 _1017_/a_634_159# acc0.A\[18\] 0
C55895 _0329_ _0328_ 0
C55896 _0853_/a_68_297# _0853_/a_150_297# 0.00477f
C55897 _0642_/a_215_297# _0827_/a_27_47# 0
C55898 _0527_/a_27_297# net11 0.17462f
C55899 _1072_/a_634_159# _1072_/a_466_413# 0.23992f
C55900 _1072_/a_193_47# _1072_/a_1059_315# 0.03405f
C55901 _1072_/a_27_47# _1072_/a_891_413# 0.03089f
C55902 net58 _0434_ 0
C55903 _0216_ _1027_/a_975_413# 0
C55904 _0830_/a_79_21# _0186_ 0.10022f
C55905 control0.reset _0214_ 0.03791f
C55906 _0841_/a_297_297# _0841_/a_215_47# 0
C55907 _0841_/a_79_21# _0841_/a_510_47# 0.00844f
C55908 net9 input11/a_75_212# 0
C55909 net88 _0183_ 0
C55910 _0328_ clknet_1_0__leaf__0460_ 0
C55911 net35 clknet_1_0__leaf__0460_ 0.03112f
C55912 VPWR _1019_/a_561_413# 0.00213f
C55913 _0714_/a_512_297# VPWR 0.00609f
C55914 B[11] net10 0.01975f
C55915 _0313_ _0732_/a_80_21# 0.12425f
C55916 _0532_/a_384_47# clknet_1_1__leaf__0457_ 0
C55917 VPWR _0694_/a_113_47# 0
C55918 _0119_ _0902_/a_27_47# 0
C55919 net1 _0381_ 0
C55920 net108 net48 0.00428f
C55921 acc0.A\[14\] _0996_/a_592_47# 0
C55922 _0218_ _0277_ 0.05976f
C55923 _1067_/a_1059_315# _1067_/a_1017_47# 0
C55924 clknet_1_0__leaf__0460_ _0599_/a_113_47# 0
C55925 _0244_ _1018_/a_466_413# 0
C55926 net44 hold95/a_49_47# 0
C55927 _0251_ acc0.A\[7\] 0.23838f
C55928 _0251_ _0989_/a_1059_315# 0.08483f
C55929 _0429_ _0989_/a_634_159# 0
C55930 _1001_/a_561_413# _0345_ 0.00157f
C55931 comp0.B\[4\] _0561_/a_51_297# 0.01146f
C55932 _1002_/a_1059_315# _0235_ 0
C55933 _0179_ acc0.A\[9\] 0.02796f
C55934 _0342_ _0999_/a_193_47# 0
C55935 _0346_ _0992_/a_1017_47# 0
C55936 _0462_ _0245_ 0.00166f
C55937 _1071_/a_891_413# _0169_ 0
C55938 _1050_/a_891_413# _0172_ 0
C55939 net45 _0773_/a_285_297# 0
C55940 hold90/a_285_47# _0219_ 0.01067f
C55941 _0449_ acc0.A\[15\] 0.00138f
C55942 _1004_/a_193_47# _0350_ 0.01497f
C55943 _1004_/a_27_47# _0380_ 0
C55944 _0216_ _0332_ 0
C55945 control0.state\[1\] _1002_/a_891_413# 0
C55946 net65 _0989_/a_1017_47# 0.00202f
C55947 _0989_/a_891_413# _0989_/a_975_413# 0.00851f
C55948 _0989_/a_381_47# _0989_/a_561_413# 0.00123f
C55949 VPWR _0807_/a_68_297# 0.15658f
C55950 _0997_/a_634_159# _0997_/a_466_413# 0.23992f
C55951 _0997_/a_193_47# _0997_/a_1059_315# 0.03405f
C55952 _0997_/a_27_47# _0997_/a_891_413# 0.03089f
C55953 _0181_ _0986_/a_891_413# 0.00262f
C55954 _0248_ _0247_ 0.00122f
C55955 net162 _0195_ 0.5222f
C55956 net36 net133 0.07439f
C55957 acc0.A\[31\] _0216_ 0
C55958 acc0.A\[16\] _0583_/a_373_47# 0.00266f
C55959 net194 net13 0.0016f
C55960 _0992_/a_891_413# _0992_/a_975_413# 0.00851f
C55961 _0992_/a_381_47# _0992_/a_561_413# 0.00123f
C55962 _0313_ _0250_ 0
C55963 VPWR _1051_/a_466_413# 0.24987f
C55964 comp0.B\[4\] _0133_ 0.02024f
C55965 _0323_ clkbuf_1_0__f__0462_/a_110_47# 0
C55966 net78 hold81/a_285_47# 0
C55967 clkbuf_1_0__f__0457_/a_110_47# _0248_ 0.00119f
C55968 _0159_ _0138_ 0
C55969 _0570_/a_109_47# acc0.A\[25\] 0
C55970 _0402_ _0808_/a_585_47# 0
C55971 hold6/a_285_47# _1042_/a_27_47# 0
C55972 hold6/a_49_47# _1042_/a_193_47# 0
C55973 VPWR _1045_/a_891_413# 0.19135f
C55974 _0402_ net79 0.00145f
C55975 acc0.A\[27\] net156 0
C55976 clknet_0__0458_ _0841_/a_215_47# 0.00246f
C55977 net202 net118 0.03826f
C55978 _0109_ _1029_/a_1059_315# 0
C55979 _0355_ _1029_/a_975_413# 0
C55980 _0354_ _1029_/a_592_47# 0
C55981 _0218_ _0808_/a_81_21# 0
C55982 control0.reset _1061_/a_1059_315# 0
C55983 hold13/a_391_47# comp0.B\[6\] 0.02069f
C55984 _0376_ _0591_/a_109_297# 0
C55985 clknet_1_1__leaf__0464_ net12 0.00572f
C55986 _0793_/a_51_297# _0405_ 0.00128f
C55987 clknet_1_1__leaf__0463_ net118 0.10398f
C55988 _0710_/a_109_297# clknet_1_1__leaf__0461_ 0
C55989 _1027_/a_27_47# _1027_/a_634_159# 0.14145f
C55990 _0743_/a_51_297# _0105_ 0.11103f
C55991 net45 _0350_ 0
C55992 _0558_/a_68_297# comp0.B\[4\] 0.00114f
C55993 output65/a_27_47# hold65/a_391_47# 0
C55994 hold46/a_285_47# hold26/a_285_47# 0.0073f
C55995 _0285_ _0811_/a_81_21# 0
C55996 net10 _0544_/a_512_297# 0
C55997 net45 _0111_ 0.05102f
C55998 hold54/a_285_47# net201 0.00974f
C55999 _1061_/a_193_47# _1061_/a_975_413# 0
C56000 _1061_/a_466_413# _1061_/a_381_47# 0.03733f
C56001 _1061_/a_1059_315# _1061_/a_891_413# 0.31086f
C56002 net51 _0754_/a_149_47# 0.00109f
C56003 net36 _0585_/a_27_297# 0
C56004 output64/a_27_47# clknet_1_1__leaf__0465_ 0
C56005 net66 _0990_/a_1059_315# 0.10827f
C56006 acc0.A\[8\] _0990_/a_466_413# 0.01652f
C56007 _0291_ _0990_/a_634_159# 0
C56008 _0257_ _0258_ 0.0166f
C56009 _0195_ net112 0
C56010 net157 net132 0
C56011 _0984_/a_193_47# net165 0
C56012 _0361_ _0731_/a_299_297# 0
C56013 _0319_ _0321_ 0.18651f
C56014 _0409_ net6 0.49047f
C56015 _1035_/a_27_47# _1035_/a_1059_315# 0.04875f
C56016 _1035_/a_193_47# _1035_/a_466_413# 0.07543f
C56017 _0399_ _0833_/a_297_297# 0.00472f
C56018 _0424_ _0288_ 0
C56019 _0734_/a_377_297# _0219_ 0
C56020 VPWR net41 3.16813f
C56021 output37/a_27_47# _0511_/a_81_21# 0
C56022 _0959_/a_217_297# _1065_/a_193_47# 0
C56023 _0959_/a_472_297# _1065_/a_27_47# 0
C56024 net156 _0364_ 0.01043f
C56025 _0956_/a_32_297# _0215_ 0.00151f
C56026 _0415_ _0414_ 0.00639f
C56027 hold75/a_49_47# acc0.A\[14\] 0
C56028 _0217_ _1014_/a_592_47# 0
C56029 _0551_/a_27_47# _0171_ 0.1634f
C56030 _0787_/a_303_47# _0091_ 0
C56031 _0489_ _1069_/a_1059_315# 0.02632f
C56032 clknet_1_0__leaf__0462_ clkbuf_0__0462_/a_110_47# 0
C56033 net36 comp0.B\[10\] 0
C56034 _0180_ _0197_ 0.37673f
C56035 _0661_/a_27_297# _0425_ 0
C56036 _1013_/a_27_47# clknet_1_1__leaf__0461_ 0.00147f
C56037 hold89/a_391_47# _0166_ 0
C56038 _0179_ _0449_ 0.00761f
C56039 net169 input12/a_75_212# 0
C56040 net70 acc0.A\[15\] 0.00479f
C56041 hold11/a_49_47# net134 0.00301f
C56042 net76 _0990_/a_891_413# 0
C56043 _0298_ _0218_ 0.02162f
C56044 _0607_/a_27_297# clknet_1_1__leaf__0461_ 0
C56045 hold20/a_49_47# _0466_ 0
C56046 hold20/a_285_47# _0488_ 0
C56047 acc0.A\[29\] _1029_/a_27_47# 0.00312f
C56048 _0268_ _0636_/a_59_75# 0.11002f
C56049 clknet_1_0__leaf__0459_ _1016_/a_193_47# 0.02522f
C56050 _1069_/a_634_159# clknet_1_0__leaf_clk 0
C56051 _1069_/a_891_413# _1069_/a_1017_47# 0.00617f
C56052 _1069_/a_193_47# _0167_ 0.26143f
C56053 _1056_/a_1059_315# net66 0.01134f
C56054 VPWR net217 0.22183f
C56055 _0854_/a_215_47# _0181_ 0.04859f
C56056 _0384_ hold73/a_49_47# 0
C56057 _0186_ _0219_ 0
C56058 _1059_/a_634_159# _0185_ 0.00106f
C56059 VPWR _0534_/a_299_297# 0.20951f
C56060 _0662_/a_384_47# _0346_ 0
C56061 comp0.B\[11\] comp0.B\[12\] 0.05869f
C56062 pp[8] _1055_/a_634_159# 0
C56063 VPWR A[11] 0.84894f
C56064 _0555_/a_240_47# net29 0
C56065 _0233_ _0600_/a_253_297# 0.00207f
C56066 _0343_ _0600_/a_253_47# 0.00587f
C56067 _0231_ _0600_/a_103_199# 0.12267f
C56068 VPWR hold62/a_285_47# 0.2871f
C56069 _0296_ _0218_ 0
C56070 _0111_ _0587_/a_27_47# 0
C56071 comp0.B\[6\] _0160_ 0.00352f
C56072 _1041_/a_1059_315# _1040_/a_891_413# 0
C56073 _1041_/a_466_413# _1040_/a_381_47# 0.00131f
C56074 _1015_/a_27_47# _0721_/a_27_47# 0.0105f
C56075 _1031_/a_592_47# _0220_ 0.00269f
C56076 _0997_/a_1059_315# _0411_ 0
C56077 net213 _0369_ 0.40477f
C56078 acc0.A\[27\] acc0.A\[26\] 0
C56079 clknet_1_1__leaf__0462_ net113 0.13126f
C56080 _0990_/a_1059_315# _0350_ 0
C56081 _0577_/a_27_297# _0577_/a_373_47# 0.01338f
C56082 hold19/a_49_47# _0219_ 0
C56083 _1027_/a_193_47# _1026_/a_1059_315# 0
C56084 _1027_/a_27_47# _1026_/a_891_413# 0
C56085 _0533_/a_27_297# _0171_ 0.0034f
C56086 hold26/a_391_47# comp0.B\[14\] 0
C56087 _0176_ net198 0
C56088 _0349_ pp[28] 0.11897f
C56089 _0137_ _0206_ 0
C56090 _1002_/a_592_47# _0181_ 0
C56091 _0959_/a_217_297# net33 0.01717f
C56092 clknet_1_0__leaf__0459_ clkbuf_0__0457_/a_110_47# 0.01784f
C56093 hold96/a_49_47# acc0.A\[24\] 0
C56094 _0343_ _1011_/a_891_413# 0
C56095 _0305_ _0679_/a_68_297# 0.00409f
C56096 _0680_/a_217_297# _0310_ 0
C56097 net237 clkbuf_1_0__f__0462_/a_110_47# 0.00671f
C56098 _0120_ _1022_/a_193_47# 0.00384f
C56099 _0217_ _1022_/a_891_413# 0
C56100 acc0.A\[22\] _1022_/a_1059_315# 0.17536f
C56101 _0816_/a_68_297# net77 0
C56102 _0228_ net51 0
C56103 _0343_ _1006_/a_27_47# 0
C56104 clknet_1_1__leaf__0458_ _0989_/a_634_159# 0
C56105 hold57/a_391_47# net160 0
C56106 hold57/a_285_47# _0210_ 0.00443f
C56107 hold1/a_391_47# clknet_1_1__leaf__0458_ 0.0246f
C56108 VPWR _0744_/a_27_47# 0.52744f
C56109 _0561_/a_240_47# hold84/a_49_47# 0
C56110 _0538_/a_51_297# _0143_ 0.10219f
C56111 _0538_/a_240_47# net183 0.08235f
C56112 _0538_/a_149_47# net21 0.00184f
C56113 _0227_ _0754_/a_51_297# 0.00101f
C56114 _0343_ _0751_/a_29_53# 0
C56115 VPWR _0760_/a_47_47# 0.37315f
C56116 clknet_1_0__leaf__0463_ _0498_/a_512_297# 0
C56117 _0135_ net26 0.00277f
C56118 _1022_/a_561_413# net151 0
C56119 hold54/a_285_47# comp0.B\[2\] 0
C56120 output53/a_27_47# _0195_ 0
C56121 pp[25] _0572_/a_109_47# 0
C56122 hold22/a_391_47# _0191_ 0.03733f
C56123 net64 _0990_/a_466_413# 0
C56124 _0343_ _0986_/a_27_47# 0
C56125 _1018_/a_381_47# _0264_ 0
C56126 clknet_0__0462_ _0219_ 0.12673f
C56127 _0325_ _0693_/a_68_297# 0.12172f
C56128 hold64/a_285_47# _0580_/a_27_297# 0
C56129 net43 net83 0.03951f
C56130 net199 _1025_/a_561_413# 0
C56131 _0994_/a_1059_315# _0994_/a_1017_47# 0
C56132 _1020_/a_1017_47# clknet_1_0__leaf__0457_ 0
C56133 acc0.A\[26\] _0364_ 0.05188f
C56134 _0284_ _0419_ 0.0274f
C56135 _0579_/a_27_297# _0099_ 0
C56136 hold74/a_285_47# _0195_ 0
C56137 _1056_/a_1059_315# _0350_ 0
C56138 clkbuf_1_1__f__0461_/a_110_47# clknet_0__0461_ 0.31019f
C56139 _0500_/a_27_47# _1048_/a_634_159# 0
C56140 _0733_/a_222_93# acc0.A\[27\] 0
C56141 _0972_/a_93_21# _0972_/a_256_47# 0.01135f
C56142 hold56/a_285_47# _0215_ 0.00383f
C56143 _1023_/a_561_413# net51 0
C56144 _0401_ _0990_/a_193_47# 0
C56145 _0720_/a_150_297# clknet_1_1__leaf__0462_ 0.00194f
C56146 _0835_/a_215_47# _0271_ 0.00157f
C56147 net70 _0179_ 0.34018f
C56148 _0346_ _0261_ 0
C56149 _0781_/a_68_297# net43 0.1387f
C56150 _0752_/a_27_413# _0222_ 0.04563f
C56151 hold14/a_49_47# comp0.B\[4\] 0.01374f
C56152 _1003_/a_592_47# _0101_ 0.00164f
C56153 comp0.B\[12\] _0202_ 0.29384f
C56154 _0993_/a_634_159# _0993_/a_466_413# 0.23992f
C56155 _0993_/a_193_47# _0993_/a_1059_315# 0.03405f
C56156 _0993_/a_27_47# _0993_/a_891_413# 0.03224f
C56157 _0816_/a_68_297# _0656_/a_59_75# 0.0083f
C56158 A[11] input4/a_75_212# 0.03221f
C56159 input3/a_75_212# A[12] 0.00154f
C56160 _1058_/a_634_159# _0156_ 0
C56161 net171 net174 0
C56162 hold45/a_49_47# net144 0.01098f
C56163 _1039_/a_1059_315# _1039_/a_891_413# 0.31086f
C56164 _1039_/a_193_47# _1039_/a_975_413# 0
C56165 _1039_/a_466_413# _1039_/a_381_47# 0.03733f
C56166 _0182_ _0531_/a_27_297# 0.12739f
C56167 hold33/a_285_47# _0138_ 0.06131f
C56168 _0578_/a_109_47# net1 0
C56169 _0280_ _0672_/a_215_47# 0.06011f
C56170 _0663_/a_27_413# _0292_ 0.00151f
C56171 _0532_/a_299_297# _0530_/a_81_21# 0
C56172 A[12] _0512_/a_373_47# 0
C56173 _1056_/a_466_413# net64 0
C56174 _0996_/a_27_47# _0400_ 0
C56175 _0172_ _1046_/a_381_47# 0.00609f
C56176 _1032_/a_193_47# _0215_ 0
C56177 _1049_/a_634_159# _0148_ 0
C56178 _1049_/a_891_413# _0196_ 0
C56179 B[3] B[4] 0.11159f
C56180 _0311_ _0240_ 0.00259f
C56181 net33 _1062_/a_592_47# 0
C56182 _1026_/a_634_159# _1026_/a_381_47# 0
C56183 hold74/a_49_47# _0369_ 0
C56184 _0733_/a_448_47# _0321_ 0.06018f
C56185 _0985_/a_381_47# clknet_1_0__leaf__0458_ 0
C56186 net69 _0347_ 0.12963f
C56187 _0311_ _0369_ 0.11198f
C56188 net36 _0848_/a_27_47# 0
C56189 _0343_ _0340_ 0.21948f
C56190 net140 _1053_/a_592_47# 0.00112f
C56191 net169 _1053_/a_975_413# 0
C56192 _0629_/a_59_75# _0261_ 0.17398f
C56193 _0216_ _0117_ 0
C56194 _0118_ _1001_/a_27_47# 0
C56195 net36 _0218_ 0.09353f
C56196 net90 acc0.A\[24\] 0.00149f
C56197 _0762_/a_79_21# _0374_ 0
C56198 _1024_/a_634_159# _0122_ 0.00401f
C56199 _1024_/a_466_413# net110 0
C56200 _0854_/a_79_21# _1018_/a_634_159# 0
C56201 _0854_/a_215_47# _1018_/a_27_47# 0
C56202 _0183_ _1067_/a_891_413# 0
C56203 _0343_ clknet_1_0__leaf__0458_ 0.00424f
C56204 _0502_/a_27_47# _0178_ 0
C56205 _0246_ acc0.A\[18\] 0
C56206 _0337_ _0338_ 0.17193f
C56207 _1014_/a_466_413# _0181_ 0
C56208 clknet_1_1__leaf__0464_ _0203_ 0
C56209 _0278_ _0646_/a_377_297# 0.00188f
C56210 _0234_ _0223_ 0
C56211 _1036_/a_1059_315# net25 0
C56212 _0439_ net66 0
C56213 _1057_/a_193_47# net143 0.016f
C56214 _0471_ _1063_/a_27_47# 0
C56215 _0090_ clknet_1_1__leaf__0465_ 0.00586f
C56216 net45 _0244_ 0.60649f
C56217 pp[16] _0997_/a_27_47# 0
C56218 clknet_1_0__leaf__0459_ net41 0
C56219 VPWR net66 1.29372f
C56220 _0199_ _1049_/a_891_413# 0
C56221 VPWR input21/a_75_212# 0.26087f
C56222 _0540_/a_512_297# _0142_ 0
C56223 _0269_ acc0.A\[3\] 0
C56224 net243 _0183_ 0
C56225 clkbuf_1_1__f__0460_/a_110_47# net96 0.00219f
C56226 net189 input2/a_75_212# 0
C56227 net168 acc0.A\[7\] 0.11747f
C56228 hold78/a_391_47# _0220_ 0
C56229 _0356_ _0568_/a_27_297# 0
C56230 _0831_/a_285_297# _0434_ 0.05826f
C56231 _0988_/a_27_47# net142 0
C56232 B[13] _1043_/a_1059_315# 0
C56233 net63 _0193_ 0
C56234 _1068_/a_381_47# _0468_ 0.01602f
C56235 net1 _0468_ 0.40067f
C56236 _1041_/a_27_47# _1041_/a_1059_315# 0.04721f
C56237 _1041_/a_193_47# _1041_/a_466_413# 0.07834f
C56238 _1048_/a_27_47# clknet_1_1__leaf__0457_ 0
C56239 _0624_/a_59_75# _0256_ 0.13373f
C56240 _0624_/a_145_75# _0270_ 0
C56241 net121 input24/a_75_212# 0
C56242 net3 clknet_1_1__leaf__0465_ 0.07809f
C56243 VPWR _0991_/a_27_47# 0.69815f
C56244 hold99/a_391_47# _0993_/a_27_47# 0
C56245 hold99/a_285_47# _0993_/a_193_47# 0
C56246 _0490_ clkbuf_0_clk/a_110_47# 0
C56247 _0232_ clkbuf_1_0__f__0460_/a_110_47# 0.00304f
C56248 _1017_/a_193_47# _0219_ 0
C56249 _0172_ _0271_ 0
C56250 _0343_ acc0.A\[16\] 0.07772f
C56251 VPWR _0773_/a_285_297# 0.26387f
C56252 hold69/a_391_47# _0352_ 0.00141f
C56253 _0341_ net60 0.80914f
C56254 _1015_/a_891_413# comp0.B\[15\] 0.0034f
C56255 _0172_ _0987_/a_891_413# 0
C56256 _0260_ acc0.A\[15\] 0
C56257 _1002_/a_193_47# net1 0.01644f
C56258 _0232_ _0250_ 0
C56259 _0415_ _0404_ 0.05549f
C56260 _0369_ hold73/a_391_47# 0.00726f
C56261 _0346_ net47 0.35937f
C56262 _0274_ _0825_/a_68_297# 0.00565f
C56263 clknet_0__0457_ hold73/a_391_47# 0
C56264 _0139_ net18 0
C56265 net32 _0140_ 0.0235f
C56266 _0569_/a_27_297# net114 0.00152f
C56267 _0170_ _0974_/a_222_93# 0
C56268 _0216_ _0368_ 0.00744f
C56269 hold2/a_391_47# net149 0.1316f
C56270 clknet_0__0464_ _1061_/a_466_413# 0
C56271 clkbuf_1_1__f__0460_/a_110_47# _0315_ 0
C56272 net163 _0220_ 0.03278f
C56273 _0707_/a_75_199# _0333_ 0.19168f
C56274 clknet_0__0460_ _1006_/a_1059_315# 0
C56275 _0305_ _0608_/a_27_47# 0
C56276 _0191_ _0255_ 0
C56277 _0644_/a_47_47# clkbuf_1_1__f__0459_/a_110_47# 0.00557f
C56278 hold44/a_285_47# _1029_/a_634_159# 0.01163f
C56279 hold44/a_391_47# _1029_/a_193_47# 0.00283f
C56280 _0439_ _0350_ 0.10887f
C56281 clknet_0__0458_ _0627_/a_297_297# 0
C56282 net103 acc0.A\[18\] 0
C56283 hold85/a_285_47# hold84/a_391_47# 0
C56284 hold85/a_391_47# hold84/a_285_47# 0
C56285 net217 _0283_ 0
C56286 net101 _0178_ 0
C56287 comp0.B\[3\] _0487_ 0
C56288 _0461_ clknet_1_0__leaf__0457_ 0.09779f
C56289 VPWR _0350_ 5.29253f
C56290 net201 _0562_/a_68_297# 0.18466f
C56291 _0111_ VPWR 0.2857f
C56292 _0285_ _0652_/a_109_297# 0
C56293 _0414_ _0347_ 0
C56294 clknet_1_0__leaf__0461_ hold60/a_391_47# 0.02839f
C56295 _0252_ _0831_/a_35_297# 0
C56296 net65 _0831_/a_285_47# 0
C56297 _0554_/a_150_297# _0210_ 0
C56298 hold68/a_285_47# _0352_ 0
C56299 _1013_/a_891_413# net60 0.00708f
C56300 VPWR _1025_/a_561_413# 0.00292f
C56301 _0293_ _0991_/a_1059_315# 0
C56302 _1055_/a_1059_315# _0186_ 0
C56303 _0258_ clknet_1_1__leaf__0458_ 0.04393f
C56304 _0257_ net72 0
C56305 net223 _0345_ 0.00223f
C56306 clknet_1_1__leaf__0462_ hold92/a_391_47# 0.00849f
C56307 net26 _0160_ 0
C56308 VPWR _0463_ 0.63865f
C56309 comp0.B\[4\] _0208_ 0.29934f
C56310 _0743_/a_51_297# _0359_ 0.1199f
C56311 _0625_/a_59_75# _0836_/a_68_297# 0.0083f
C56312 net21 clkbuf_0__0464_/a_110_47# 0.00446f
C56313 _0430_ _0438_ 0.04052f
C56314 _0476_ _0559_/a_240_47# 0.00544f
C56315 _0473_ _1040_/a_1059_315# 0
C56316 _0195_ net111 0
C56317 VPWR _0621_/a_35_297# 0.22589f
C56318 _0625_/a_59_75# net212 0.00225f
C56319 hold66/a_49_47# net150 0.0124f
C56320 VPWR net80 0.36473f
C56321 _0305_ net229 0.07107f
C56322 net155 _0570_/a_27_297# 0
C56323 _0195_ _0570_/a_109_297# 0.05702f
C56324 net102 _0347_ 0
C56325 _0720_/a_68_297# net116 0.00353f
C56326 _0140_ _1042_/a_1059_315# 0
C56327 _0460_ hold93/a_285_47# 0.02689f
C56328 VPWR _1044_/a_1059_315# 0.39816f
C56329 _0179_ _0260_ 0
C56330 hold100/a_49_47# _0219_ 0
C56331 VPWR _0149_ 0.46348f
C56332 _0225_ _0600_/a_103_199# 0.13775f
C56333 _0476_ net29 0
C56334 _0732_/a_80_21# clkbuf_0__0460_/a_110_47# 0.00119f
C56335 _1020_/a_193_47# acc0.A\[21\] 0
C56336 _0982_/a_891_413# _0345_ 0.01909f
C56337 net36 _0177_ 0.19128f
C56338 _0390_ _0773_/a_285_297# 0
C56339 _1000_/a_1059_315# _0216_ 0
C56340 _1001_/a_1059_315# _0461_ 0.00876f
C56341 _0643_/a_253_297# _0643_/a_253_47# 0.00137f
C56342 _0786_/a_217_297# _0421_ 0
C56343 _0606_/a_109_53# _0754_/a_240_47# 0
C56344 _1027_/a_891_413# _1027_/a_975_413# 0.00851f
C56345 _1027_/a_381_47# _1027_/a_561_413# 0.00123f
C56346 _0181_ _1067_/a_193_47# 0
C56347 hold8/a_285_47# clknet_1_1__leaf__0462_ 0.00568f
C56348 acc0.A\[16\] _0998_/a_193_47# 0
C56349 net10 _0140_ 0.14842f
C56350 net101 _1019_/a_27_47# 0
C56351 _0233_ _0222_ 0.10723f
C56352 _0749_/a_81_21# _0749_/a_299_297# 0.08213f
C56353 net36 _0112_ 0
C56354 clknet_1_0__leaf__0462_ _1023_/a_634_159# 0.00275f
C56355 acc0.A\[8\] _0088_ 0.02301f
C56356 hold57/a_285_47# clknet_1_0__leaf__0463_ 0
C56357 _0143_ net11 0
C56358 net248 _0442_ 0
C56359 _0195_ hold50/a_285_47# 0
C56360 clknet_1_1__leaf__0460_ acc0.A\[27\] 0.83836f
C56361 clknet_1_0__leaf__0464_ _1061_/a_634_159# 0
C56362 net133 _1061_/a_27_47# 0
C56363 net119 comp0.B\[3\] 0
C56364 clkbuf_0__0460_/a_110_47# clkbuf_1_0__f__0460_/a_110_47# 0.00994f
C56365 clkload2/a_110_47# net135 0
C56366 hold20/a_285_47# hold12/a_391_47# 0
C56367 clknet_0__0458_ _0272_ 0.00117f
C56368 _0678_/a_68_297# _0678_/a_150_297# 0.00477f
C56369 _1065_/a_466_413# _0161_ 0.00151f
C56370 control0.reset _1063_/a_27_47# 0
C56371 _1035_/a_891_413# _1035_/a_1017_47# 0.00617f
C56372 _1035_/a_193_47# _0133_ 0.51757f
C56373 _1035_/a_634_159# net121 0
C56374 _0949_/a_59_75# VPWR 0.20564f
C56375 clknet_1_0__leaf__0465_ _0835_/a_215_47# 0.00305f
C56376 _0358_ _0729_/a_68_297# 0.11143f
C56377 _0390_ _0350_ 0.09763f
C56378 hold39/a_285_47# _1034_/a_193_47# 0.00758f
C56379 hold39/a_49_47# _1034_/a_634_159# 0.00124f
C56380 hold39/a_391_47# _1034_/a_27_47# 0
C56381 _1035_/a_381_47# B[15] 0
C56382 _0410_ _0219_ 0
C56383 _1058_/a_27_47# _1058_/a_193_47# 0.96639f
C56384 _0218_ _0308_ 0
C56385 clkbuf_0__0460_/a_110_47# _0250_ 0.02331f
C56386 _0322_ _0690_/a_68_297# 0.15846f
C56387 input23/a_75_212# B[15] 0.18534f
C56388 _1000_/a_975_413# _0247_ 0
C56389 _1000_/a_891_413# _0240_ 0
C56390 _1051_/a_634_159# _0172_ 0.04621f
C56391 comp0.B\[2\] _0562_/a_68_297# 0
C56392 _0789_/a_75_199# net41 0
C56393 _0172_ _1045_/a_1059_315# 0
C56394 _0293_ _0425_ 0.00104f
C56395 _0983_/a_27_47# _0082_ 0
C56396 _0558_/a_68_297# _1035_/a_193_47# 0
C56397 _0450_ _0219_ 0.02195f
C56398 _1030_/a_466_413# _0334_ 0
C56399 _0252_ _0988_/a_381_47# 0
C56400 net44 _0607_/a_109_297# 0.01493f
C56401 _1011_/a_466_413# _0726_/a_240_47# 0
C56402 _0343_ hold91/a_285_47# 0.00386f
C56403 clknet_1_0__leaf__0465_ _0523_/a_299_297# 0.00164f
C56404 _1033_/a_634_159# _1065_/a_1059_315# 0
C56405 clknet_1_1__leaf__0460_ _0364_ 0.00513f
C56406 net152 _1043_/a_466_413# 0
C56407 _0402_ _0301_ 0.00187f
C56408 _0182_ _1015_/a_27_47# 0
C56409 _0387_ clkbuf_0__0461_/a_110_47# 0
C56410 _0966_/a_109_297# _0482_ 0
C56411 _1052_/a_193_47# net148 0
C56412 _0786_/a_80_21# _0809_/a_299_297# 0
C56413 net145 _0185_ 0.00375f
C56414 pp[8] net141 0.06223f
C56415 net55 hold77/a_49_47# 0.35361f
C56416 _0160_ hold84/a_285_47# 0.00477f
C56417 net22 _0159_ 0
C56418 _1041_/a_381_47# net174 0
C56419 net56 _0727_/a_193_47# 0
C56420 _0179_ _0524_/a_27_297# 0.00984f
C56421 _0255_ clkbuf_1_0__f__0465_/a_110_47# 0.12663f
C56422 net125 _1061_/a_561_413# 0
C56423 _0839_/a_109_297# VPWR 0.0043f
C56424 pp[15] _0218_ 0.04412f
C56425 _0398_ _1016_/a_1059_315# 0
C56426 _0466_ _0162_ 0
C56427 clknet_1_1__leaf__0460_ _0110_ 0
C56428 net150 acc0.A\[22\] 0
C56429 clknet_1_0__leaf__0460_ _0161_ 0
C56430 _0577_/a_373_47# _0120_ 0
C56431 comp0.B\[10\] _1061_/a_27_47# 0.00274f
C56432 net156 _1026_/a_634_159# 0
C56433 hold65/a_49_47# _0369_ 0.01373f
C56434 _0195_ _1018_/a_466_413# 0.02373f
C56435 _0553_/a_149_47# net171 0.01241f
C56436 net58 _0988_/a_466_413# 0.0047f
C56437 _0199_ _0171_ 0.00439f
C56438 _0467_ _1067_/a_1059_315# 0
C56439 _0794_/a_326_47# _0405_ 0
C56440 _0277_ _0792_/a_80_21# 0
C56441 net208 hold62/a_391_47# 0.039f
C56442 _0195_ _1049_/a_193_47# 0
C56443 hold15/a_49_47# net162 0
C56444 hold15/a_391_47# acc0.A\[31\] 0
C56445 _1038_/a_27_47# _0176_ 0.03734f
C56446 _0645_/a_285_47# _0302_ 0.00861f
C56447 _0183_ net151 0.089f
C56448 output43/a_27_47# pp[16] 0.15883f
C56449 _0426_ net67 0
C56450 _0563_/a_240_47# _0173_ 0.01647f
C56451 _0563_/a_245_297# _0208_ 0.00291f
C56452 net55 _0353_ 0
C56453 _0227_ _0219_ 0.19777f
C56454 _0996_/a_27_47# clkbuf_0__0459_/a_110_47# 0.0161f
C56455 clknet_1_0__leaf__0463_ _0159_ 0.04716f
C56456 _0326_ _0462_ 0.00202f
C56457 net148 net12 0
C56458 net175 net170 0
C56459 clknet_1_0__leaf__0459_ _0350_ 0.04004f
C56460 net59 _1012_/a_27_47# 0.00306f
C56461 _0635_/a_27_47# _0465_ 0.00337f
C56462 _0296_ net228 0
C56463 net64 _0088_ 0
C56464 clkbuf_1_0__f__0462_/a_110_47# _0320_ 0
C56465 _0475_ _0214_ 0.08711f
C56466 net211 _1019_/a_1059_315# 0.02973f
C56467 _0995_/a_27_47# pp[14] 0.00265f
C56468 _0995_/a_891_413# output41/a_27_47# 0
C56469 _0995_/a_634_159# net41 0
C56470 _0800_/a_240_47# _0400_ 0
C56471 net180 B[7] 0
C56472 _0520_/a_109_297# net168 0.0015f
C56473 _0798_/a_113_297# _0345_ 0.00145f
C56474 _0538_/a_51_297# _0174_ 0.09446f
C56475 _0343_ _0670_/a_215_47# 0
C56476 _0401_ clknet_1_1__leaf__0465_ 0.08044f
C56477 _0696_/a_109_297# _0328_ 0.01233f
C56478 net45 _1013_/a_975_413# 0
C56479 net67 _0185_ 0.00349f
C56480 _1018_/a_891_413# _0247_ 0
C56481 hold91/a_49_47# net5 0.03309f
C56482 hold35/a_391_47# net66 0
C56483 _0972_/a_250_297# _0164_ 0
C56484 _0336_ hold61/a_391_47# 0.01588f
C56485 clknet_1_0__leaf__0465_ _0172_ 0.05502f
C56486 _1043_/a_193_47# _1042_/a_891_413# 0
C56487 _1043_/a_466_413# _1042_/a_466_413# 0.00504f
C56488 _1043_/a_891_413# _1042_/a_193_47# 0
C56489 net116 hold92/a_285_47# 0
C56490 net236 _0162_ 0
C56491 clkbuf_0__0463_/a_110_47# net29 0
C56492 _0244_ VPWR 1.06061f
C56493 _0343_ _0247_ 0.02031f
C56494 _0642_/a_215_297# _0989_/a_193_47# 0
C56495 _0642_/a_298_297# _0989_/a_27_47# 0
C56496 _0759_/a_113_47# _0219_ 0
C56497 pp[27] _1030_/a_634_159# 0
C56498 net144 _0156_ 0.01235f
C56499 _0181_ net229 0
C56500 _1020_/a_27_47# hold55/a_391_47# 0
C56501 _0627_/a_215_53# _0627_/a_369_297# 0.00854f
C56502 _0627_/a_109_93# _0627_/a_297_297# 0
C56503 _0404_ _0347_ 0.11776f
C56504 _0352_ _0754_/a_51_297# 0.12157f
C56505 _0984_/a_27_47# _0983_/a_193_47# 0
C56506 _0984_/a_193_47# _0983_/a_27_47# 0
C56507 _0742_/a_384_47# _0315_ 0.0093f
C56508 net46 _1006_/a_193_47# 0
C56509 _0751_/a_111_297# net46 0
C56510 _1039_/a_27_47# comp0.B\[10\] 0
C56511 clknet_1_1__leaf__0460_ _1010_/a_193_47# 0.04634f
C56512 acc0.A\[29\] hold95/a_285_47# 0.04981f
C56513 _0677_/a_285_47# _0240_ 0
C56514 _0343_ _0707_/a_315_47# 0
C56515 net10 _1043_/a_634_159# 0.00423f
C56516 hold21/a_49_47# hold22/a_49_47# 0.0024f
C56517 _0234_ _0596_/a_59_75# 0
C56518 _0107_ _0371_ 0
C56519 _0472_ control0.reset 0
C56520 _0453_ _0350_ 0
C56521 _0714_/a_240_47# _1031_/a_27_47# 0
C56522 net63 _0830_/a_510_47# 0
C56523 _0485_ _1064_/a_1059_315# 0.01196f
C56524 _0487_ _1064_/a_466_413# 0
C56525 hold92/a_49_47# hold92/a_391_47# 0.00188f
C56526 _0162_ _1064_/a_193_47# 0.2458f
C56527 net135 _0148_ 0
C56528 _0549_/a_150_297# _0208_ 0
C56529 hold52/a_49_47# _0123_ 0.02533f
C56530 _0747_/a_215_47# _0219_ 0.00115f
C56531 clknet_1_1__leaf__0463_ _0175_ 0.68961f
C56532 _1059_/a_561_413# VPWR 0.00322f
C56533 _1026_/a_381_47# net112 0
C56534 _1026_/a_634_159# acc0.A\[26\] 0
C56535 control0.count\[3\] _1005_/a_193_47# 0
C56536 _0465_ _1047_/a_891_413# 0.00676f
C56537 hold10/a_49_47# _0145_ 0
C56538 _1072_/a_466_413# _0486_ 0
C56539 _0376_ net91 0
C56540 _0472_ _1061_/a_891_413# 0
C56541 hold14/a_285_47# _1035_/a_27_47# 0
C56542 hold14/a_49_47# _1035_/a_193_47# 0
C56543 _0356_ _0725_/a_80_21# 0
C56544 _0415_ _0419_ 0
C56545 _0817_/a_368_297# _0817_/a_266_47# 0.00153f
C56546 clknet_1_1__leaf__0460_ _1009_/a_634_159# 0.01274f
C56547 _0337_ _0348_ 0.28328f
C56548 acc0.A\[19\] _0771_/a_215_297# 0.01616f
C56549 _1020_/a_1059_315# _0099_ 0
C56550 _0118_ _0772_/a_79_21# 0
C56551 clknet_1_1__leaf__0458_ _0988_/a_193_47# 0
C56552 _0323_ _0324_ 0.2698f
C56553 _0399_ clkbuf_1_1__f__0458_/a_110_47# 0.00475f
C56554 acc0.A\[2\] _1047_/a_891_413# 0
C56555 net110 _0122_ 0.00195f
C56556 _1024_/a_1017_47# acc0.A\[24\] 0
C56557 _0542_/a_149_47# net20 0.02838f
C56558 _0141_ _0540_/a_51_297# 0
C56559 _0854_/a_79_21# net104 0
C56560 _0081_ _1018_/a_466_413# 0
C56561 _0294_ _0346_ 0.0306f
C56562 pp[26] _0571_/a_27_297# 0.05721f
C56563 clknet_0__0465_ acc0.A\[6\] 0.00265f
C56564 hold66/a_391_47# net213 0.13565f
C56565 hold76/a_49_47# _0241_ 0.00215f
C56566 _0226_ _0345_ 0
C56567 _0789_/a_544_297# _0405_ 0
C56568 _0850_/a_68_297# _0465_ 0.00344f
C56569 _0736_/a_56_297# _0370_ 0
C56570 net182 net66 0
C56571 _0662_/a_384_47# _0259_ 0.00921f
C56572 _0343_ _0455_ 0
C56573 _0251_ _0186_ 0
C56574 acc0.A\[11\] net37 1.03632f
C56575 net8 _0175_ 0
C56576 _0174_ _1040_/a_381_47# 0.00133f
C56577 _0136_ _1040_/a_193_47# 0
C56578 _1037_/a_1059_315# _1037_/a_891_413# 0.31086f
C56579 _1037_/a_193_47# _1037_/a_975_413# 0
C56580 _1037_/a_466_413# _1037_/a_381_47# 0.03733f
C56581 hold21/a_285_47# net140 0
C56582 _0716_/a_27_47# _0302_ 0
C56583 _0305_ _0678_/a_68_297# 0
C56584 _0183_ _0378_ 0
C56585 comp0.B\[10\] _1040_/a_975_413# 0.00106f
C56586 net59 _1030_/a_27_47# 0.00401f
C56587 input11/a_75_212# A[7] 0
C56588 _0195_ net85 0
C56589 VPWR _1005_/a_1059_315# 0.409f
C56590 clkbuf_1_0__f__0459_/a_110_47# acc0.A\[16\] 0.00322f
C56591 _0234_ _0216_ 0
C56592 _0790_/a_117_297# _0406_ 0
C56593 _0731_/a_299_297# VPWR 0.28408f
C56594 _0790_/a_285_47# acc0.A\[15\] 0
C56595 net183 _0473_ 0.00572f
C56596 VPWR _0519_/a_384_47# 0.00139f
C56597 acc0.A\[18\] _0774_/a_68_297# 0.001f
C56598 _0228_ hold3/a_391_47# 0.01674f
C56599 clknet_1_1__leaf__0458_ net72 0.12116f
C56600 VPWR _0847_/a_109_297# 0.0043f
C56601 _0369_ _0114_ 0.00158f
C56602 _1054_/a_381_47# _0180_ 0.01645f
C56603 _0336_ clknet_1_1__leaf__0462_ 0
C56604 hold30/a_285_47# _1023_/a_466_413# 0
C56605 hold30/a_49_47# _1023_/a_1059_315# 0
C56606 hold30/a_391_47# _1023_/a_634_159# 0
C56607 clknet_1_0__leaf__0462_ _0377_ 0
C56608 _0555_/a_240_47# net26 0
C56609 _0579_/a_27_297# _0721_/a_27_47# 0
C56610 _0243_ _0386_ 0.00443f
C56611 _0390_ _0244_ 0
C56612 output56/a_27_47# _1030_/a_381_47# 0
C56613 pp[28] _1030_/a_193_47# 0
C56614 _1038_/a_1059_315# net8 0
C56615 net224 _0370_ 0
C56616 _0176_ _1043_/a_592_47# 0
C56617 _0337_ acc0.A\[31\] 0.00376f
C56618 net58 _0186_ 0.02058f
C56619 VPWR _0765_/a_79_21# 0.44727f
C56620 _1039_/a_561_413# _0473_ 0.00114f
C56621 _0625_/a_59_75# _0989_/a_891_413# 0
C56622 _0127_ net114 0.00226f
C56623 _0958_/a_197_47# _0471_ 0.00749f
C56624 _0216_ clknet_0__0460_ 0.00242f
C56625 net9 net10 0.12368f
C56626 _0366_ acc0.A\[26\] 0
C56627 _0338_ _0333_ 0.00572f
C56628 _0811_/a_81_21# net228 0.00503f
C56629 _0963_/a_35_297# _0977_/a_75_212# 0.08511f
C56630 _0275_ _0817_/a_81_21# 0
C56631 _0198_ _0531_/a_109_297# 0.01875f
C56632 _0532_/a_81_21# net175 0.04844f
C56633 _0833_/a_79_21# _0434_ 0
C56634 _1049_/a_193_47# _1048_/a_193_47# 0.00549f
C56635 _1049_/a_27_47# _1048_/a_634_159# 0.00133f
C56636 _1049_/a_634_159# _1048_/a_27_47# 0
C56637 net53 _1026_/a_466_413# 0
C56638 hold33/a_285_47# clknet_1_0__leaf__0463_ 0.00753f
C56639 hold44/a_49_47# net191 0
C56640 VPWR _1011_/a_561_413# 0.00213f
C56641 hold97/a_391_47# net244 0.14844f
C56642 clkbuf_0__0457_/a_110_47# _0345_ 0.00945f
C56643 VPWR _1006_/a_634_159# 0.20288f
C56644 _0476_ comp0.B\[6\] 0.08328f
C56645 _0266_ acc0.A\[1\] 0.10867f
C56646 _0751_/a_183_297# VPWR 0
C56647 net37 hold81/a_391_47# 0.05456f
C56648 _1055_/a_634_159# A[10] 0
C56649 _0736_/a_311_297# _0350_ 0.00109f
C56650 _0307_ _0396_ 0
C56651 _0195_ _1030_/a_1059_315# 0.00224f
C56652 _0216_ _1030_/a_634_159# 0
C56653 net48 _1005_/a_1059_315# 0.01636f
C56654 VPWR _0986_/a_634_159# 0.18625f
C56655 _0289_ net67 0.21038f
C56656 _0550_/a_245_297# _0176_ 0
C56657 _0714_/a_512_297# _0345_ 0
C56658 _1019_/a_561_413# _0345_ 0.0021f
C56659 net117 _0567_/a_109_297# 0
C56660 pp[9] _1058_/a_27_47# 0
C56661 _0742_/a_81_21# _0742_/a_384_47# 0.00138f
C56662 _0951_/a_109_93# _0951_/a_209_311# 0.16762f
C56663 net237 _0324_ 0
C56664 _1013_/a_27_47# _0567_/a_27_297# 0
C56665 _0769_/a_81_21# _0462_ 0
C56666 _0715_/a_27_47# _0218_ 0
C56667 net101 comp0.B\[1\] 0
C56668 _0275_ _0084_ 0.20033f
C56669 clknet_1_0__leaf__0458_ _0842_/a_59_75# 0
C56670 control0.state\[0\] _0972_/a_346_47# 0
C56671 net48 _0765_/a_79_21# 0.14446f
C56672 _1072_/a_27_47# _1068_/a_27_47# 0
C56673 _0244_ clknet_1_0__leaf__0459_ 0.02969f
C56674 _1021_/a_27_47# net23 0
C56675 _0180_ _0522_/a_27_297# 0.10439f
C56676 _0532_/a_299_297# _0147_ 0
C56677 _0372_ control0.add 0
C56678 acc0.A\[3\] clkbuf_0__0458_/a_110_47# 0
C56679 control0.sh _0560_/a_68_297# 0
C56680 _0807_/a_68_297# _0345_ 0
C56681 _0571_/a_109_297# VPWR 0.17528f
C56682 comp0.B\[13\] _0538_/a_51_297# 0.04831f
C56683 _1001_/a_891_413# _0869_/a_27_47# 0.00229f
C56684 net95 _1009_/a_1059_315# 0
C56685 _0483_ _0468_ 0
C56686 VPWR clkbuf_1_0__f__0463_/a_110_47# 1.32044f
C56687 _0292_ acc0.A\[9\] 0.07845f
C56688 _1003_/a_1059_315# acc0.A\[21\] 0.01254f
C56689 net45 _0195_ 0.07686f
C56690 _0316_ _0323_ 0.00179f
C56691 hold75/a_285_47# _0350_ 0
C56692 _1035_/a_1059_315# _0173_ 0
C56693 _1035_/a_193_47# _0208_ 0
C56694 _0830_/a_215_47# clkbuf_1_0__f__0465_/a_110_47# 0
C56695 _1047_/a_27_47# _1047_/a_634_159# 0.14145f
C56696 net61 clkload1/Y 0.02868f
C56697 _0985_/a_1059_315# clkbuf_1_0__f__0458_/a_110_47# 0
C56698 net1 _1014_/a_381_47# 0
C56699 comp0.B\[8\] _1040_/a_1059_315# 0.12812f
C56700 _0206_ _1040_/a_466_413# 0.03279f
C56701 net178 _0181_ 0
C56702 hold97/a_49_47# _0317_ 0
C56703 clknet_1_1__leaf__0465_ hold70/a_49_47# 0
C56704 _0957_/a_32_297# _0473_ 0.1133f
C56705 net53 _0315_ 0.3321f
C56706 _0137_ clkbuf_0__0463_/a_110_47# 0.00809f
C56707 control0.add hold40/a_49_47# 0
C56708 clknet_1_0__leaf__0462_ net109 0.14186f
C56709 net60 acc0.A\[30\] 0
C56710 _1041_/a_193_47# _0174_ 0.01401f
C56711 clknet_1_0__leaf__0460_ _0758_/a_510_47# 0.00144f
C56712 _0664_/a_79_21# _0664_/a_382_297# 0.00145f
C56713 hold82/a_391_47# net229 0.13105f
C56714 _0582_/a_109_47# net221 0
C56715 clknet_1_0__leaf__0464_ net147 0
C56716 hold98/a_49_47# output60/a_27_47# 0
C56717 _0328_ hold90/a_285_47# 0
C56718 _0855_/a_81_21# _1014_/a_1059_315# 0.01733f
C56719 _0080_ hold2/a_391_47# 0
C56720 _1001_/a_193_47# clknet_1_0__leaf__0461_ 0
C56721 _0216_ net201 0.00207f
C56722 _0478_ _1071_/a_975_413# 0
C56723 _0324_ _0686_/a_27_53# 0.01038f
C56724 _1007_/a_634_159# _1007_/a_381_47# 0
C56725 _1052_/a_193_47# _1052_/a_592_47# 0
C56726 _1052_/a_466_413# _1052_/a_561_413# 0.00772f
C56727 _1052_/a_634_159# _1052_/a_975_413# 0
C56728 _0089_ clknet_1_1__leaf__0465_ 0
C56729 hold96/a_285_47# _1004_/a_27_47# 0.00197f
C56730 hold96/a_49_47# _1004_/a_193_47# 0.00129f
C56731 VPWR _0737_/a_285_297# 0.25176f
C56732 _0243_ _1006_/a_466_413# 0
C56733 _0663_/a_27_413# clkbuf_1_1__f__0465_/a_110_47# 0
C56734 _0177_ _1061_/a_27_47# 0
C56735 net186 _1034_/a_381_47# 0.11897f
C56736 _0837_/a_81_21# _0837_/a_266_47# 0.04342f
C56737 _1058_/a_634_159# _1058_/a_1017_47# 0
C56738 _1058_/a_466_413# _1058_/a_592_47# 0.00553f
C56739 _0172_ _1044_/a_466_413# 0.06385f
C56740 _1020_/a_27_47# _0352_ 0.01359f
C56741 hold69/a_49_47# _1006_/a_27_47# 0
C56742 _0477_ hold84/a_391_47# 0.00462f
C56743 _0179_ _1052_/a_466_413# 0.0363f
C56744 _0499_/a_59_75# _0465_ 0
C56745 net149 control0.reset 0
C56746 _0259_ net47 0.02284f
C56747 net216 clknet_1_0__leaf__0460_ 0
C56748 _0432_ _0829_/a_109_297# 0
C56749 net137 _0172_ 0.04956f
C56750 _0345_ net41 0.28155f
C56751 _0399_ _0408_ 0
C56752 _0212_ _1035_/a_891_413# 0.0012f
C56753 net188 acc0.A\[12\] 0
C56754 _1050_/a_466_413# net154 0.0061f
C56755 _1050_/a_27_47# net11 0.02819f
C56756 net185 input23/a_75_212# 0
C56757 hold86/a_285_47# _0346_ 0
C56758 net36 hold27/a_285_47# 0
C56759 VPWR _0722_/a_510_47# 0
C56760 _0608_/a_27_47# clknet_1_1__leaf__0461_ 0
C56761 _0262_ _0186_ 0.00322f
C56762 clk _0167_ 0
C56763 _1011_/a_592_47# _0355_ 0
C56764 _1011_/a_891_413# _0109_ 0.0502f
C56765 VPWR _1013_/a_975_413# 0.00464f
C56766 _0258_ _0218_ 0
C56767 net119 _1065_/a_1059_315# 0
C56768 _1033_/a_27_47# control0.reset 0.01875f
C56769 _1002_/a_381_47# VPWR 0.07694f
C56770 _0637_/a_56_297# _0219_ 0
C56771 hold21/a_285_47# input14/a_75_212# 0
C56772 _0195_ _0587_/a_27_47# 0
C56773 net152 net196 0
C56774 hold74/a_285_47# _0183_ 0
C56775 _0399_ _0291_ 0
C56776 _0230_ clknet_1_0__leaf__0460_ 0.00701f
C56777 _0656_/a_145_75# clknet_1_1__leaf__0465_ 0.00162f
C56778 acc0.A\[17\] _0779_/a_79_21# 0
C56779 _1054_/a_1059_315# _0152_ 0.00854f
C56780 clknet_1_0__leaf__0462_ pp[24] 0
C56781 _0369_ _0828_/a_199_47# 0
C56782 _0220_ net116 0
C56783 _0689_/a_68_297# acc0.A\[26\] 0.00149f
C56784 _1063_/a_27_47# _1063_/a_193_47# 0.96163f
C56785 net217 _0345_ 0.00303f
C56786 net206 _0611_/a_68_297# 0
C56787 _0331_ _0356_ 0
C56788 _1058_/a_466_413# _0186_ 0
C56789 _0179_ _0194_ 0
C56790 _0176_ B[6] 0.00299f
C56791 _0310_ acc0.A\[17\] 0
C56792 acc0.A\[16\] clkbuf_0__0461_/a_110_47# 0.02076f
C56793 _0399_ net166 0
C56794 clkbuf_0__0463_/a_110_47# comp0.B\[6\] 0.00138f
C56795 _0345_ hold62/a_285_47# 0.00264f
C56796 _1027_/a_1017_47# acc0.A\[26\] 0
C56797 _0422_ _0304_ 0
C56798 _0136_ _0207_ 0.1274f
C56799 net125 clknet_1_0__leaf__0464_ 0
C56800 hold80/a_49_47# hold80/a_391_47# 0.00188f
C56801 _1063_/a_891_413# _0880_/a_27_47# 0.00229f
C56802 _0592_/a_68_297# VPWR 0.15373f
C56803 net37 _0281_ 0.25626f
C56804 net46 _0103_ 0
C56805 _0974_/a_79_199# net159 0.00586f
C56806 _0197_ _1048_/a_891_413# 0
C56807 _1039_/a_27_47# _0177_ 0
C56808 net205 _1034_/a_975_413# 0
C56809 _1050_/a_27_47# hold7/a_391_47# 0
C56810 net64 _0516_/a_109_297# 0
C56811 _0217_ _0235_ 0
C56812 _0727_/a_277_47# _0221_ 0
C56813 _0984_/a_381_47# VPWR 0.07689f
C56814 net63 _0989_/a_193_47# 0.03203f
C56815 _0336_ hold92/a_49_47# 0
C56816 _0220_ hold92/a_285_47# 0.00332f
C56817 _0693_/a_68_297# _1006_/a_891_413# 0
C56818 net63 hold1/a_285_47# 0.0244f
C56819 _0172_ _0546_/a_240_47# 0.0851f
C56820 _0994_/a_975_413# _0218_ 0
C56821 _0538_/a_51_297# comp0.B\[9\] 0
C56822 pp[8] pp[9] 0.75233f
C56823 _0237_ _0754_/a_51_297# 0
C56824 hold30/a_391_47# _0377_ 0
C56825 net67 _0418_ 0
C56826 net221 net47 0
C56827 net111 _1026_/a_381_47# 0
C56828 _1011_/a_193_47# acc0.A\[29\] 0.00773f
C56829 pp[27] pp[17] 0
C56830 hold44/a_391_47# acc0.A\[28\] 0
C56831 _1004_/a_193_47# net90 0.01355f
C56832 net168 _0186_ 0.09964f
C56833 _0183_ _0583_/a_109_297# 0.05848f
C56834 hold41/a_285_47# acc0.A\[10\] 0.02416f
C56835 _0516_/a_27_297# _0290_ 0.0011f
C56836 _0369_ _0990_/a_466_413# 0
C56837 clkbuf_1_0__f__0462_/a_110_47# _1007_/a_1059_315# 0.02051f
C56838 _1002_/a_381_47# net48 0
C56839 _0429_ _0642_/a_298_297# 0
C56840 VPWR _1042_/a_1017_47# 0
C56841 _1060_/a_27_47# _1060_/a_193_47# 0.96639f
C56842 _0982_/a_561_413# _0346_ 0.0014f
C56843 hold97/a_285_47# clknet_1_1__leaf__0460_ 0.01241f
C56844 hold43/a_49_47# _1028_/a_193_47# 0
C56845 hold43/a_285_47# _1028_/a_27_47# 0
C56846 _1070_/a_193_47# _0979_/a_109_297# 0
C56847 _1070_/a_27_47# _0979_/a_109_47# 0
C56848 _0191_ _0620_/a_113_47# 0
C56849 _0191_ _0989_/a_27_47# 0
C56850 pp[26] net210 0
C56851 net54 net155 0
C56852 _1043_/a_1059_315# net128 0
C56853 _0694_/a_113_47# net52 0
C56854 _1030_/a_561_413# acc0.A\[30\] 0
C56855 _0273_ _0989_/a_891_413# 0
C56856 clknet_1_1__leaf__0463_ _0955_/a_114_297# 0
C56857 hold56/a_391_47# _1065_/a_27_47# 0
C56858 hold56/a_285_47# _1065_/a_193_47# 0
C56859 _0343_ hold31/a_391_47# 0
C56860 hold16/a_285_47# hold62/a_49_47# 0
C56861 _0988_/a_634_159# _0988_/a_592_47# 0
C56862 _0553_/a_51_297# _0553_/a_149_47# 0.02487f
C56863 output57/a_27_47# _0355_ 0
C56864 _0352_ _0219_ 0.10353f
C56865 _0181_ clkbuf_1_1__f__0457_/a_110_47# 0.15409f
C56866 _1039_/a_1059_315# _0136_ 0
C56867 output55/a_27_47# _0568_/a_109_297# 0
C56868 _1053_/a_634_159# acc0.A\[7\] 0
C56869 hold100/a_285_47# _0465_ 0.00645f
C56870 clkbuf_0_clk/a_110_47# _1062_/a_466_413# 0
C56871 clk _1062_/a_27_47# 0
C56872 net1 _1067_/a_1059_315# 0
C56873 _0357_ _0358_ 0.09288f
C56874 _0305_ _0675_/a_68_297# 0.00375f
C56875 net56 _0350_ 0.0035f
C56876 _0476_ net26 0.03812f
C56877 _0511_/a_81_21# net143 0
C56878 clknet_1_0__leaf__0461_ net107 0.23859f
C56879 _0982_/a_634_159# _0465_ 0.00233f
C56880 _0953_/a_32_297# comp0.B\[10\] 0.1511f
C56881 net10 net129 0
C56882 _1063_/a_27_47# _1062_/a_891_413# 0
C56883 _1063_/a_193_47# _1062_/a_1059_315# 0
C56884 VPWR _1014_/a_27_47# 0.61873f
C56885 net58 hold100/a_49_47# 0.02838f
C56886 acc0.A\[2\] hold100/a_285_47# 0
C56887 _0312_ _0326_ 0.40536f
C56888 _0785_/a_299_297# acc0.A\[9\] 0
C56889 _0542_/a_240_47# _0203_ 0
C56890 _0542_/a_245_297# net19 0
C56891 _0111_ _1031_/a_634_159# 0
C56892 net227 _0334_ 0.00285f
C56893 hold101/a_285_47# VPWR 0.29725f
C56894 _1056_/a_466_413# _0369_ 0
C56895 hold96/a_49_47# net199 0
C56896 net112 acc0.A\[26\] 0
C56897 _0432_ _0840_/a_150_297# 0
C56898 _0982_/a_634_159# acc0.A\[2\] 0
C56899 _0328_ clknet_0__0462_ 0.82029f
C56900 _0999_/a_381_47# _0097_ 0.11632f
C56901 _0460_ _1062_/a_1059_315# 0
C56902 _0684_/a_59_75# _0318_ 0.00285f
C56903 _0316_ _0686_/a_27_53# 0.12f
C56904 _0640_/a_109_53# net62 0
C56905 _0674_/a_113_47# net43 0
C56906 _1021_/a_634_159# _0460_ 0.00504f
C56907 _0399_ _0290_ 0.0318f
C56908 _1021_/a_1059_315# clknet_1_0__leaf__0457_ 0.00987f
C56909 _0490_ _0487_ 0
C56910 _0316_ _1008_/a_891_413# 0
C56911 _0701_/a_80_21# _0701_/a_209_297# 0.06257f
C56912 net133 _1047_/a_634_159# 0
C56913 A[14] pp[13] 0
C56914 net36 _0268_ 0
C56915 pp[26] _0125_ 0.17933f
C56916 clkbuf_0__0462_/a_110_47# _0737_/a_35_297# 0
C56917 _0626_/a_68_297# _0271_ 0.01607f
C56918 _0626_/a_150_297# _0256_ 0.0017f
C56919 acc0.A\[20\] _0218_ 0.01722f
C56920 _0580_/a_109_297# acc0.A\[19\] 0.01859f
C56921 hold67/a_49_47# _0179_ 0.00498f
C56922 net44 net59 0.52132f
C56923 _0279_ _0994_/a_381_47# 0
C56924 _0461_ _0246_ 0
C56925 _1050_/a_27_47# clknet_1_1__leaf__0458_ 0
C56926 _1008_/a_1059_315# _0739_/a_79_21# 0.00344f
C56927 clknet_1_1__leaf__0460_ _0366_ 0.15477f
C56928 _0144_ _1061_/a_193_47# 0
C56929 _0557_/a_512_297# _0175_ 0.00291f
C56930 net43 _0406_ 0
C56931 _0347_ _1008_/a_891_413# 0.00783f
C56932 _1037_/a_381_47# _0135_ 0.13111f
C56933 hold45/a_49_47# A[11] 0
C56934 _0996_/a_27_47# hold91/a_391_47# 0
C56935 _0996_/a_193_47# hold91/a_285_47# 0
C56936 _0531_/a_109_297# _1048_/a_466_413# 0
C56937 _0531_/a_27_297# _1048_/a_1059_315# 0.00131f
C56938 hold97/a_391_47# clkbuf_1_1__f__0462_/a_110_47# 0
C56939 pp[0] B[7] 0
C56940 _0195_ _0998_/a_1017_47# 0
C56941 _0236_ clknet_1_0__leaf__0460_ 0
C56942 _0644_/a_47_47# _0277_ 0.17523f
C56943 pp[30] _1030_/a_592_47# 0
C56944 hold34/a_285_47# hold34/a_391_47# 0.41909f
C56945 _0986_/a_27_47# acc0.A\[6\] 0
C56946 hold13/a_285_47# _0957_/a_32_297# 0
C56947 _0557_/a_149_47# control0.sh 0.00423f
C56948 net58 net62 0.09343f
C56949 _0664_/a_79_21# _0402_ 0.04465f
C56950 _0642_/a_215_297# _0988_/a_27_47# 0
C56951 hold9/a_49_47# clknet_1_1__leaf__0462_ 0.01484f
C56952 net58 _0450_ 0.03581f
C56953 clknet_0__0457_ _0584_/a_27_297# 0
C56954 hold18/a_391_47# VPWR 0.18821f
C56955 _0083_ _0844_/a_79_21# 0.0023f
C56956 _0728_/a_59_75# net115 0
C56957 clkbuf_1_1__f__0462_/a_110_47# net96 0
C56958 hold30/a_285_47# net177 0.01139f
C56959 _1001_/a_27_47# _0772_/a_79_21# 0.00999f
C56960 _1001_/a_634_159# _1001_/a_592_47# 0
C56961 _0235_ _0248_ 0
C56962 _0253_ net47 0
C56963 _0991_/a_27_47# _0345_ 0.00139f
C56964 _0399_ acc0.A\[1\] 0
C56965 net189 _0189_ 0
C56966 clknet_1_0__leaf__0464_ _0186_ 0.03163f
C56967 _1062_/a_1059_315# _1062_/a_891_413# 0.31086f
C56968 _1062_/a_193_47# _1062_/a_975_413# 0
C56969 _1062_/a_466_413# _1062_/a_381_47# 0.03733f
C56970 _0708_/a_150_297# pp[31] 0
C56971 _0239_ acc0.A\[17\] 0.03965f
C56972 _0348_ _0333_ 0.02008f
C56973 output56/a_27_47# _0568_/a_27_297# 0
C56974 _0487_ hold93/a_49_47# 0
C56975 clkbuf_1_1__f__0463_/a_110_47# comp0.B\[0\] 0
C56976 _1029_/a_27_47# clknet_1_1__leaf__0462_ 0.00782f
C56977 _1011_/a_891_413# _0725_/a_80_21# 0
C56978 _1011_/a_1059_315# _0725_/a_209_297# 0.00125f
C56979 _0675_/a_68_297# _0675_/a_150_297# 0.00477f
C56980 _0992_/a_634_159# net228 0.00125f
C56981 _0869_/a_27_47# net149 0
C56982 net199 net90 0
C56983 _1021_/a_27_47# _1021_/a_891_413# 0.03224f
C56984 _1021_/a_193_47# _1021_/a_1059_315# 0.03405f
C56985 _1021_/a_634_159# _1021_/a_466_413# 0.23992f
C56986 _0831_/a_285_47# _0253_ 0
C56987 pp[17] _0216_ 0
C56988 _1003_/a_891_413# net49 0.00823f
C56989 _0518_/a_27_297# clknet_1_1__leaf__0458_ 0.0154f
C56990 _0146_ net9 0.02192f
C56991 _1049_/a_27_47# net134 0.04128f
C56992 clkbuf_1_0__f__0459_/a_110_47# _0506_/a_299_297# 0
C56993 net144 output37/a_27_47# 0.00114f
C56994 _0195_ VPWR 10.62823f
C56995 _1037_/a_1059_315# net27 0
C56996 _0476_ hold84/a_285_47# 0.02821f
C56997 control0.state\[1\] _0971_/a_299_297# 0
C56998 VPWR net92 0.35047f
C56999 _0791_/a_113_297# net41 0
C57000 net191 _1008_/a_193_47# 0
C57001 _0205_ _0545_/a_68_297# 0.12369f
C57002 hold43/a_285_47# _1029_/a_381_47# 0
C57003 _0536_/a_149_47# _0953_/a_32_297# 0
C57004 hold87/a_49_47# hold59/a_391_47# 0
C57005 net117 _1031_/a_27_47# 0.22435f
C57006 _0963_/a_285_297# control0.count\[0\] 0.06868f
C57007 net194 net21 0
C57008 A[12] net37 0.10612f
C57009 VPWR _0548_/a_245_297# 0.00515f
C57010 _0856_/a_510_47# VPWR 0
C57011 clkbuf_1_0__f__0465_/a_110_47# _0989_/a_27_47# 0
C57012 clkbuf_1_0__f__0465_/a_110_47# hold1/a_49_47# 0.00147f
C57013 net34 _0975_/a_145_75# 0
C57014 _0968_/a_193_297# _0486_ 0.01657f
C57015 clknet_1_1__leaf__0464_ _1043_/a_891_413# 0.05311f
C57016 _0350_ _0345_ 0.58465f
C57017 _0752_/a_27_413# _0378_ 0
C57018 _0234_ _0756_/a_377_297# 0
C57019 _0216_ _1015_/a_193_47# 0
C57020 clkload1/Y _0431_ 0.00305f
C57021 _0433_ _0825_/a_68_297# 0.11687f
C57022 _0111_ _0345_ 0.00101f
C57023 _0083_ _0846_/a_240_47# 0
C57024 _0317_ _0685_/a_150_297# 0
C57025 net45 _0779_/a_510_47# 0
C57026 _0763_/a_109_47# _0462_ 0
C57027 A[13] _0668_/a_382_297# 0
C57028 clknet_1_0__leaf__0465_ _0437_ 0
C57029 _0092_ _0994_/a_1059_315# 0
C57030 _0185_ net6 0.02915f
C57031 _1034_/a_634_159# clkbuf_1_1__f__0463_/a_110_47# 0.00576f
C57032 _0951_/a_368_53# comp0.B\[0\] 0.00514f
C57033 _0333_ _0332_ 0.30586f
C57034 _0343_ _0444_ 0
C57035 hold38/a_285_47# _1034_/a_27_47# 0
C57036 net187 _0902_/a_27_47# 0.00369f
C57037 _0371_ _0346_ 0.06499f
C57038 hold40/a_391_47# hold73/a_391_47# 0
C57039 _0218_ hold92/a_391_47# 0
C57040 net213 _0374_ 0
C57041 _0714_/a_149_47# _0344_ 0.00753f
C57042 hold34/a_285_47# _0181_ 0
C57043 net160 _0552_/a_68_297# 0
C57044 _0368_ _0319_ 0
C57045 acc0.A\[5\] _0150_ 0
C57046 _0307_ net43 0.25906f
C57047 net34 _0164_ 0.00115f
C57048 _0717_/a_209_297# output44/a_27_47# 0
C57049 hold29/a_49_47# _1022_/a_27_47# 0
C57050 _0324_ _0320_ 0
C57051 _0180_ _0193_ 0.02876f
C57052 _0259_ _0294_ 0.10582f
C57053 _0982_/a_193_47# _0262_ 0
C57054 _0675_/a_68_297# _0181_ 0.00984f
C57055 _0121_ clknet_1_0__leaf__0460_ 0
C57056 _1020_/a_27_47# net106 0.22672f
C57057 hold20/a_391_47# clknet_1_0__leaf_clk 0
C57058 net11 _0987_/a_27_47# 0.03793f
C57059 _0618_/a_79_21# _0618_/a_297_297# 0.01735f
C57060 _0473_ _0213_ 0.12467f
C57061 _0957_/a_32_297# _0132_ 0
C57062 _1036_/a_381_47# clknet_1_1__leaf__0463_ 0.01223f
C57063 _1036_/a_1059_315# net122 0
C57064 _1052_/a_466_413# hold83/a_49_47# 0
C57065 _0343_ _0367_ 0
C57066 _0233_ _0366_ 0.00198f
C57067 _0999_/a_27_47# _0307_ 0
C57068 _0461_ _1019_/a_1059_315# 0.01442f
C57069 hold68/a_285_47# _0222_ 0
C57070 _0101_ _0227_ 0
C57071 _0218_ net72 0.10234f
C57072 hold96/a_49_47# VPWR 0.27895f
C57073 _0678_/a_68_297# clknet_1_1__leaf__0461_ 0
C57074 VPWR _0852_/a_35_297# 0.16009f
C57075 clknet_0__0458_ _0990_/a_193_47# 0
C57076 _0644_/a_47_47# _0296_ 0
C57077 _1001_/a_193_47# _0218_ 0
C57078 _1041_/a_193_47# comp0.B\[9\] 0
C57079 _1041_/a_1059_315# net153 0
C57080 _1041_/a_891_413# net127 0
C57081 _1047_/a_891_413# _1047_/a_975_413# 0.00851f
C57082 _1047_/a_381_47# _1047_/a_561_413# 0.00123f
C57083 net23 _0132_ 0
C57084 _1037_/a_1059_315# _0136_ 0
C57085 _1030_/a_592_47# _0339_ 0
C57086 _0206_ net174 0.01164f
C57087 _0305_ _0780_/a_285_47# 0.00135f
C57088 _0472_ _0475_ 0.12855f
C57089 _0290_ _0295_ 0.03768f
C57090 _0264_ acc0.A\[18\] 0.00217f
C57091 hold25/a_285_47# VPWR 0.30138f
C57092 net47 net74 0
C57093 _0401_ _0296_ 0
C57094 clknet_1_0__leaf_clk _0970_/a_27_297# 0
C57095 clknet_0__0465_ _0826_/a_219_297# 0.00394f
C57096 comp0.B\[1\] _0563_/a_512_297# 0
C57097 net185 _0561_/a_149_47# 0.0066f
C57098 _0270_ _0465_ 0
C57099 _0212_ _0561_/a_512_297# 0
C57100 _0961_/a_113_297# _0480_ 0.01005f
C57101 _0849_/a_79_21# _0219_ 0.13069f
C57102 _0230_ hold94/a_285_47# 0
C57103 pp[28] _0354_ 0.00748f
C57104 _0343_ _0718_/a_285_47# 0.01005f
C57105 comp0.B\[5\] _0176_ 0.21833f
C57106 hold41/a_285_47# _0188_ 0.05275f
C57107 _0217_ _1018_/a_891_413# 0.0151f
C57108 _0183_ _1018_/a_466_413# 0
C57109 input28/a_75_212# _0175_ 0
C57110 _0567_/a_109_297# _0704_/a_68_297# 0
C57111 hold85/a_49_47# _0959_/a_80_21# 0
C57112 _1007_/a_381_47# net93 0
C57113 hold22/a_285_47# _0152_ 0.00315f
C57114 _0389_ _0216_ 0.0266f
C57115 _0464_ _0196_ 0
C57116 _0536_/a_245_297# _0473_ 0.00125f
C57117 _0858_/a_27_47# _0465_ 0.00544f
C57118 _0680_/a_80_21# net95 0
C57119 net243 _1004_/a_891_413# 0.04439f
C57120 VPWR _0081_ 0.35761f
C57121 net12 hold83/a_391_47# 0.0158f
C57122 _0525_/a_299_297# acc0.A\[6\] 0
C57123 _0194_ hold83/a_49_47# 0
C57124 _0837_/a_585_47# _0442_ 0
C57125 net186 comp0.B\[2\] 0.0032f
C57126 _0411_ _0798_/a_113_297# 0.00761f
C57127 _0343_ _0217_ 0.39693f
C57128 _0305_ _0677_/a_47_47# 0.01689f
C57129 _0446_ _0261_ 0.22858f
C57130 _0502_/a_27_47# _0180_ 0.24195f
C57131 _0570_/a_109_297# net156 0.00104f
C57132 _0126_ _1027_/a_1059_315# 0
C57133 input19/a_75_212# net19 0.10859f
C57134 B[11] _0203_ 0
C57135 _0767_/a_59_75# _0306_ 0
C57136 _0502_/a_27_47# net218 0
C57137 hold7/a_285_47# _0987_/a_193_47# 0.00166f
C57138 hold7/a_49_47# _0987_/a_634_159# 0.0037f
C57139 hold7/a_391_47# _0987_/a_27_47# 0.00109f
C57140 _0629_/a_59_75# _0458_ 0.00247f
C57141 acc0.A\[2\] _0858_/a_27_47# 0
C57142 _1057_/a_193_47# net37 0
C57143 net30 clkbuf_1_0__f__0463_/a_110_47# 0
C57144 _0267_ _0265_ 0.14694f
C57145 net208 _0334_ 0
C57146 _0216_ _0355_ 0.00178f
C57147 hold58/a_285_47# _0175_ 0
C57148 VPWR _0505_/a_373_47# 0
C57149 _0172_ _0148_ 0
C57150 _0294_ net221 0.02723f
C57151 hold24/a_49_47# VPWR 0.33101f
C57152 hold42/a_49_47# net67 0
C57153 clknet_1_0__leaf__0461_ _0208_ 0.13359f
C57154 _1057_/a_466_413# net67 0.01658f
C57155 _0757_/a_68_297# acc0.A\[23\] 0.01322f
C57156 hold25/a_49_47# _0550_/a_51_297# 0
C57157 _1038_/a_27_47# net28 0
C57158 net61 _0989_/a_1017_47# 0
C57159 _0243_ _0240_ 0.06274f
C57160 _0179_ _0517_/a_299_297# 0.0536f
C57161 _0983_/a_381_47# _0081_ 0.13242f
C57162 net36 clkbuf_1_0__f__0461_/a_110_47# 0
C57163 _0243_ _0369_ 0
C57164 _1063_/a_466_413# _1063_/a_592_47# 0.00553f
C57165 _1063_/a_634_159# _1063_/a_1017_47# 0
C57166 _0833_/a_215_47# _0988_/a_193_47# 0
C57167 _0573_/a_27_47# _0584_/a_109_297# 0
C57168 _0965_/a_285_47# _1072_/a_27_47# 0
C57169 net233 _0465_ 0.01576f
C57170 VPWR net90 0.94676f
C57171 _0636_/a_59_75# _0844_/a_297_47# 0
C57172 _0399_ net77 0
C57173 hold19/a_285_47# _0115_ 0
C57174 _1037_/a_592_47# _0208_ 0
C57175 net133 _0174_ 0
C57176 _0400_ _0791_/a_199_47# 0.01074f
C57177 acc0.A\[20\] _0099_ 0
C57178 _0626_/a_68_297# clknet_1_0__leaf__0465_ 0
C57179 _0985_/a_1059_315# acc0.A\[15\] 0
C57180 _0839_/a_109_297# _0345_ 0.00382f
C57181 _0585_/a_27_297# _0585_/a_109_47# 0.00393f
C57182 _0121_ _0576_/a_109_297# 0.0036f
C57183 _1071_/a_27_47# _0976_/a_76_199# 0
C57184 _0556_/a_68_297# _0175_ 0.10319f
C57185 _0982_/a_27_47# net47 0
C57186 hold76/a_49_47# _0352_ 0
C57187 net233 acc0.A\[2\] 0
C57188 _0172_ input31/a_75_212# 0
C57189 clknet_1_0__leaf__0464_ _1050_/a_634_159# 0.00109f
C57190 _0305_ hold82/a_285_47# 0.01664f
C57191 _0349_ _1012_/a_27_47# 0
C57192 VPWR _1048_/a_193_47# 0.3116f
C57193 _0535_/a_68_297# comp0.B\[10\] 0.00271f
C57194 _0349_ _0330_ 0
C57195 net198 _0542_/a_51_297# 0.10395f
C57196 _0544_/a_512_297# _0203_ 0
C57197 _0183_ acc0.A\[13\] 0.09129f
C57198 net232 _1062_/a_193_47# 0.0031f
C57199 _0144_ clkbuf_0__0464_/a_110_47# 0
C57200 _0195_ clknet_1_0__leaf__0459_ 0.02725f
C57201 _1028_/a_466_413# net113 0
C57202 _1028_/a_891_413# clknet_1_1__leaf__0462_ 0.00801f
C57203 hold57/a_49_47# _0175_ 0
C57204 hold46/a_285_47# _0473_ 0
C57205 clknet_0__0459_ _0302_ 0.1782f
C57206 _0191_ net11 0
C57207 net214 acc0.A\[8\] 0
C57208 _0483_ _1071_/a_466_413# 0
C57209 _0530_/a_299_297# clknet_1_1__leaf__0457_ 0
C57210 _0556_/a_150_297# control0.sh 0
C57211 _0237_ _0219_ 0.35678f
C57212 _0429_ _0191_ 0
C57213 hold47/a_391_47# _0186_ 0
C57214 _0427_ clkbuf_0__0465_/a_110_47# 0
C57215 _0819_/a_384_47# clknet_0__0465_ 0
C57216 net111 acc0.A\[26\] 0
C57217 clknet_1_1__leaf__0460_ acc0.A\[24\] 0.03192f
C57218 _0195_ _0569_/a_109_47# 0.00382f
C57219 _0216_ _0569_/a_27_297# 0.19926f
C57220 _0570_/a_109_297# acc0.A\[26\] 0.00413f
C57221 _0369_ _0088_ 0.02952f
C57222 VPWR _1010_/a_891_413# 0.21503f
C57223 _0190_ _0290_ 0
C57224 _1000_/a_27_47# _1000_/a_891_413# 0.03089f
C57225 _1000_/a_193_47# _1000_/a_1059_315# 0.03405f
C57226 _1000_/a_634_159# _1000_/a_466_413# 0.23992f
C57227 _1060_/a_466_413# _1060_/a_592_47# 0.00553f
C57228 _1060_/a_634_159# _1060_/a_1017_47# 0
C57229 _0350_ net52 0.02715f
C57230 _1051_/a_27_47# net154 0.02098f
C57231 hold57/a_285_47# control0.sh 0.04397f
C57232 net114 _1008_/a_561_413# 0
C57233 net4 acc0.A\[10\] 0.31579f
C57234 VPWR _0979_/a_109_297# 0.19578f
C57235 _1051_/a_891_413# _0346_ 0
C57236 _0192_ _0520_/a_373_47# 0
C57237 _0151_ _0520_/a_27_297# 0.05365f
C57238 net230 _0520_/a_109_47# 0
C57239 _0462_ _0616_/a_215_47# 0.0016f
C57240 _0457_ net149 0
C57241 _0346_ clkbuf_1_1__f__0458_/a_110_47# 0
C57242 _1039_/a_592_47# comp0.B\[9\] 0
C57243 _0257_ clkbuf_1_0__f__0465_/a_110_47# 0.02921f
C57244 clknet_1_1__leaf__0458_ _0987_/a_27_47# 0.00146f
C57245 VPWR _0846_/a_149_47# 0
C57246 _0343_ _0742_/a_299_297# 0.00955f
C57247 _0467_ _0163_ 0.06756f
C57248 _0568_/a_109_297# acc0.A\[30\] 0
C57249 _0805_/a_109_47# VPWR 0
C57250 _0553_/a_245_297# _0136_ 0
C57251 _0399_ _0986_/a_1059_315# 0.00229f
C57252 _0347_ _0320_ 0.01844f
C57253 _0973_/a_27_297# _1063_/a_1059_315# 0.01884f
C57254 VPWR _1009_/a_381_47# 0.07658f
C57255 hold36/a_285_47# clknet_1_1__leaf__0464_ 0
C57256 hold14/a_285_47# _0173_ 0
C57257 acc0.A\[12\] hold81/a_49_47# 0.31715f
C57258 _0446_ net47 0
C57259 _0174_ comp0.B\[10\] 0.83077f
C57260 clkbuf_1_0__f__0457_/a_110_47# net87 0
C57261 _0857_/a_27_47# _1033_/a_891_413# 0
C57262 _0457_ _1033_/a_27_47# 0
C57263 clknet_1_0__leaf__0460_ _0380_ 0.00723f
C57264 _0963_/a_35_297# _0963_/a_117_297# 0.00641f
C57265 _0401_ _0811_/a_81_21# 0
C57266 hold27/a_285_47# _1039_/a_27_47# 0
C57267 net68 _0465_ 0.00113f
C57268 _0195_ _0453_ 0.0017f
C57269 _0216_ _0266_ 0
C57270 _0227_ net35 0.00173f
C57271 _0233_ _0378_ 0.00878f
C57272 _0375_ _0183_ 0
C57273 _0583_/a_27_297# net165 0.05973f
C57274 _0236_ hold94/a_285_47# 0.00465f
C57275 _1071_/a_975_413# VPWR 0.00485f
C57276 net240 _0880_/a_27_47# 0
C57277 _0973_/a_373_47# _0460_ 0
C57278 net195 _0141_ 0
C57279 _1056_/a_193_47# net178 0
C57280 hold37/a_391_47# clkbuf_0__0464_/a_110_47# 0.00111f
C57281 _0343_ _0248_ 0.42185f
C57282 _0330_ _0701_/a_209_297# 0.03541f
C57283 _0216_ _0567_/a_109_297# 0.00669f
C57284 _0573_/a_27_47# VPWR 0.4025f
C57285 _0195_ _0567_/a_373_47# 0.00228f
C57286 _0985_/a_1059_315# _0179_ 0.02353f
C57287 acc0.A\[26\] hold50/a_285_47# 0
C57288 clknet_1_0__leaf__0457_ net223 0.08277f
C57289 acc0.A\[15\] acc0.A\[13\] 0.21716f
C57290 clknet_1_1__leaf__0462_ _0739_/a_79_21# 0.00805f
C57291 _0163_ comp0.B\[0\] 0.36109f
C57292 _0179_ _1049_/a_193_47# 0.29096f
C57293 _0707_/a_75_199# acc0.A\[29\] 0.00369f
C57294 _1059_/a_466_413# _0219_ 0
C57295 clknet_0__0458_ _0438_ 0.0128f
C57296 net36 _0182_ 0.01982f
C57297 _0701_/a_209_47# _0333_ 0
C57298 clkbuf_1_0__f__0458_/a_110_47# VPWR 1.18661f
C57299 _0997_/a_193_47# net41 0.04955f
C57300 _0997_/a_1059_315# output41/a_27_47# 0
C57301 _0222_ _0754_/a_51_297# 0.00757f
C57302 _0309_ acc0.A\[17\] 0.07119f
C57303 clknet_0__0464_ _1046_/a_1059_315# 0.00118f
C57304 hold11/a_49_47# net157 0.05889f
C57305 _1071_/a_193_47# clknet_0_clk 0.00414f
C57306 clknet_0__0458_ _0636_/a_59_75# 0
C57307 _1008_/a_891_413# _0106_ 0.04091f
C57308 A[11] _0156_ 0
C57309 VPWR _0954_/a_304_297# 0.00535f
C57310 hold13/a_285_47# _0213_ 0.0012f
C57311 hold13/a_49_47# _0173_ 0.00218f
C57312 _0134_ _0175_ 0.06396f
C57313 _0585_/a_27_297# _0208_ 0
C57314 _0349_ _1030_/a_27_47# 0
C57315 net9 _1048_/a_381_47# 0
C57316 _0178_ _1047_/a_193_47# 0.04168f
C57317 clknet_1_0__leaf__0459_ _0081_ 0.00139f
C57318 _0683_/a_113_47# clknet_1_0__leaf__0460_ 0
C57319 comp0.B\[11\] _1043_/a_1059_315# 0.10769f
C57320 clkbuf_1_1__f__0465_/a_110_47# acc0.A\[9\] 0.02842f
C57321 _0677_/a_47_47# _0181_ 0.00851f
C57322 _0328_ _0687_/a_59_75# 0.00177f
C57323 _1020_/a_466_413# _0578_/a_27_297# 0
C57324 output56/a_27_47# _0725_/a_80_21# 0
C57325 clknet_0__0459_ net6 0.50209f
C57326 _0998_/a_1059_315# _0790_/a_285_297# 0
C57327 net21 _1045_/a_27_47# 0.02697f
C57328 net183 _1045_/a_193_47# 0.00154f
C57329 _0531_/a_27_297# clkbuf_1_1__f__0457_/a_110_47# 0
C57330 clknet_1_1__leaf__0459_ _0097_ 0.00287f
C57331 VPWR _1022_/a_561_413# 0.00292f
C57332 pp[30] _0568_/a_373_47# 0
C57333 hold101/a_49_47# _0172_ 0.00915f
C57334 _0650_/a_68_297# hold81/a_49_47# 0.0141f
C57335 VPWR _0779_/a_510_47# 0
C57336 _0637_/a_311_297# _0465_ 0
C57337 _0852_/a_35_297# _0453_ 0.21351f
C57338 clknet_1_1__leaf__0459_ _0993_/a_381_47# 0
C57339 _0852_/a_285_47# _0452_ 0
C57340 _0852_/a_285_297# _0266_ 0.00189f
C57341 _0993_/a_975_413# net38 0
C57342 B[14] hold6/a_391_47# 0
C57343 net22 hold6/a_285_47# 0
C57344 _0999_/a_634_159# _0999_/a_381_47# 0
C57345 _0854_/a_297_297# _0399_ 0.00153f
C57346 net17 _1063_/a_1059_315# 0.05489f
C57347 _0992_/a_634_159# _0090_ 0
C57348 _1001_/a_27_47# _1019_/a_27_47# 0.00135f
C57349 _1017_/a_634_159# _0115_ 0.00107f
C57350 _0461_ _0774_/a_68_297# 0
C57351 _0957_/a_32_297# net25 0
C57352 _0972_/a_256_47# clknet_1_1__leaf_clk 0
C57353 _0833_/a_79_21# _0186_ 0.04731f
C57354 _1001_/a_193_47# _0099_ 0.1749f
C57355 hold26/a_391_47# clkbuf_1_0__f__0463_/a_110_47# 0
C57356 _1001_/a_1059_315# net223 0.05968f
C57357 _0340_ _1031_/a_1059_315# 0
C57358 clknet_1_0__leaf__0465_ _0252_ 0
C57359 hold35/a_285_47# _0369_ 0
C57360 _0665_/a_109_297# net6 0.00357f
C57361 _0555_/a_149_47# _0957_/a_32_297# 0
C57362 net58 _0637_/a_56_297# 0
C57363 acc0.A\[3\] _0447_ 0
C57364 net120 _1034_/a_381_47# 0
C57365 _1004_/a_466_413# _0217_ 0
C57366 net205 VPWR 0.56788f
C57367 net159 net17 0
C57368 _1033_/a_27_47# _0475_ 0
C57369 _0423_ _0813_/a_109_297# 0.01406f
C57370 net61 _0261_ 0.57634f
C57371 _1062_/a_381_47# _0160_ 0.12896f
C57372 net23 net25 0
C57373 output56/a_27_47# _0128_ 0
C57374 clknet_1_1__leaf__0465_ net229 0.00466f
C57375 _1020_/a_634_159# net202 0
C57376 net244 hold50/a_391_47# 0
C57377 _0343_ _0424_ 0
C57378 _0179_ acc0.A\[13\] 0.00392f
C57379 _0724_/a_113_297# net208 0
C57380 _0600_/a_253_297# _0219_ 0
C57381 B[9] _0544_/a_245_297# 0
C57382 hold98/a_391_47# net43 0.00357f
C57383 _0603_/a_68_297# _0249_ 0
C57384 _1021_/a_634_159# _0119_ 0.0216f
C57385 _0231_ net213 0
C57386 _0191_ clknet_1_1__leaf__0458_ 0.0237f
C57387 _0081_ _0453_ 0.00148f
C57388 _0558_/a_68_297# input25/a_75_212# 0
C57389 _1017_/a_592_47# _0459_ 0
C57390 _0394_ _0350_ 0
C57391 _0576_/a_109_297# _0380_ 0
C57392 _0147_ _1048_/a_1017_47# 0
C57393 hold55/a_391_47# net23 0.0017f
C57394 _0174_ _0536_/a_149_47# 0.02087f
C57395 _0648_/a_27_297# _0648_/a_277_297# 0.00876f
C57396 _0266_ net247 0
C57397 _0732_/a_80_21# _0368_ 0.09151f
C57398 net168 input12/a_75_212# 0.00208f
C57399 _0510_/a_109_297# net4 0.00625f
C57400 VPWR _0540_/a_240_47# 0.00265f
C57401 hold17/a_285_47# _0979_/a_109_297# 0
C57402 hold17/a_391_47# _0979_/a_27_297# 0.01653f
C57403 clknet_1_1__leaf__0460_ _0698_/a_113_297# 0.0252f
C57404 net115 net94 0.00768f
C57405 _1017_/a_27_47# _0294_ 0
C57406 _0733_/a_222_93# _0361_ 0.00478f
C57407 _1056_/a_891_413# acc0.A\[12\] 0
C57408 net45 _0183_ 0.14505f
C57409 _0477_ net23 0.10324f
C57410 acc0.A\[20\] hold3/a_285_47# 0.00129f
C57411 _1043_/a_193_47# net20 0
C57412 net62 _0988_/a_975_413# 0
C57413 _1011_/a_466_413# _0219_ 0
C57414 _0675_/a_68_297# clknet_1_1__leaf__0461_ 0
C57415 net126 _1041_/a_193_47# 0.00836f
C57416 pp[26] _1026_/a_891_413# 0
C57417 _0467_ _1066_/a_27_47# 0
C57418 _0195_ _0113_ 0
C57419 net132 _1061_/a_975_413# 0
C57420 _0467_ _1068_/a_27_47# 0
C57421 _0217_ _0224_ 0
C57422 _0713_/a_27_47# _0216_ 0
C57423 net157 _0159_ 0
C57424 _0554_/a_68_297# _0175_ 0.10454f
C57425 _0985_/a_27_47# _0985_/a_193_47# 0.96696f
C57426 _0673_/a_253_297# _0288_ 0
C57427 _0411_ net41 0
C57428 _0986_/a_634_159# _0345_ 0
C57429 hold39/a_49_47# _0955_/a_32_297# 0.00133f
C57430 _0368_ clkbuf_1_0__f__0460_/a_110_47# 0
C57431 hold85/a_49_47# net232 0.00252f
C57432 acc0.A\[8\] _0434_ 0.02691f
C57433 _0243_ hold64/a_49_47# 0.04398f
C57434 control0.count\[2\] _1071_/a_1059_315# 0.1282f
C57435 _0642_/a_27_413# _0642_/a_298_297# 0.00498f
C57436 _1055_/a_891_413# _0189_ 0
C57437 net178 _0438_ 0
C57438 hold47/a_49_47# _1050_/a_1059_315# 0.01257f
C57439 _0213_ _0132_ 0.14122f
C57440 VPWR _1067_/a_592_47# 0
C57441 net61 _0509_/a_27_47# 0
C57442 net176 _1022_/a_1059_315# 0
C57443 _0368_ _0250_ 0.00783f
C57444 clknet_0__0460_ _0319_ 0
C57445 _1050_/a_561_413# _0186_ 0.00148f
C57446 _0181_ _0242_ 0
C57447 _0554_/a_150_297# control0.sh 0
C57448 input11/a_75_212# net11 0.10955f
C57449 _0618_/a_215_47# clkbuf_1_0__f__0460_/a_110_47# 0
C57450 _0254_ net235 0
C57451 _0216_ _0612_/a_59_75# 0.02872f
C57452 pp[9] A[10] 0.2001f
C57453 _0582_/a_109_297# net219 0.01148f
C57454 _1019_/a_27_47# _0459_ 0
C57455 _0359_ _1007_/a_891_413# 0
C57456 _0753_/a_297_297# _0753_/a_381_47# 0
C57457 _0753_/a_79_21# _0753_/a_465_47# 0
C57458 net185 _0160_ 0
C57459 hold55/a_49_47# clknet_1_0__leaf__0461_ 0.0336f
C57460 clknet_1_1__leaf__0460_ _0691_/a_68_297# 0
C57461 net154 _0085_ 0
C57462 _0618_/a_215_47# _0250_ 0
C57463 comp0.B\[4\] clknet_1_1__leaf__0463_ 0.11197f
C57464 _0348_ _1030_/a_1017_47# 0
C57465 _0172_ _0548_/a_51_297# 0.1518f
C57466 net180 _0548_/a_512_297# 0
C57467 hold27/a_49_47# clkbuf_0__0464_/a_110_47# 0
C57468 VPWR _1027_/a_466_413# 0.26268f
C57469 net21 net132 0
C57470 _0218_ _0772_/a_297_297# 0.00577f
C57471 B[4] net27 0.00558f
C57472 net45 acc0.A\[15\] 0
C57473 _1003_/a_1059_315# _0381_ 0.00351f
C57474 net17 _0173_ 0.00207f
C57475 _0805_/a_27_47# _0286_ 0.10178f
C57476 _0805_/a_109_47# _0283_ 0
C57477 clknet_1_1__leaf__0462_ hold95/a_285_47# 0
C57478 _0339_ _0568_/a_373_47# 0
C57479 _1031_/a_27_47# _0704_/a_68_297# 0
C57480 _0153_ _0510_/a_27_297# 0
C57481 _0346_ _0291_ 0.15446f
C57482 _0623_/a_109_297# _0186_ 0
C57483 _0869_/a_27_47# net206 0
C57484 _0459_ _0581_/a_373_47# 0
C57485 clk _0970_/a_114_47# 0.00176f
C57486 hold61/a_285_47# net209 0
C57487 _1042_/a_193_47# hold51/a_285_47# 0
C57488 _1042_/a_27_47# hold51/a_391_47# 0
C57489 _0216_ net50 0.33351f
C57490 _0212_ _0132_ 0.01192f
C57491 comp0.B\[13\] comp0.B\[10\] 0
C57492 net240 net107 0.00191f
C57493 _0557_/a_240_47# _1036_/a_1059_315# 0
C57494 _0677_/a_47_47# _0677_/a_377_297# 0.00899f
C57495 _0399_ _1014_/a_634_159# 0
C57496 VPWR _0764_/a_299_297# 0.22004f
C57497 _0422_ _0421_ 0
C57498 _1019_/a_193_47# clknet_1_0__leaf__0461_ 0
C57499 _0559_/a_149_47# net28 0
C57500 _0645_/a_129_47# acc0.A\[13\] 0.00297f
C57501 _1004_/a_891_413# _0378_ 0
C57502 _1004_/a_634_159# _0379_ 0
C57503 acc0.A\[7\] acc0.A\[8\] 0.13085f
C57504 net55 _0730_/a_510_47# 0.00504f
C57505 acc0.A\[8\] _0989_/a_1059_315# 0.03485f
C57506 _0343_ _0755_/a_109_297# 0
C57507 _0188_ net4 0.02834f
C57508 hold54/a_285_47# _0563_/a_240_47# 0
C57509 hold74/a_391_47# acc0.A\[17\] 0.00194f
C57510 pp[17] hold15/a_391_47# 0.02082f
C57511 _0346_ _0991_/a_634_159# 0.00269f
C57512 _0994_/a_27_47# net80 0.26272f
C57513 _0996_/a_1059_315# net6 0
C57514 _0712_/a_561_47# _0340_ 0.01197f
C57515 _0667_/a_113_47# VPWR 0
C57516 _0994_/a_381_47# net246 0
C57517 _0101_ _0352_ 0.00455f
C57518 _0487_ clknet_1_0__leaf__0457_ 0.02769f
C57519 hold88/a_285_47# _0988_/a_1059_315# 0.00319f
C57520 _0544_/a_149_47# _0544_/a_240_47# 0.06872f
C57521 _0544_/a_51_297# _0204_ 0.19811f
C57522 _0811_/a_81_21# hold70/a_49_47# 0.00276f
C57523 clkbuf_1_0__f__0464_/a_110_47# _0186_ 0.00128f
C57524 _0345_ _0737_/a_285_297# 0.00101f
C57525 hold15/a_49_47# VPWR 0.32498f
C57526 hold7/a_49_47# net73 0
C57527 hold74/a_49_47# clkbuf_1_1__f__0461_/a_110_47# 0
C57528 hold30/a_285_47# hold4/a_49_47# 0
C57529 input17/a_75_212# net17 0.10861f
C57530 comp0.B\[15\] control0.reset 0.01761f
C57531 _0730_/a_215_47# _0347_ 0.05723f
C57532 _0313_ _0686_/a_219_297# 0
C57533 hold44/a_285_47# acc0.A\[27\] 0.00186f
C57534 net2 net142 0
C57535 _1034_/a_1059_315# _1034_/a_891_413# 0.31086f
C57536 _1034_/a_193_47# _1034_/a_975_413# 0
C57537 _1034_/a_466_413# _1034_/a_381_47# 0.03733f
C57538 hold6/a_391_47# _0544_/a_51_297# 0.00338f
C57539 _0796_/a_215_47# _0410_ 0.01038f
C57540 _0796_/a_79_21# _0094_ 0.05847f
C57541 _0462_ _0771_/a_215_297# 0
C57542 _0313_ _1008_/a_1059_315# 0
C57543 net162 _1030_/a_975_413# 0
C57544 _1021_/a_381_47# acc0.A\[21\] 0
C57545 _0607_/a_27_297# _0308_ 0
C57546 _0559_/a_245_297# net205 0.00305f
C57547 _0837_/a_81_21# _0433_ 0
C57548 net64 _0434_ 0.01021f
C57549 _0258_ _0268_ 0
C57550 _0464_ _0498_/a_149_47# 0
C57551 clknet_1_0__leaf__0458_ hold2/a_391_47# 0.03229f
C57552 net189 net67 0.25207f
C57553 hold25/a_285_47# net30 0.01422f
C57554 _0982_/a_1017_47# clknet_1_0__leaf__0461_ 0
C57555 _0398_ _0781_/a_150_297# 0
C57556 _0770_/a_79_21# control0.add 0.18903f
C57557 _1051_/a_27_47# clknet_0__0464_ 0
C57558 _0399_ _0781_/a_68_297# 0.00566f
C57559 clkbuf_1_0__f__0465_/a_110_47# clknet_1_1__leaf__0458_ 0.0281f
C57560 _0570_/a_27_297# net197 0.1463f
C57561 _0343_ _0583_/a_373_47# 0
C57562 _0416_ _0285_ 0
C57563 _0229_ _0460_ 0.00159f
C57564 clknet_0__0464_ _1045_/a_634_159# 0
C57565 _0731_/a_299_297# net52 0
C57566 _0226_ clknet_1_0__leaf__0457_ 0.00214f
C57567 _1063_/a_592_47# _0161_ 0
C57568 _0086_ _0988_/a_1059_315# 0
C57569 _0981_/a_109_297# _0468_ 0
C57570 _0483_ _0480_ 0.00748f
C57571 control0.state\[0\] _1068_/a_891_413# 0
C57572 _0842_/a_59_75# _0444_ 0
C57573 _0324_ clkbuf_1_0__f__0462_/a_110_47# 0.02626f
C57574 VPWR _1026_/a_381_47# 0.07615f
C57575 _0454_ acc0.A\[18\] 0.00855f
C57576 _0585_/a_109_297# _0178_ 0
C57577 _0483_ _1072_/a_891_413# 0
C57578 control0.count\[3\] _1072_/a_561_413# 0.00204f
C57579 hold96/a_391_47# net50 0.03967f
C57580 net48 _0764_/a_299_297# 0
C57581 net35 pp[21] 0
C57582 acc0.A\[22\] net46 0.05143f
C57583 _0547_/a_68_297# comp0.B\[8\] 0.18449f
C57584 VPWR _1024_/a_1017_47# 0
C57585 net86 _0181_ 0
C57586 pp[15] _1013_/a_27_47# 0
C57587 hold66/a_285_47# VPWR 0.36105f
C57588 _0559_/a_51_297# _0211_ 0.0013f
C57589 net242 hold95/a_285_47# 0.0102f
C57590 _1018_/a_27_47# _0242_ 0
C57591 _1071_/a_27_47# _0488_ 0.00233f
C57592 clknet_1_0__leaf__0464_ net136 0.21253f
C57593 _0174_ _0177_ 0.06896f
C57594 net18 net19 0.02454f
C57595 hold8/a_49_47# _0347_ 0
C57596 clknet_1_0__leaf__0460_ _1005_/a_891_413# 0.00417f
C57597 hold52/a_391_47# acc0.A\[25\] 0.01293f
C57598 _1017_/a_193_47# _1017_/a_381_47# 0.09799f
C57599 _1017_/a_634_159# _1017_/a_891_413# 0.03684f
C57600 _1017_/a_27_47# _1017_/a_561_413# 0.00163f
C57601 _0487_ _1062_/a_466_413# 0
C57602 pp[18] pp[31] 0.19495f
C57603 _0357_ _0727_/a_109_47# 0.00132f
C57604 _1058_/a_891_413# _0512_/a_27_297# 0
C57605 _1058_/a_1059_315# _0512_/a_109_297# 0
C57606 _0753_/a_79_21# _0234_ 0.00433f
C57607 net178 clknet_1_1__leaf__0465_ 0.03107f
C57608 _1052_/a_193_47# net9 0.04102f
C57609 output65/a_27_47# _0437_ 0
C57610 hold24/a_285_47# net180 0
C57611 _0313_ acc0.A\[23\] 0
C57612 _0473_ _1046_/a_975_413# 0
C57613 _0984_/a_634_159# _0219_ 0
C57614 _1016_/a_27_47# _1060_/a_27_47# 0
C57615 _0216_ _0127_ 0.09505f
C57616 _0179_ _0531_/a_373_47# 0
C57617 _1006_/a_634_159# net52 0
C57618 _1000_/a_466_413# net86 0
C57619 _1000_/a_634_159# _0098_ 0
C57620 _1060_/a_592_47# _0158_ 0
C57621 _0958_/a_27_47# _0161_ 0
C57622 _1056_/a_193_47# hold34/a_285_47# 0.00146f
C57623 _1056_/a_634_159# hold34/a_49_47# 0.00128f
C57624 _1056_/a_27_47# hold34/a_391_47# 0
C57625 _1051_/a_975_413# net11 0
C57626 _0216_ _0399_ 0.013f
C57627 _0129_ _1013_/a_466_413# 0
C57628 control0.count\[1\] _0480_ 0.48586f
C57629 _0346_ _0290_ 0.04559f
C57630 _1072_/a_1017_47# VPWR 0
C57631 net131 net154 0
C57632 hold46/a_285_47# _0200_ 0.04183f
C57633 _0804_/a_297_297# _0804_/a_215_47# 0
C57634 _0804_/a_79_21# _0804_/a_510_47# 0.00844f
C57635 clkbuf_0__0463_/a_110_47# _0465_ 0.00108f
C57636 net160 VPWR 0.42643f
C57637 comp0.B\[10\] comp0.B\[9\] 0.25941f
C57638 _1033_/a_27_47# _1033_/a_193_47# 0.96976f
C57639 _0536_/a_149_47# _1046_/a_193_47# 0
C57640 _0536_/a_240_47# _1046_/a_27_47# 0
C57641 _0536_/a_51_297# _1046_/a_1059_315# 0
C57642 net203 control0.reset 0
C57643 _0320_ _0106_ 0.0023f
C57644 _0985_/a_193_47# _0197_ 0.00206f
C57645 _0520_/a_373_47# clknet_1_0__leaf__0465_ 0.00153f
C57646 _1012_/a_27_47# _1012_/a_193_47# 0.97441f
C57647 acc0.A\[5\] _0989_/a_634_159# 0
C57648 acc0.A\[5\] hold1/a_391_47# 0.00727f
C57649 _0463_ net171 0
C57650 _0293_ _0817_/a_266_47# 0.00417f
C57651 _0165_ _1063_/a_1059_315# 0.00215f
C57652 _0973_/a_109_297# _0161_ 0.01056f
C57653 _0528_/a_299_297# _0527_/a_27_297# 0
C57654 _0528_/a_81_21# _0527_/a_109_297# 0
C57655 net243 hold68/a_285_47# 0
C57656 hold96/a_285_47# net215 0
C57657 hold82/a_285_47# hold82/a_391_47# 0.41909f
C57658 _0195_ net56 0.75257f
C57659 _0401_ _0992_/a_634_159# 0
C57660 net9 net12 0.02416f
C57661 _0102_ _1007_/a_27_47# 0
C57662 _0347_ _1007_/a_1059_315# 0
C57663 _0352_ _1007_/a_193_47# 0
C57664 _1056_/a_27_47# _0510_/a_27_297# 0
C57665 net158 hold36/a_285_47# 0
C57666 clknet_1_0__leaf__0460_ _1006_/a_466_413# 0
C57667 _0363_ _1009_/a_27_47# 0.00221f
C57668 _0963_/a_285_47# _0481_ 0.00308f
C57669 _0216_ _1031_/a_27_47# 0.01309f
C57670 _0195_ _1031_/a_634_159# 0.04558f
C57671 acc0.A\[20\] _1032_/a_193_47# 0
C57672 _0376_ _0755_/a_109_297# 0.00263f
C57673 _0231_ _0618_/a_510_47# 0.005f
C57674 net23 _0352_ 0
C57675 hold70/a_285_47# _0419_ 0
C57676 _0548_/a_149_47# _0545_/a_68_297# 0
C57677 clknet_0__0457_ _0579_/a_109_47# 0.00473f
C57678 VPWR _0650_/a_150_297# 0.00208f
C57679 A[13] _0218_ 0
C57680 net165 _0114_ 0
C57681 _0347_ _0420_ 0
C57682 net164 clkbuf_1_0__f_clk/a_110_47# 0
C57683 clknet_1_1__leaf__0460_ _0361_ 0.00276f
C57684 _1072_/a_466_413# clknet_0_clk 0.01944f
C57685 _1050_/a_1059_315# _1050_/a_891_413# 0.31086f
C57686 _1050_/a_193_47# _1050_/a_975_413# 0
C57687 _1050_/a_466_413# _1050_/a_381_47# 0.03733f
C57688 _0179_ _0990_/a_1059_315# 0
C57689 hold27/a_285_47# _0953_/a_32_297# 0
C57690 hold59/a_49_47# _0454_ 0
C57691 _0990_/a_27_47# _0181_ 0.01099f
C57692 net36 _0854_/a_215_47# 0
C57693 _1041_/a_27_47# _0546_/a_51_297# 0
C57694 _0463_ net24 0
C57695 net232 net17 0.06408f
C57696 hold85/a_391_47# _0946_/a_30_53# 0
C57697 _1014_/a_27_47# _0345_ 0
C57698 net213 _0225_ 0
C57699 _1024_/a_193_47# net50 0.04137f
C57700 _0221_ _1011_/a_975_413# 0
C57701 _0459_ _0347_ 0.05508f
C57702 _0750_/a_27_47# _0227_ 0.00107f
C57703 net44 _0305_ 0.03801f
C57704 hold29/a_49_47# _0122_ 0
C57705 _0428_ _0401_ 0.09031f
C57706 _0427_ _0425_ 0
C57707 _0349_ net44 0
C57708 _0337_ pp[17] 0
C57709 _0338_ acc0.A\[29\] 0
C57710 _0157_ _0219_ 0
C57711 _0465_ _0849_/a_297_297# 0
C57712 _0279_ _0218_ 0.00166f
C57713 _0565_/a_51_297# _0565_/a_240_47# 0.03076f
C57714 _0241_ _0391_ 0.0221f
C57715 _0573_/a_27_47# _0113_ 0
C57716 net116 hold95/a_49_47# 0
C57717 acc0.A\[1\] _0346_ 0.16184f
C57718 _0680_/a_472_297# VPWR 0.01347f
C57719 _0461_ _0769_/a_384_47# 0
C57720 _0595_/a_109_297# acc0.A\[21\] 0.00448f
C57721 _0222_ _0219_ 0.0858f
C57722 _0582_/a_27_297# _0774_/a_68_297# 0
C57723 _0998_/a_891_413# net43 0.01039f
C57724 _0598_/a_79_21# net51 0.03014f
C57725 net58 _0849_/a_79_21# 0
C57726 _0294_ _0245_ 0.05921f
C57727 _1054_/a_193_47# _1052_/a_891_413# 0.00445f
C57728 _1054_/a_634_159# _1052_/a_1059_315# 0.00187f
C57729 hold88/a_391_47# _0186_ 0.04367f
C57730 _0302_ _0297_ 0
C57731 clknet_1_1__leaf__0459_ _0403_ 0.08034f
C57732 _0328_ _0352_ 0
C57733 _0112_ _0208_ 0
C57734 _0982_/a_1059_315# net149 0.00216f
C57735 _0176_ _1040_/a_634_159# 0.02207f
C57736 net1 _0163_ 0
C57737 _1014_/a_27_47# hold2/a_49_47# 0.00167f
C57738 _1039_/a_466_413# _0463_ 0.00729f
C57739 _1039_/a_381_47# clkbuf_0__0463_/a_110_47# 0.00105f
C57740 _0183_ VPWR 5.52683f
C57741 comp0.B\[12\] net196 0.00592f
C57742 net46 _0379_ 0.04061f
C57743 _1056_/a_1059_315# _0179_ 0.06575f
C57744 _0477_ _1062_/a_561_413# 0
C57745 pp[28] _0353_ 0.15374f
C57746 _0833_/a_79_21# net62 0.00189f
C57747 hold46/a_285_47# net193 0.04017f
C57748 net45 _0780_/a_35_297# 0
C57749 _1056_/a_27_47# _0181_ 0
C57750 clknet_1_1__leaf__0461_ _0507_/a_109_47# 0
C57751 _0201_ net184 0
C57752 net205 _1036_/a_27_47# 0
C57753 net46 _0372_ 0.03172f
C57754 net175 clknet_1_1__leaf__0457_ 0.00762f
C57755 _0999_/a_27_47# _0998_/a_891_413# 0
C57756 hold46/a_49_47# _1046_/a_1059_315# 0
C57757 hold92/a_285_47# hold95/a_49_47# 0
C57758 VPWR output63/a_27_47# 0.40221f
C57759 _0533_/a_109_297# _0465_ 0
C57760 hold10/a_391_47# _0180_ 0
C57761 hold10/a_285_47# net8 0
C57762 _1033_/a_891_413# _0208_ 0
C57763 hold67/a_49_47# _0292_ 0
C57764 _0465_ hold71/a_49_47# 0.01435f
C57765 _1012_/a_27_47# clknet_1_1__leaf__0461_ 0.00531f
C57766 _0999_/a_381_47# net85 0.00165f
C57767 _0412_ _0795_/a_299_297# 0
C57768 _0639_/a_109_297# _0218_ 0.002f
C57769 net103 _0115_ 0.14324f
C57770 _0772_/a_510_47# _0391_ 0.00122f
C57771 VPWR _0993_/a_1017_47# 0
C57772 _0629_/a_59_75# acc0.A\[1\] 0
C57773 _0399_ net247 0
C57774 _1016_/a_466_413# net221 0.03246f
C57775 _0752_/a_27_413# _0375_ 0.00294f
C57776 acc0.A\[2\] hold71/a_49_47# 0
C57777 net120 comp0.B\[2\] 0.02135f
C57778 net215 _1024_/a_27_47# 0
C57779 clknet_1_0__leaf__0462_ _1007_/a_1017_47# 0
C57780 _0715_/a_27_47# _0401_ 0.0201f
C57781 _0477_ _0213_ 0
C57782 _0732_/a_80_21# _0732_/a_303_47# 0.01146f
C57783 _0732_/a_209_297# _0732_/a_209_47# 0
C57784 hold18/a_391_47# _0345_ 0.00736f
C57785 _0278_ input5/a_75_212# 0
C57786 _0131_ _0473_ 0
C57787 hold31/a_391_47# acc0.A\[6\] 0.02949f
C57788 VPWR _0542_/a_512_297# 0.00655f
C57789 output66/a_27_47# net2 0.00146f
C57790 clkbuf_1_0__f__0462_/a_110_47# _0347_ 0
C57791 _0323_ _0360_ 0
C57792 _0996_/a_27_47# net42 0
C57793 clknet_0__0463_ _0564_/a_150_297# 0
C57794 hold91/a_49_47# _0669_/a_29_53# 0
C57795 _1043_/a_27_47# net195 0
C57796 _1043_/a_634_159# _0203_ 0.00315f
C57797 clkbuf_1_0__f__0458_/a_110_47# hold75/a_285_47# 0.02258f
C57798 _0186_ _0823_/a_109_297# 0
C57799 net220 _0219_ 0
C57800 _0212_ net25 0.36001f
C57801 _1033_/a_1059_315# net17 0.03182f
C57802 _0563_/a_51_297# _0560_/a_68_297# 0
C57803 _1016_/a_891_413# _0459_ 0.00521f
C57804 _0648_/a_277_297# _0280_ 0
C57805 _0500_/a_27_47# net157 0
C57806 _0183_ net48 0.02794f
C57807 clkbuf_1_1__f__0463_/a_110_47# control0.sh 0
C57808 hold17/a_391_47# _0169_ 0.01467f
C57809 control0.count\[2\] net164 0.18403f
C57810 _0234_ clkbuf_1_0__f__0460_/a_110_47# 0
C57811 _0732_/a_80_21# clknet_0__0460_ 0
C57812 _0443_ _0428_ 0
C57813 VPWR acc0.A\[15\] 2.67842f
C57814 _0206_ _0543_/a_68_297# 0
C57815 _1052_/a_27_47# _0522_/a_27_297# 0
C57816 _0195_ _0345_ 0.43276f
C57817 _1002_/a_561_413# clknet_1_0__leaf__0460_ 0
C57818 _0234_ _0250_ 0
C57819 net92 _0345_ 0
C57820 _0221_ _0334_ 0.18466f
C57821 _0416_ _0218_ 0.02534f
C57822 acc0.A\[12\] _0286_ 0.02927f
C57823 net188 acc0.A\[11\] 0.39406f
C57824 _0518_/a_27_297# net15 0.19131f
C57825 net10 _0541_/a_150_297# 0
C57826 _0614_/a_111_297# _0246_ 0
C57827 hold86/a_285_47# _0446_ 0.0516f
C57828 _0856_/a_510_47# _0345_ 0.00153f
C57829 _0712_/a_79_21# _0216_ 0
C57830 _0712_/a_381_47# _0195_ 0
C57831 _0985_/a_634_159# _0985_/a_1017_47# 0
C57832 _0985_/a_466_413# _0985_/a_592_47# 0.00553f
C57833 hold100/a_49_47# acc0.A\[14\] 0.28434f
C57834 hold39/a_391_47# comp0.B\[6\] 0.00628f
C57835 clkbuf_1_0__f__0463_/a_110_47# _1040_/a_27_47# 0.00586f
C57836 _0563_/a_240_47# _0562_/a_68_297# 0
C57837 clknet_1_1__leaf__0458_ _0824_/a_145_75# 0
C57838 _0326_ _1007_/a_634_159# 0
C57839 _0998_/a_381_47# _0181_ 0
C57840 _1020_/a_27_47# net88 0
C57841 _1018_/a_466_413# _1018_/a_561_413# 0.00772f
C57842 _1018_/a_634_159# _1018_/a_975_413# 0
C57843 _0297_ net6 0.0361f
C57844 net36 _1014_/a_466_413# 0
C57845 hold85/a_391_47# _0967_/a_109_93# 0
C57846 hold85/a_285_47# _0967_/a_215_297# 0.00115f
C57847 clkbuf_1_0__f__0460_/a_110_47# clknet_0__0460_ 0.31131f
C57848 hold19/a_391_47# _1016_/a_27_47# 0
C57849 hold19/a_285_47# _1016_/a_193_47# 0.00369f
C57850 hold19/a_49_47# _1016_/a_634_159# 0.00169f
C57851 hold11/a_285_47# _0464_ 0.00198f
C57852 _0390_ _0183_ 0
C57853 comp0.B\[14\] _1046_/a_1059_315# 0.08741f
C57854 _0670_/a_79_21# _0219_ 0
C57855 _0195_ hold2/a_49_47# 0
C57856 _0982_/a_27_47# _0982_/a_561_413# 0.0027f
C57857 _0982_/a_634_159# _0982_/a_891_413# 0.03684f
C57858 _0982_/a_193_47# _0982_/a_381_47# 0.09503f
C57859 _0592_/a_150_297# clknet_1_0__leaf__0460_ 0
C57860 _1011_/a_193_47# clknet_1_1__leaf__0462_ 0
C57861 _1049_/a_634_159# _1049_/a_1059_315# 0
C57862 _1049_/a_27_47# _1049_/a_381_47# 0.06222f
C57863 _1049_/a_193_47# _1049_/a_891_413# 0.19489f
C57864 _0343_ _1018_/a_891_413# 0.00667f
C57865 _0725_/a_303_47# _0339_ 0
C57866 _0324_ net51 0
C57867 _0250_ clknet_0__0460_ 0.03913f
C57868 _0284_ _0347_ 0
C57869 _0983_/a_381_47# acc0.A\[15\] 0
C57870 _0430_ _0258_ 0
C57871 net148 _0522_/a_109_47# 0
C57872 _0659_/a_68_297# net47 0
C57873 output37/a_27_47# A[11] 0.05117f
C57874 _0753_/a_561_47# _0231_ 0.00969f
C57875 _0666_/a_113_47# _0297_ 0
C57876 _0465_ _0529_/a_109_297# 0
C57877 _0289_ _0657_/a_109_297# 0.01181f
C57878 _0399_ _0841_/a_79_21# 0.19678f
C57879 comp0.B\[5\] net28 0.29896f
C57880 net180 _0138_ 0.30165f
C57881 _0412_ net6 0
C57882 _1019_/a_193_47# _0218_ 0
C57883 hold56/a_285_47# _0133_ 0
C57884 VPWR net156 0.2999f
C57885 hold98/a_391_47# net40 0
C57886 hold98/a_49_47# net245 0.00115f
C57887 hold79/a_391_47# net226 0.15711f
C57888 _0369_ _0304_ 0
C57889 _0258_ acc0.A\[5\] 0
C57890 hold16/a_49_47# _0195_ 0.0131f
C57891 _0268_ net72 0
C57892 acc0.A\[27\] _0219_ 0.12958f
C57893 _1066_/a_634_159# _1066_/a_1059_315# 0
C57894 _1066_/a_27_47# _1066_/a_381_47# 0.06222f
C57895 _1066_/a_193_47# _1066_/a_891_413# 0.19497f
C57896 hold37/a_391_47# _1050_/a_193_47# 0
C57897 net56 _1010_/a_891_413# 0.00329f
C57898 pp[10] _0512_/a_109_297# 0
C57899 net58 _0529_/a_27_297# 0
C57900 acc0.A\[14\] _0410_ 0.04497f
C57901 net1 _1066_/a_27_47# 0
C57902 _0098_ _0242_ 0
C57903 _0101_ _0237_ 0.02885f
C57904 net45 _0999_/a_381_47# 0.00271f
C57905 VPWR _1052_/a_561_413# 0.00213f
C57906 _0538_/a_51_297# _1042_/a_1059_315# 0
C57907 _0852_/a_35_297# _0345_ 0.0055f
C57908 _1031_/a_891_413# acc0.A\[30\] 0
C57909 _1023_/a_466_413# _1022_/a_1059_315# 0
C57910 _0476_ clkbuf_0_clk/a_110_47# 0
C57911 clkload3/a_268_47# clkload3/Y 0.00587f
C57912 _1068_/a_634_159# _1068_/a_1059_315# 0
C57913 _1068_/a_27_47# _1068_/a_381_47# 0.05658f
C57914 _1068_/a_193_47# _1068_/a_891_413# 0.19226f
C57915 net44 _0181_ 0.00351f
C57916 _1030_/a_27_47# _1030_/a_193_47# 0.9705f
C57917 _0179_ VPWR 5.39517f
C57918 acc0.A\[14\] _0450_ 0.02146f
C57919 _0557_/a_512_297# comp0.B\[4\] 0.00116f
C57920 net71 _0844_/a_79_21# 0
C57921 net237 _0360_ 0.08002f
C57922 _0487_ _1063_/a_1017_47# 0
C57923 VPWR _0971_/a_384_47# 0
C57924 _0286_ _0650_/a_68_297# 0
C57925 _0283_ _0650_/a_150_297# 0
C57926 VPWR B[14] 0.2463f
C57927 _1034_/a_27_47# clknet_1_1__leaf_clk 0
C57928 net205 comp0.B\[3\] 0.00297f
C57929 pp[29] _0219_ 0
C57930 output67/a_27_47# net3 0.05725f
C57931 VPWR hold40/a_285_47# 0.28265f
C57932 _1032_/a_891_413# net23 0
C57933 _0312_ _1009_/a_193_47# 0
C57934 _0313_ clknet_1_1__leaf__0462_ 0.0012f
C57935 _0449_ _0219_ 0.04318f
C57936 _0346_ net77 0
C57937 _1035_/a_193_47# clknet_1_1__leaf__0463_ 0.01124f
C57938 _0232_ acc0.A\[23\] 0
C57939 _0992_/a_193_47# hold70/a_285_47# 0.00171f
C57940 _0992_/a_27_47# hold70/a_391_47# 0
C57941 _0344_ _0342_ 0.29154f
C57942 comp0.B\[10\] hold5/a_285_47# 0.09469f
C57943 hold53/a_49_47# _0123_ 0.2937f
C57944 _0183_ clknet_1_0__leaf__0459_ 1.48425f
C57945 _0217_ net87 0.10366f
C57946 _0519_/a_299_297# _0252_ 0.06522f
C57947 _0108_ _0352_ 0
C57948 hold47/a_285_47# _1051_/a_27_47# 0
C57949 hold47/a_49_47# _1051_/a_193_47# 0
C57950 _0269_ _0261_ 0.16855f
C57951 _1051_/a_1059_315# _0186_ 0.00448f
C57952 _1034_/a_466_413# comp0.B\[2\] 0.03589f
C57953 _0155_ acc0.A\[11\] 0.02636f
C57954 output65/a_27_47# _0252_ 0
C57955 pp[7] _0989_/a_193_47# 0
C57956 acc0.A\[27\] _1008_/a_634_159# 0.01768f
C57957 VPWR _0513_/a_81_21# 0.20063f
C57958 hold98/a_49_47# net45 0
C57959 _0979_/a_373_47# _0466_ 0
C57960 hold64/a_285_47# _0399_ 0
C57961 _0110_ _0219_ 0
C57962 clknet_0__0464_ _1044_/a_193_47# 0
C57963 _1072_/a_193_47# _0466_ 0.00175f
C57964 net43 _0793_/a_240_47# 0.03887f
C57965 _0816_/a_150_297# _0426_ 0
C57966 net45 clkload3/a_110_47# 0
C57967 hold89/a_285_47# clkbuf_0_clk/a_110_47# 0
C57968 _0958_/a_109_47# _0487_ 0
C57969 _0225_ _0618_/a_510_47# 0.00141f
C57970 net197 _0126_ 0.23385f
C57971 clknet_0__0464_ net131 0.18652f
C57972 _0534_/a_299_297# _1047_/a_891_413# 0
C57973 _0481_ net226 0.20007f
C57974 _0346_ _1006_/a_1059_315# 0.05593f
C57975 _0346_ _0656_/a_59_75# 0
C57976 _0247_ _0611_/a_68_297# 0
C57977 hold57/a_285_47# _0474_ 0
C57978 _0267_ _0347_ 0
C57979 _0369_ _0619_/a_150_297# 0
C57980 net34 _0166_ 0
C57981 net126 comp0.B\[10\] 0
C57982 _0756_/a_377_297# net50 0.00156f
C57983 VPWR acc0.A\[26\] 0.86428f
C57984 _0293_ _0181_ 0.00602f
C57985 net168 hold21/a_49_47# 0
C57986 _0179_ input4/a_75_212# 0
C57987 pp[30] _1031_/a_561_413# 0
C57988 _1058_/a_1059_315# _0189_ 0
C57989 _0346_ _0986_/a_1059_315# 0
C57990 _1032_/a_466_413# clknet_1_0__leaf__0461_ 0.02082f
C57991 _0686_/a_219_297# _0321_ 0
C57992 net144 input3/a_75_212# 0
C57993 _0258_ _0443_ 0.02848f
C57994 _0973_/a_109_47# _0487_ 0.00269f
C57995 _0805_/a_27_47# net79 0
C57996 net104 acc0.A\[19\] 0
C57997 _0183_ _0453_ 0
C57998 _1071_/a_1017_47# _0466_ 0
C57999 _0343_ _0998_/a_193_47# 0.00384f
C58000 _1021_/a_891_413# _0352_ 0.00272f
C58001 _1008_/a_1059_315# _0321_ 0
C58002 net54 _0317_ 0
C58003 _0645_/a_47_47# _0996_/a_193_47# 0
C58004 _0476_ _1062_/a_381_47# 0
C58005 _1017_/a_891_413# net103 0
C58006 _0487_ _0160_ 0
C58007 net106 net23 0.02435f
C58008 _0602_/a_113_47# _0232_ 0
C58009 acc0.A\[12\] _0672_/a_79_21# 0.07921f
C58010 _0642_/a_27_413# clkbuf_1_0__f__0465_/a_110_47# 0
C58011 _1017_/a_193_47# _1016_/a_634_159# 0
C58012 _1017_/a_634_159# _1016_/a_193_47# 0.00136f
C58013 _1017_/a_466_413# _1016_/a_27_47# 0.0047f
C58014 _1017_/a_27_47# _1016_/a_466_413# 0
C58015 _0343_ _0376_ 0.05506f
C58016 _0233_ _0375_ 0.11311f
C58017 _0661_/a_27_297# _0661_/a_109_297# 0.00695f
C58018 clknet_1_0__leaf__0459_ acc0.A\[15\] 0.01641f
C58019 acc0.A\[8\] _0988_/a_466_413# 0
C58020 _0998_/a_27_47# acc0.A\[17\] 0
C58021 _0181_ _0566_/a_27_47# 0.01599f
C58022 net70 _0219_ 0
C58023 _0201_ _0176_ 0.00696f
C58024 _0253_ clkbuf_1_1__f__0458_/a_110_47# 0.00673f
C58025 net92 net52 0
C58026 net86 _0098_ 0.03196f
C58027 _0101_ _1005_/a_27_47# 0
C58028 _0477_ _0161_ 0.02186f
C58029 _0565_/a_51_297# _0171_ 0
C58030 input4/a_75_212# _0513_/a_81_21# 0
C58031 clkload0/a_27_47# _1071_/a_1059_315# 0.00502f
C58032 _0733_/a_222_93# VPWR 0.0829f
C58033 _1067_/a_193_47# _1065_/a_193_47# 0.00249f
C58034 _0837_/a_81_21# _0835_/a_78_199# 0
C58035 _0465_ _0264_ 0.01434f
C58036 _0298_ _0797_/a_27_413# 0
C58037 _0404_ _0797_/a_207_413# 0
C58038 _0521_/a_299_297# _0151_ 0.0681f
C58039 _1033_/a_466_413# _1033_/a_592_47# 0.00553f
C58040 _1033_/a_634_159# _1033_/a_1017_47# 0
C58041 _0457_ comp0.B\[15\] 0.0029f
C58042 _0286_ net42 0
C58043 hold3/a_391_47# net51 0
C58044 _0283_ acc0.A\[15\] 0
C58045 _0259_ _0291_ 0.07834f
C58046 _0221_ _0724_/a_113_297# 0.05024f
C58047 _0347_ net51 0
C58048 net194 hold37/a_391_47# 0.00959f
C58049 _1012_/a_466_413# _1012_/a_592_47# 0.00553f
C58050 _1012_/a_634_159# _1012_/a_1017_47# 0
C58051 _1039_/a_891_413# _0176_ 0.03051f
C58052 VPWR _0780_/a_35_297# 0.22461f
C58053 _0130_ _1033_/a_27_47# 0
C58054 _0216_ _0327_ 0
C58055 clknet_1_1__leaf__0460_ _0726_/a_51_297# 0.00157f
C58056 _0846_/a_149_47# _0345_ 0.00154f
C58057 _0985_/a_27_47# _0636_/a_59_75# 0
C58058 _0529_/a_27_297# _0262_ 0
C58059 _0530_/a_81_21# _0147_ 0.11488f
C58060 hold79/a_285_47# _0162_ 0
C58061 _1056_/a_27_47# _0187_ 0
C58062 pp[1] A[9] 0
C58063 net76 _0988_/a_891_413# 0
C58064 _0285_ net246 0
C58065 _0343_ A[14] 0
C58066 _0805_/a_109_47# _0345_ 0
C58067 _0243_ _1000_/a_27_47# 0
C58068 hold27/a_285_47# _0174_ 0
C58069 clknet_1_0__leaf__0458_ _0853_/a_150_297# 0
C58070 _1009_/a_634_159# _0219_ 0.04517f
C58071 hold86/a_285_47# net61 0.00319f
C58072 _0220_ hold95/a_49_47# 0
C58073 clknet_1_0__leaf__0457_ _0350_ 0.09408f
C58074 net44 _0677_/a_377_297# 0.0058f
C58075 _1050_/a_466_413# acc0.A\[4\] 0.03097f
C58076 net15 _0987_/a_27_47# 0
C58077 _0453_ acc0.A\[15\] 0
C58078 clknet_1_1__leaf__0464_ hold51/a_285_47# 0
C58079 _0348_ acc0.A\[29\] 0
C58080 net35 _0237_ 0
C58081 _1055_/a_1059_315# acc0.A\[9\] 0.10942f
C58082 _1041_/a_1059_315# _0205_ 0.00362f
C58083 _1041_/a_193_47# net32 0
C58084 _1041_/a_634_159# net152 0
C58085 comp0.B\[2\] net118 0
C58086 hold88/a_391_47# net62 0.03271f
C58087 _0162_ net17 0
C58088 clknet_0_clk _0951_/a_209_311# 0
C58089 clkbuf_1_0__f__0465_/a_110_47# _0218_ 0.04132f
C58090 _1033_/a_1059_315# _0165_ 0
C58091 _0350_ _0988_/a_1059_315# 0
C58092 net36 net7 0
C58093 VPWR _0441_ 0.3725f
C58094 hold26/a_285_47# _0138_ 0.00385f
C58095 _0508_/a_299_297# _0508_/a_384_47# 0
C58096 _0465_ net170 0
C58097 clkbuf_1_0__f__0463_/a_110_47# net171 0.00181f
C58098 comp0.B\[4\] input28/a_75_212# 0
C58099 VPWR _0544_/a_51_297# 0.44292f
C58100 net158 hold26/a_49_47# 0
C58101 _0476_ net185 0.12698f
C58102 _0983_/a_27_47# _1018_/a_634_159# 0
C58103 hold96/a_49_47# net52 0.01744f
C58104 VPWR _1034_/a_193_47# 0.28439f
C58105 _0204_ _1043_/a_27_47# 0
C58106 _0544_/a_240_47# _1043_/a_466_413# 0
C58107 _0960_/a_181_47# VPWR 0
C58108 _1004_/a_634_159# _0575_/a_27_297# 0
C58109 _1004_/a_193_47# _0575_/a_109_297# 0
C58110 hold34/a_49_47# hold35/a_49_47# 0.00686f
C58111 _0369_ clknet_1_0__leaf__0460_ 0.06191f
C58112 acc0.A\[2\] net170 0.00784f
C58113 _1017_/a_193_47# _0116_ 0
C58114 _0465_ _0845_/a_109_297# 0
C58115 clkload3/Y clkbuf_1_1__f__0461_/a_110_47# 0.00248f
C58116 hold65/a_285_47# _0435_ 0
C58117 hold65/a_49_47# _0436_ 0
C58118 clkbuf_1_0__f__0458_/a_110_47# _0345_ 0.03368f
C58119 _0553_/a_51_297# _0463_ 0
C58120 _0179_ _1054_/a_1017_47# 0
C58121 net21 _1044_/a_1017_47# 0
C58122 _0998_/a_27_47# _0998_/a_634_159# 0.13601f
C58123 _0956_/a_32_297# _0208_ 0.05665f
C58124 net64 _0988_/a_466_413# 0.02313f
C58125 _1059_/a_27_47# _0459_ 0.01257f
C58126 _1031_/a_561_413# _0339_ 0.0017f
C58127 _1031_/a_975_413# _0338_ 0
C58128 hold96/a_285_47# clknet_1_0__leaf__0460_ 0
C58129 hold58/a_285_47# comp0.B\[4\] 0.10313f
C58130 clknet_1_1__leaf__0459_ acc0.A\[13\] 0.02427f
C58131 net214 _0369_ 0.38978f
C58132 clkbuf_1_1__f__0463_/a_110_47# _0955_/a_32_297# 0
C58133 _0179_ _0283_ 0
C58134 _0750_/a_27_47# _0352_ 0
C58135 _0734_/a_377_297# _0370_ 0
C58136 acc0.A\[29\] _0332_ 0.00836f
C58137 _0432_ _0640_/a_465_297# 0
C58138 _0183_ _0113_ 0
C58139 _1001_/a_1059_315# _0350_ 0.02404f
C58140 _1046_/a_634_159# _1046_/a_592_47# 0
C58141 net44 _1012_/a_193_47# 0.00182f
C58142 _0475_ comp0.B\[15\] 0.00339f
C58143 _1019_/a_193_47# _0099_ 0
C58144 acc0.A\[21\] hold3/a_49_47# 0.31354f
C58145 _0557_/a_149_47# _0549_/a_68_297# 0
C58146 net203 _0457_ 0
C58147 net54 net197 0.06805f
C58148 _1056_/a_193_47# _0153_ 0.00188f
C58149 clkbuf_1_1__f__0458_/a_110_47# net74 0
C58150 clknet_1_0__leaf__0464_ _0533_/a_27_297# 0
C58151 clknet_1_0__leaf__0463_ input29/a_75_212# 0.01007f
C58152 _1032_/a_592_47# clknet_1_0__leaf__0457_ 0
C58153 _0458_ _0446_ 0.05406f
C58154 net166 net221 0.02255f
C58155 _1016_/a_592_47# _0115_ 0.00121f
C58156 _0753_/a_561_47# _0225_ 0
C58157 net154 _0525_/a_81_21# 0.05916f
C58158 _1051_/a_891_413# _1050_/a_193_47# 0
C58159 _1051_/a_466_413# _1050_/a_466_413# 0.01154f
C58160 _1051_/a_193_47# _1050_/a_891_413# 0
C58161 _1039_/a_466_413# clkbuf_1_0__f__0463_/a_110_47# 0.00169f
C58162 _0985_/a_891_413# net175 0
C58163 VPWR _0141_ 0.41206f
C58164 _0748_/a_81_21# _0370_ 0
C58165 _0982_/a_634_159# clkbuf_0__0457_/a_110_47# 0
C58166 _0996_/a_1017_47# acc0.A\[15\] 0
C58167 hold91/a_391_47# _0301_ 0
C58168 _0556_/a_68_297# comp0.B\[4\] 0.18776f
C58169 hold34/a_49_47# A[9] 0.00388f
C58170 net175 _1049_/a_634_159# 0
C58171 hold87/a_49_47# net47 0.02582f
C58172 acc0.A\[12\] _1057_/a_1017_47# 0.00126f
C58173 _0272_ _0840_/a_150_297# 0
C58174 _0998_/a_381_47# clknet_1_1__leaf__0461_ 0
C58175 _0259_ _0290_ 0.04794f
C58176 _0661_/a_277_297# _0426_ 0
C58177 _0576_/a_27_297# _0216_ 0
C58178 _0775_/a_79_21# _0352_ 0.16778f
C58179 clkload1/Y net248 0.0524f
C58180 _0775_/a_510_47# _0347_ 0.00122f
C58181 _0627_/a_215_53# _0399_ 0
C58182 _0457_ _1032_/a_561_413# 0
C58183 _1041_/a_193_47# net10 0
C58184 control0.state\[0\] clkbuf_1_0__f_clk/a_110_47# 0
C58185 clknet_1_1__leaf__0459_ net85 0.09664f
C58186 pp[30] _0129_ 0.00461f
C58187 net59 net163 0
C58188 acc0.A\[8\] _0186_ 0.45691f
C58189 _0707_/a_75_199# hold61/a_391_47# 0
C58190 net90 net52 0.19664f
C58191 _0758_/a_79_21# _0758_/a_297_297# 0.01735f
C58192 _0179_ hold35/a_391_47# 0
C58193 VPWR _0999_/a_381_47# 0.07033f
C58194 hold27/a_391_47# _0536_/a_240_47# 0
C58195 _1052_/a_891_413# acc0.A\[6\] 0.05455f
C58196 _1052_/a_27_47# _0193_ 0
C58197 _0752_/a_27_413# VPWR 0.22575f
C58198 _0614_/a_183_297# _0352_ 0
C58199 _0581_/a_27_297# net219 0.07519f
C58200 _0990_/a_27_47# _0990_/a_193_47# 0.96574f
C58201 _0230_ _0227_ 0.19431f
C58202 hold22/a_285_47# A[8] 0
C58203 _0789_/a_75_199# acc0.A\[15\] 0
C58204 _0534_/a_81_21# net149 0.06946f
C58205 net15 _0191_ 0.5f
C58206 net10 net11 0
C58207 _0697_/a_217_297# clkbuf_1_1__f__0460_/a_110_47# 0
C58208 _1039_/a_592_47# net8 0
C58209 _0985_/a_592_47# _0083_ 0
C58210 _0984_/a_634_159# net58 0
C58211 _0501_/a_27_47# _0465_ 0.00367f
C58212 _0672_/a_79_21# net42 0.05288f
C58213 _0850_/a_68_297# _0350_ 0.01375f
C58214 net150 _0605_/a_109_297# 0
C58215 _0343_ _0990_/a_381_47# 0.01283f
C58216 _0985_/a_466_413# acc0.A\[3\] 0.00319f
C58217 _0260_ _0219_ 0
C58218 _0346_ _1014_/a_634_159# 0.00365f
C58219 _0970_/a_285_47# _0162_ 0.00799f
C58220 _0484_ _0485_ 0.3093f
C58221 _0343_ _0793_/a_51_297# 0.02295f
C58222 net44 clknet_1_1__leaf__0461_ 0.02681f
C58223 _1053_/a_1059_315# _0191_ 0.00113f
C58224 _0982_/a_1059_315# _0080_ 0
C58225 _0982_/a_891_413# net68 0
C58226 VPWR hold83/a_49_47# 0.27316f
C58227 _0343_ clkbuf_1_0__f__0459_/a_110_47# 0.02966f
C58228 hold88/a_285_47# net235 0.00885f
C58229 _1049_/a_27_47# acc0.A\[3\] 0
C58230 _1049_/a_466_413# _0147_ 0.02084f
C58231 _1049_/a_1059_315# net135 0
C58232 hold25/a_49_47# _1040_/a_193_47# 0
C58233 hold25/a_285_47# _1040_/a_27_47# 0
C58234 _1011_/a_27_47# hold80/a_285_47# 0
C58235 _1011_/a_193_47# hold80/a_49_47# 0
C58236 net203 _0475_ 0.08996f
C58237 net245 clknet_1_1__leaf__0459_ 0.02162f
C58238 _0747_/a_215_47# net216 0.04611f
C58239 _0229_ _0373_ 0.10789f
C58240 _0598_/a_297_47# hold3/a_49_47# 0.03824f
C58241 hold96/a_285_47# _0576_/a_109_297# 0
C58242 _0606_/a_215_297# _0606_/a_465_297# 0.00827f
C58243 _0473_ _1044_/a_891_413# 0
C58244 _0381_ net159 0
C58245 VPWR _0530_/a_384_47# 0
C58246 _1070_/a_634_159# _1070_/a_1059_315# 0
C58247 _1070_/a_27_47# _1070_/a_381_47# 0.06222f
C58248 _1070_/a_193_47# _1070_/a_891_413# 0.19685f
C58249 _1053_/a_193_47# _1053_/a_592_47# 0.00135f
C58250 _1053_/a_466_413# _1053_/a_561_413# 0.00772f
C58251 _1053_/a_634_159# _1053_/a_975_413# 0
C58252 hold42/a_285_47# acc0.A\[10\] 0
C58253 output44/a_27_47# _1030_/a_1059_315# 0.00107f
C58254 net44 _1030_/a_193_47# 0.25803f
C58255 _0382_ _0460_ 0.00242f
C58256 hold98/a_49_47# VPWR 0.32619f
C58257 _0647_/a_47_47# _0647_/a_285_47# 0.01755f
C58258 _0575_/a_109_297# net199 0.01296f
C58259 _0578_/a_373_47# net23 0
C58260 clknet_1_0__leaf__0465_ _1050_/a_1059_315# 0.00712f
C58261 _1015_/a_193_47# net118 0
C58262 _0532_/a_81_21# _0465_ 0.00516f
C58263 net45 _0998_/a_466_413# 0.00401f
C58264 _0198_ _1061_/a_193_47# 0.00124f
C58265 _1032_/a_193_47# _0208_ 0
C58266 _1032_/a_1059_315# _0173_ 0
C58267 acc0.A\[22\] _1023_/a_193_47# 0
C58268 _0996_/a_381_47# _0181_ 0
C58269 _0294_ _0326_ 0
C58270 hold43/a_285_47# _0195_ 0.00189f
C58271 _1066_/a_1059_315# clknet_1_1__leaf_clk 0
C58272 _1066_/a_27_47# control0.sh 0.01172f
C58273 _0179_ _0523_/a_81_21# 0.01138f
C58274 clkload3/a_110_47# VPWR 0
C58275 hold75/a_285_47# acc0.A\[15\] 0.00781f
C58276 _0314_ _1007_/a_1059_315# 0.04445f
C58277 _0991_/a_381_47# net47 0
C58278 _1037_/a_891_413# _0176_ 0
C58279 _0378_ _0754_/a_51_297# 0
C58280 _0082_ _0261_ 0
C58281 _1034_/a_381_47# _0175_ 0.017f
C58282 _0752_/a_27_413# net48 0.00398f
C58283 _0179_ net182 0.08669f
C58284 hold32/a_391_47# clknet_1_1__leaf__0465_ 0.00876f
C58285 hold10/a_285_47# _0492_/a_27_47# 0
C58286 _0309_ _0777_/a_129_47# 0.00159f
C58287 acc0.A\[2\] _0532_/a_81_21# 0
C58288 net109 _1022_/a_891_413# 0.00263f
C58289 net177 _1022_/a_1059_315# 0.04013f
C58290 net235 _0086_ 0.0083f
C58291 _0311_ _0462_ 0.03694f
C58292 _1068_/a_466_413# _0166_ 0.00167f
C58293 _1030_/a_466_413# _1030_/a_592_47# 0.00553f
C58294 _1030_/a_634_159# _1030_/a_1017_47# 0
C58295 clkbuf_1_1__f__0464_/a_110_47# _1044_/a_891_413# 0.01528f
C58296 VPWR input13/a_75_212# 0.27221f
C58297 hold5/a_391_47# net153 0
C58298 _0134_ comp0.B\[4\] 0
C58299 clknet_1_1__leaf__0460_ VPWR 4.07772f
C58300 _0218_ net246 0.08097f
C58301 net188 A[12] 0
C58302 _0244_ clknet_1_0__leaf__0457_ 0
C58303 clknet_1_0__leaf__0462_ _0758_/a_297_297# 0
C58304 _0256_ _0271_ 0.24367f
C58305 _0376_ _0224_ 0
C58306 _0443_ net72 0.02645f
C58307 _0330_ _0354_ 0
C58308 hold27/a_49_47# _1046_/a_634_159# 0
C58309 hold27/a_391_47# _1046_/a_27_47# 0
C58310 hold27/a_285_47# _1046_/a_193_47# 0
C58311 _1014_/a_1059_315# hold60/a_285_47# 0.00319f
C58312 net64 _0186_ 0.02763f
C58313 acc0.A\[12\] net79 0
C58314 acc0.A\[14\] _0637_/a_56_297# 0.04353f
C58315 _0764_/a_299_297# _0345_ 0.00339f
C58316 _1035_/a_1017_47# net122 0
C58317 _1056_/a_27_47# _1056_/a_193_47# 0.96639f
C58318 _0992_/a_975_413# net37 0
C58319 _0415_ _0347_ 0.14775f
C58320 _1032_/a_27_47# net17 0.00919f
C58321 net122 net23 0
C58322 _0671_/a_113_297# _0671_/a_199_47# 0
C58323 _0243_ acc0.A\[19\] 1.08538f
C58324 control0.state\[0\] control0.count\[2\] 0
C58325 _1015_/a_1017_47# _0181_ 0.00134f
C58326 _0320_ _0360_ 0
C58327 _0987_/a_466_413# _0987_/a_381_47# 0.03733f
C58328 _0987_/a_193_47# _0987_/a_975_413# 0
C58329 _0987_/a_1059_315# _0987_/a_891_413# 0.31086f
C58330 _0721_/a_27_47# _0208_ 0.22735f
C58331 net194 _1051_/a_891_413# 0
C58332 _0355_ _0333_ 0.05047f
C58333 _0579_/a_373_47# _0183_ 0
C58334 _0604_/a_113_47# _0462_ 0
C58335 net45 clknet_1_1__leaf__0459_ 0.07688f
C58336 _0855_/a_81_21# _0855_/a_299_297# 0.08213f
C58337 _0180_ _1047_/a_193_47# 0
C58338 acc0.A\[1\] _1047_/a_466_413# 0
C58339 _0182_ _1047_/a_634_159# 0.00576f
C58340 _0608_/a_109_297# _0306_ 0
C58341 _0608_/a_27_47# _0308_ 0.05044f
C58342 hold15/a_49_47# _0345_ 0
C58343 acc0.A\[20\] _0765_/a_510_47# 0.00608f
C58344 acc0.A\[27\] net94 0.00441f
C58345 _0992_/a_1017_47# net67 0
C58346 _1000_/a_1017_47# VPWR 0
C58347 _1004_/a_193_47# _1004_/a_891_413# 0.19489f
C58348 _1004_/a_27_47# _1004_/a_381_47# 0.06222f
C58349 _1004_/a_634_159# _1004_/a_1059_315# 0
C58350 _0729_/a_68_297# net57 0.00295f
C58351 _0129_ _0339_ 0.04624f
C58352 net69 _0181_ 0
C58353 _1027_/a_193_47# _1008_/a_27_47# 0
C58354 _1027_/a_27_47# _1008_/a_193_47# 0
C58355 _0557_/a_51_297# _1035_/a_466_413# 0
C58356 net157 _1049_/a_27_47# 0.00496f
C58357 _0788_/a_68_297# _0399_ 0.01961f
C58358 _0369_ _0434_ 0.06236f
C58359 hold15/a_285_47# _0712_/a_297_297# 0
C58360 _0967_/a_215_297# _0477_ 0.00197f
C58361 rst _1064_/a_193_47# 0
C58362 _0493_/a_27_47# _0171_ 0.03743f
C58363 _0216_ _0346_ 0.04253f
C58364 clknet_1_1__leaf__0462_ _0321_ 0
C58365 net180 net22 0
C58366 _0603_/a_68_297# _0462_ 0.00242f
C58367 _1029_/a_1059_315# _1029_/a_891_413# 0.31086f
C58368 _1029_/a_193_47# _1029_/a_975_413# 0
C58369 _1029_/a_466_413# _1029_/a_381_47# 0.03733f
C58370 hold75/a_285_47# _0179_ 0
C58371 _0462_ hold73/a_391_47# 0.00622f
C58372 hold37/a_285_47# _1045_/a_193_47# 0
C58373 hold37/a_391_47# _1045_/a_27_47# 0.00179f
C58374 net1 _0584_/a_27_297# 0
C58375 _0834_/a_109_297# _0433_ 0
C58376 net211 _0580_/a_373_47# 0
C58377 _0352_ _0391_ 0.12694f
C58378 VPWR _0565_/a_240_47# 0.00319f
C58379 _0243_ _0249_ 0
C58380 clknet_0__0464_ net170 0
C58381 _0195_ _0997_/a_193_47# 0
C58382 comp0.B\[11\] hold51/a_49_47# 0.30972f
C58383 net202 clknet_1_0__leaf__0461_ 0.00304f
C58384 _0316_ _0324_ 0
C58385 A[7] net12 0.1369f
C58386 acc0.A\[4\] _0270_ 0.15792f
C58387 clknet_1_1__leaf__0463_ clknet_1_0__leaf__0461_ 0.04028f
C58388 _0351_ clknet_1_1__leaf__0462_ 0.01167f
C58389 clkload0/X _1072_/a_193_47# 0
C58390 _0314_ clkbuf_1_0__f__0462_/a_110_47# 0.10284f
C58391 hold67/a_49_47# clkbuf_1_1__f__0465_/a_110_47# 0
C58392 comp0.B\[13\] _1045_/a_975_413# 0
C58393 _0621_/a_285_297# _0253_ 0.11503f
C58394 acc0.A\[4\] _0987_/a_466_413# 0.01935f
C58395 comp0.B\[1\] _0178_ 0
C58396 hold66/a_285_47# _0345_ 0
C58397 _0984_/a_27_47# _0263_ 0
C58398 _0650_/a_68_297# net79 0
C58399 net61 _0458_ 0.25276f
C58400 clknet_1_0__leaf__0463_ net180 0.32169f
C58401 _0324_ _0347_ 0
C58402 _0482_ _0946_/a_30_53# 0
C58403 acc0.A\[29\] _0701_/a_209_47# 0
C58404 _1046_/a_891_413# _1045_/a_1059_315# 0
C58405 net14 _0180_ 0.08165f
C58406 _0661_/a_277_297# _0289_ 0.00141f
C58407 _0661_/a_205_297# _0287_ 0
C58408 pp[16] _1013_/a_1059_315# 0.00206f
C58409 _1017_/a_27_47# net166 0.01384f
C58410 net103 _1016_/a_193_47# 0.03462f
C58411 _0581_/a_27_297# _0352_ 0
C58412 _0399_ _0674_/a_113_47# 0
C58413 _0554_/a_68_297# comp0.B\[4\] 0.02761f
C58414 clknet_1_1__leaf__0459_ _0587_/a_27_47# 0.00265f
C58415 _0174_ B[13] 0
C58416 _0856_/a_79_21# _0465_ 0.0105f
C58417 _0274_ _0255_ 0.14115f
C58418 _0082_ net47 0.07631f
C58419 _0483_ _1068_/a_27_47# 0.002f
C58420 control0.count\[3\] _1068_/a_634_159# 0
C58421 _0222_ hold4/a_285_47# 0.00715f
C58422 hold81/a_49_47# hold81/a_391_47# 0.00188f
C58423 _0782_/a_27_47# acc0.A\[1\] 0
C58424 _1028_/a_634_159# _1028_/a_381_47# 0
C58425 _1030_/a_27_47# _0354_ 0
C58426 _0473_ _1042_/a_27_47# 0
C58427 acc0.A\[2\] _0856_/a_79_21# 0
C58428 _0343_ _0996_/a_193_47# 0.00352f
C58429 acc0.A\[7\] _0369_ 0.00125f
C58430 _0369_ _0989_/a_1059_315# 0.00781f
C58431 _0399_ _0406_ 0
C58432 _0441_ _0835_/a_493_297# 0
C58433 clknet_1_0__leaf__0458_ _0633_/a_109_297# 0
C58434 _0671_/a_113_297# clkbuf_1_1__f__0459_/a_110_47# 0.00167f
C58435 _0115_ hold72/a_391_47# 0.00309f
C58436 _0765_/a_79_21# clknet_1_0__leaf__0457_ 0.00119f
C58437 _0306_ _1009_/a_975_413# 0
C58438 _0144_ net132 0.00104f
C58439 _0852_/a_285_297# _0346_ 0.06388f
C58440 hold57/a_285_47# _0549_/a_68_297# 0
C58441 _0985_/a_975_413# VPWR 0.00464f
C58442 hold27/a_285_47# comp0.B\[9\] 0.00125f
C58443 pp[30] hold61/a_285_47# 0.0088f
C58444 VPWR _1018_/a_561_413# 0.00225f
C58445 _0722_/a_215_47# net239 0
C58446 output39/a_27_47# net80 0
C58447 net211 control0.add 0
C58448 _0557_/a_51_297# _1037_/a_27_47# 0
C58449 VPWR _1049_/a_891_413# 0.18994f
C58450 net15 input11/a_75_212# 0.00144f
C58451 clknet_0__0459_ clkload3/Y 0
C58452 _0233_ VPWR 0.53475f
C58453 _0593_/a_113_47# _0225_ 0.00992f
C58454 _0123_ _0352_ 0
C58455 _0575_/a_109_297# VPWR 0.19822f
C58456 _1041_/a_466_413# net31 0.02584f
C58457 pp[15] _0797_/a_27_413# 0.00187f
C58458 _0460_ _1006_/a_27_47# 0.04409f
C58459 hold97/a_285_47# _1008_/a_634_159# 0
C58460 hold97/a_391_47# _1008_/a_193_47# 0
C58461 _0751_/a_29_53# _0460_ 0
C58462 VPWR _1066_/a_891_413# 0.20826f
C58463 _0981_/a_109_297# _0480_ 0
C58464 _0137_ clknet_1_1__leaf__0457_ 0
C58465 _0745_/a_109_47# _0324_ 0
C58466 VPWR _1068_/a_891_413# 0.17471f
C58467 _0968_/a_109_297# _0488_ 0
C58468 _0455_ _0853_/a_150_297# 0
C58469 _1053_/a_1059_315# input11/a_75_212# 0
C58470 _0476_ _0946_/a_30_53# 0
C58471 _0366_ _0219_ 0.00812f
C58472 _0153_ clknet_1_1__leaf__0465_ 0.01389f
C58473 _1051_/a_891_413# _0987_/a_193_47# 0
C58474 _0346_ net247 0
C58475 _0993_/a_193_47# _0091_ 0.23509f
C58476 _0993_/a_466_413# _0419_ 0
C58477 _0993_/a_891_413# _0417_ 0
C58478 net69 _1018_/a_27_47# 0
C58479 _0518_/a_109_47# acc0.A\[8\] 0
C58480 comp0.B\[14\] net131 0.00104f
C58481 _0828_/a_199_47# _0436_ 0.00151f
C58482 _0661_/a_27_297# clknet_1_1__leaf__0465_ 0.01579f
C58483 _0750_/a_27_47# _0237_ 0.0283f
C58484 hold32/a_285_47# A[9] 0.08267f
C58485 _0140_ _1043_/a_891_413# 0.00617f
C58486 net198 _1043_/a_592_47# 0
C58487 hold39/a_49_47# _1035_/a_27_47# 0
C58488 hold76/a_391_47# _0771_/a_27_413# 0.00346f
C58489 hold76/a_285_47# _0771_/a_215_297# 0.0023f
C58490 clknet_1_0__leaf__0464_ _0196_ 0.06118f
C58491 clknet_1_0__leaf__0465_ _1046_/a_891_413# 0.00186f
C58492 _0531_/a_109_297# net9 0.01479f
C58493 _0343_ _0983_/a_975_413# 0
C58494 _0292_ _0990_/a_1059_315# 0
C58495 _0767_/a_59_75# _0245_ 0
C58496 hold25/a_285_47# net171 0.0011f
C58497 hold25/a_49_47# _0207_ 0.00708f
C58498 _0996_/a_27_47# net5 0.05651f
C58499 clkbuf_1_0__f_clk/a_110_47# _1068_/a_193_47# 0
C58500 output64/a_27_47# output58/a_27_47# 0
C58501 _0662_/a_299_297# acc0.A\[9\] 0.00343f
C58502 _1002_/a_592_47# acc0.A\[20\] 0
C58503 _0998_/a_891_413# _0998_/a_975_413# 0.00851f
C58504 _0998_/a_27_47# net84 0.30014f
C58505 _0998_/a_381_47# _0998_/a_561_413# 0.00123f
C58506 net45 _0793_/a_512_297# 0
C58507 _0710_/a_109_47# _0220_ 0
C58508 _0803_/a_150_297# _0403_ 0
C58509 _0649_/a_113_47# acc0.A\[10\] 0
C58510 net58 _0449_ 0
C58511 _0804_/a_79_21# net80 0
C58512 _1009_/a_466_413# _0318_ 0
C58513 clknet_1_0__leaf__0460_ _0756_/a_47_47# 0.00348f
C58514 _0621_/a_285_297# net74 0
C58515 acc0.A\[12\] hold45/a_285_47# 0
C58516 net247 _0935_/a_27_47# 0.02994f
C58517 _1003_/a_592_47# _0369_ 0
C58518 _0101_ _0762_/a_297_297# 0
C58519 _0346_ _0825_/a_68_297# 0
C58520 net7 _1061_/a_27_47# 0.02619f
C58521 net247 _1061_/a_193_47# 0.00126f
C58522 _0094_ _0400_ 0
C58523 _0183_ _0345_ 0.41363f
C58524 _1024_/a_1059_315# acc0.A\[23\] 0
C58525 net203 _1033_/a_193_47# 0.03196f
C58526 _0259_ _0986_/a_1059_315# 0
C58527 clknet_0__0463_ comp0.B\[5\] 0
C58528 clkbuf_1_1__f__0463_/a_110_47# _0474_ 0
C58529 _0984_/a_193_47# net47 0.02906f
C58530 _0346_ _0844_/a_382_297# 0
C58531 hold38/a_285_47# comp0.B\[6\] 0.0069f
C58532 hold38/a_391_47# comp0.B\[5\] 0
C58533 _0478_ clkbuf_1_0__f_clk/a_110_47# 0.02633f
C58534 _1019_/a_634_159# _1019_/a_592_47# 0
C58535 _0714_/a_51_297# _0714_/a_245_297# 0.01218f
C58536 _1058_/a_634_159# net37 0
C58537 _0629_/a_59_75# net247 0.00814f
C58538 _0123_ _0574_/a_109_297# 0.00469f
C58539 _0965_/a_47_47# _0965_/a_377_297# 0.00899f
C58540 hold42/a_285_47# _0188_ 0.06826f
C58541 net65 _0825_/a_68_297# 0.00125f
C58542 clknet_1_1__leaf__0463_ _0959_/a_217_297# 0
C58543 net72 _0986_/a_891_413# 0
C58544 _0440_ _0172_ 0.08775f
C58545 clknet_1_0__leaf__0464_ _0199_ 0
C58546 VPWR _1012_/a_975_413# 0.00549f
C58547 _0097_ _0219_ 0
C58548 _0553_/a_51_297# clkbuf_1_0__f__0463_/a_110_47# 0
C58549 hold54/a_391_47# _0208_ 0.07783f
C58550 _0482_ _0487_ 0
C58551 _1004_/a_1059_315# net46 0
C58552 net22 _0545_/a_150_297# 0.00128f
C58553 _1030_/a_27_47# _0567_/a_27_297# 0
C58554 _1051_/a_27_47# acc0.A\[4\] 0.00132f
C58555 acc0.A\[5\] _1050_/a_27_47# 0.00128f
C58556 _0399_ _0307_ 0.04213f
C58557 net201 _0175_ 0.08251f
C58558 net61 clkbuf_1_1__f__0458_/a_110_47# 0
C58559 _0475_ _0176_ 0.09283f
C58560 _0726_/a_51_297# _0726_/a_240_47# 0.03076f
C58561 acc0.A\[4\] _1045_/a_634_159# 0
C58562 _1050_/a_891_413# net184 0
C58563 hold9/a_285_47# net114 0
C58564 _0183_ hold2/a_49_47# 0.00421f
C58565 acc0.A\[8\] net62 0.02756f
C58566 _1058_/a_1059_315# net67 0.00292f
C58567 hold24/a_49_47# net171 0.03504f
C58568 net68 clkbuf_0__0457_/a_110_47# 0
C58569 _1033_/a_1059_315# _1032_/a_1059_315# 0
C58570 _0729_/a_68_297# _1010_/a_1059_315# 0.01105f
C58571 net36 clkbuf_1_1__f__0457_/a_110_47# 0.08112f
C58572 hold100/a_285_47# _0350_ 0.0149f
C58573 net9 _1049_/a_1017_47# 0.00116f
C58574 net175 net135 0
C58575 _1013_/a_193_47# _0220_ 0
C58576 clknet_1_0__leaf__0458_ _1060_/a_193_47# 0
C58577 hold55/a_49_47# _1032_/a_193_47# 0
C58578 hold55/a_285_47# _1032_/a_27_47# 0.00319f
C58579 _0316_ _0347_ 0.00143f
C58580 _0717_/a_80_21# hold61/a_285_47# 0
C58581 _0717_/a_209_297# hold61/a_49_47# 0
C58582 _0718_/a_47_47# _0129_ 0
C58583 _0222_ _0599_/a_113_47# 0
C58584 _1050_/a_27_47# _0528_/a_299_297# 0
C58585 _1050_/a_193_47# _0528_/a_81_21# 0
C58586 clknet_1_0__leaf__0465_ _0256_ 0.00265f
C58587 hold26/a_285_47# net22 0.03914f
C58588 _0180_ _0585_/a_109_297# 0
C58589 net159 _0468_ 0
C58590 VPWR _0998_/a_466_413# 0.25441f
C58591 _0338_ hold61/a_391_47# 0.05135f
C58592 clknet_1_0__leaf__0465_ _0987_/a_1059_315# 0.00965f
C58593 clknet_1_0__leaf__0463_ _0545_/a_150_297# 0
C58594 _0991_/a_193_47# _0450_ 0
C58595 _0990_/a_27_47# clknet_1_1__leaf__0465_ 0
C58596 _0758_/a_510_47# _0352_ 0.00142f
C58597 _0758_/a_215_47# _0102_ 0
C58598 acc0.A\[20\] _0384_ 0
C58599 _1024_/a_1017_47# net52 0
C58600 _0991_/a_891_413# _0218_ 0
C58601 net219 _0116_ 0.00573f
C58602 net145 net47 0
C58603 _0990_/a_466_413# _0990_/a_592_47# 0.00553f
C58604 _0990_/a_634_159# _0990_/a_1017_47# 0
C58605 _0343_ _0109_ 0.00442f
C58606 _0461_ _0771_/a_382_47# 0
C58607 hold81/a_49_47# _0281_ 0.01109f
C58608 acc0.A\[15\] _0345_ 0.04428f
C58609 _0790_/a_285_47# _0219_ 0.00301f
C58610 _0546_/a_51_297# net153 0
C58611 _0955_/a_32_297# _1066_/a_27_47# 0
C58612 _1002_/a_381_47# clknet_1_0__leaf__0457_ 0
C58613 _1056_/a_1017_47# _0187_ 0
C58614 _1002_/a_1059_315# _0460_ 0.01934f
C58615 _1032_/a_27_47# _0165_ 0
C58616 _0537_/a_68_297# _1043_/a_193_47# 0
C58617 _0537_/a_150_297# _1043_/a_27_47# 0
C58618 net70 net58 0
C58619 clknet_1_0__leaf__0463_ hold26/a_285_47# 0.00423f
C58620 net59 _0720_/a_68_297# 0
C58621 _0556_/a_68_297# _1035_/a_193_47# 0
C58622 net8 comp0.B\[10\] 0
C58623 net216 _0352_ 0.05096f
C58624 acc0.A\[16\] _1060_/a_193_47# 0
C58625 _0518_/a_27_297# acc0.A\[5\] 0
C58626 _0083_ acc0.A\[3\] 0.00844f
C58627 hold86/a_285_47# _0269_ 0.00184f
C58628 _0967_/a_109_93# _0476_ 0.08656f
C58629 _0770_/a_79_21# net46 0.06277f
C58630 _0476_ _0487_ 0
C58631 _0346_ net100 0
C58632 _1065_/a_27_47# _0951_/a_209_311# 0
C58633 _0488_ _0486_ 0.21135f
C58634 _0466_ control0.state\[2\] 0.99831f
C58635 comp0.B\[10\] net32 0.02263f
C58636 hold75/a_49_47# net165 0
C58637 net200 _1025_/a_193_47# 0.34157f
C58638 hold66/a_391_47# clknet_1_0__leaf__0460_ 0.00482f
C58639 _0802_/a_59_75# _0802_/a_145_75# 0.00658f
C58640 _0217_ _0611_/a_68_297# 0
C58641 _0743_/a_245_297# _0319_ 0
C58642 _0465_ _0846_/a_51_297# 0.01062f
C58643 hold2/a_49_47# acc0.A\[15\] 0
C58644 _0216_ _0778_/a_68_297# 0
C58645 _1051_/a_27_47# _1051_/a_466_413# 0.27314f
C58646 _1051_/a_193_47# _1051_/a_634_159# 0.11897f
C58647 hold9/a_285_47# _0365_ 0
C58648 output44/a_27_47# VPWR 0.25155f
C58649 _1056_/a_27_47# clknet_1_1__leaf__0465_ 0.00872f
C58650 clknet_1_1__leaf__0459_ VPWR 4.55368f
C58651 acc0.A\[14\] _0849_/a_79_21# 0.06206f
C58652 _0294_ clknet_0__0461_ 0.02449f
C58653 _1070_/a_466_413# _0168_ 0.00321f
C58654 _0230_ _0352_ 0.06712f
C58655 _1070_/a_891_413# VPWR 0.19113f
C58656 _1070_/a_27_47# control0.count\[1\] 0.00129f
C58657 net106 _1033_/a_466_413# 0
C58658 _1045_/a_193_47# _1045_/a_381_47# 0.10164f
C58659 _1045_/a_634_159# _1045_/a_891_413# 0.03684f
C58660 _1045_/a_27_47# _1045_/a_561_413# 0.0027f
C58661 _0480_ _1069_/a_27_47# 0
C58662 _1003_/a_27_47# hold66/a_49_47# 0
C58663 _0478_ control0.count\[2\] 0.0639f
C58664 _0217_ net109 0.02194f
C58665 net150 net177 0
C58666 VPWR _1043_/a_27_47# 0.69674f
C58667 _0678_/a_68_297# _0308_ 0.17708f
C58668 _1014_/a_975_413# _0465_ 0
C58669 _0552_/a_150_297# net29 0
C58670 VPWR _1030_/a_975_413# 0.00441f
C58671 net67 net47 0
C58672 _0313_ _0105_ 0.14286f
C58673 _0783_/a_215_47# _0397_ 0.04866f
C58674 _0378_ _0219_ 0.00202f
C58675 _0733_/a_222_93# _0697_/a_80_21# 0
C58676 _1043_/a_193_47# _1043_/a_381_47# 0.09503f
C58677 _1043_/a_634_159# _1043_/a_891_413# 0.03684f
C58678 _1043_/a_27_47# _1043_/a_561_413# 0.0027f
C58679 comp0.B\[2\] _0175_ 0.80541f
C58680 hold32/a_285_47# _0516_/a_27_297# 0
C58681 net64 net62 0.0269f
C58682 hold64/a_285_47# _0346_ 0
C58683 _0502_/a_27_47# _0181_ 0.33408f
C58684 clknet_1_1__leaf__0459_ _0654_/a_27_413# 0.01844f
C58685 _1038_/a_381_47# _0209_ 0
C58686 net236 control0.state\[2\] 0.02811f
C58687 clkbuf_0__0464_/a_110_47# clknet_1_1__leaf__0464_ 0.00118f
C58688 _1004_/a_891_413# VPWR 0.19368f
C58689 _1021_/a_193_47# _1002_/a_381_47# 0
C58690 hold89/a_285_47# _0487_ 0.05559f
C58691 _0775_/a_79_21# _0392_ 0.05518f
C58692 _1054_/a_27_47# _1054_/a_634_159# 0.14145f
C58693 net187 _0586_/a_27_47# 0
C58694 _0736_/a_311_297# clknet_1_1__leaf__0460_ 0
C58695 _1071_/a_193_47# clknet_1_0__leaf_clk 0.01121f
C58696 _0179_ _0345_ 0.17986f
C58697 VPWR _0171_ 1.03904f
C58698 _0730_/a_79_21# _1010_/a_27_47# 0
C58699 _0182_ _0208_ 0.13426f
C58700 _0982_/a_27_47# acc0.A\[1\] 0
C58701 comp0.B\[10\] _1042_/a_1059_315# 0.08555f
C58702 net194 _1044_/a_381_47# 0.115f
C58703 _0241_ _0386_ 0
C58704 _0792_/a_80_21# _0792_/a_209_47# 0.01013f
C58705 _0987_/a_381_47# _0085_ 0.13418f
C58706 _0345_ hold40/a_285_47# 0
C58707 net53 _0697_/a_217_297# 0
C58708 _0849_/a_215_47# _0451_ 0.00837f
C58709 _0292_ VPWR 0.78155f
C58710 acc0.A\[1\] _0145_ 0
C58711 _0476_ net119 0
C58712 control0.state\[2\] _1064_/a_193_47# 0
C58713 _0458_ _0431_ 0.00385f
C58714 net162 _0219_ 0
C58715 acc0.A\[27\] _0328_ 0
C58716 _0217_ pp[24] 0
C58717 _0684_/a_59_75# _0350_ 0
C58718 _0972_/a_250_297# _0471_ 0.01421f
C58719 input9/a_27_47# A[2] 0.20222f
C58720 _0343_ _0794_/a_326_47# 0
C58721 _0557_/a_51_297# _0133_ 0
C58722 _0557_/a_245_297# net121 0
C58723 _0134_ _1035_/a_193_47# 0
C58724 _0727_/a_109_47# _0356_ 0
C58725 clkbuf_0__0465_/a_110_47# _0347_ 0
C58726 hold47/a_391_47# _0196_ 0
C58727 comp0.B\[10\] net10 0.05938f
C58728 _0642_/a_215_297# _0432_ 0
C58729 _1059_/a_466_413# _0158_ 0
C58730 _0820_/a_79_21# hold67/a_285_47# 0
C58731 _0541_/a_68_297# net20 0
C58732 net27 _0176_ 0
C58733 _0983_/a_27_47# _0983_/a_891_413# 0.03089f
C58734 _0983_/a_193_47# _0983_/a_1059_315# 0.03405f
C58735 _0983_/a_634_159# _0983_/a_466_413# 0.23992f
C58736 _0311_ _0312_ 0.01533f
C58737 hold34/a_391_47# net16 0
C58738 clknet_1_0__leaf__0465_ _1051_/a_193_47# 0.00843f
C58739 output41/a_27_47# net41 0.19769f
C58740 clknet_1_0__leaf__0465_ _1045_/a_466_413# 0.00265f
C58741 hold98/a_285_47# _0995_/a_193_47# 0.00185f
C58742 hold98/a_391_47# _0995_/a_27_47# 0
C58743 _0558_/a_68_297# _0557_/a_51_297# 0
C58744 _1029_/a_381_47# net191 0.12065f
C58745 hold37/a_49_47# net131 0
C58746 _0246_ _0350_ 0
C58747 net88 net23 0
C58748 net46 pp[19] 0.05079f
C58749 net59 net116 0.07298f
C58750 _0770_/a_382_297# VPWR 0.00511f
C58751 VPWR _0435_ 0.31521f
C58752 net55 hold95/a_285_47# 0
C58753 _0343_ acc0.A\[6\] 0.09205f
C58754 acc0.A\[1\] _0446_ 0
C58755 acc0.A\[26\] _0345_ 0
C58756 net17 _0950_/a_75_212# 0
C58757 net101 _0181_ 0.00206f
C58758 _0328_ _0364_ 0.00479f
C58759 _0581_/a_27_297# hold72/a_285_47# 0
C58760 _1015_/a_193_47# _0526_/a_27_47# 0
C58761 acc0.A\[24\] _0219_ 0.06439f
C58762 _0260_ _0640_/a_109_53# 0.00133f
C58763 _1015_/a_27_47# _0566_/a_27_47# 0
C58764 acc0.A\[4\] _0085_ 0.04804f
C58765 acc0.A\[12\] _0301_ 0.02683f
C58766 clknet_1_0__leaf__0459_ _0998_/a_466_413# 0
C58767 A[11] net143 0
C58768 _0113_ _0565_/a_240_47# 0
C58769 _1020_/a_561_413# _0183_ 0.00157f
C58770 clknet_0__0465_ _0271_ 0.04337f
C58771 _1003_/a_193_47# _0217_ 0.00713f
C58772 _0371_ _0326_ 0.01697f
C58773 _0956_/a_32_297# _0956_/a_220_297# 0.00132f
C58774 _0806_/a_199_47# _0418_ 0.00151f
C58775 _1013_/a_634_159# _0218_ 0.01586f
C58776 net235 _0350_ 0.00298f
C58777 _1016_/a_466_413# _1016_/a_561_413# 0.00772f
C58778 _1016_/a_634_159# _1016_/a_975_413# 0
C58779 hold25/a_285_47# _1037_/a_466_413# 0
C58780 hold25/a_49_47# _1037_/a_1059_315# 0
C58781 _0251_ hold31/a_49_47# 0.01252f
C58782 _0548_/a_512_297# net147 0
C58783 VPWR _0726_/a_240_47# 0.00167f
C58784 net205 net24 0
C58785 net59 hold92/a_285_47# 0.13073f
C58786 acc0.A\[20\] _0383_ 0
C58787 hold87/a_285_47# acc0.A\[14\] 0
C58788 comp0.B\[1\] _0956_/a_114_297# 0.00153f
C58789 clknet_1_1__leaf__0462_ _1026_/a_27_47# 0.00538f
C58790 _1028_/a_381_47# net114 0
C58791 _1028_/a_634_159# acc0.A\[28\] 0
C58792 net49 _0760_/a_285_47# 0
C58793 net9 A[2] 0.0701f
C58794 _0130_ comp0.B\[15\] 0.11777f
C58795 _0236_ _0352_ 0
C58796 _1057_/a_891_413# _0187_ 0.03292f
C58797 _0213_ _0560_/a_150_297# 0
C58798 _0744_/a_27_47# net143 0.00189f
C58799 _0173_ _0560_/a_68_297# 0.00317f
C58800 net99 clknet_1_1__leaf__0462_ 0
C58801 VPWR _0990_/a_975_413# 0.00467f
C58802 _0812_/a_510_47# _0422_ 0.00254f
C58803 _0542_/a_240_47# hold51/a_285_47# 0
C58804 _0343_ _0725_/a_80_21# 0.12424f
C58805 VPWR _0793_/a_512_297# 0.00735f
C58806 pp[10] net67 0.01202f
C58807 _0733_/a_222_93# _0345_ 0
C58808 _0136_ _0176_ 0.04955f
C58809 clkbuf_1_0__f__0462_/a_110_47# _0360_ 0
C58810 _0626_/a_68_297# _0445_ 0
C58811 net58 _0260_ 0
C58812 net39 _0994_/a_634_159# 0.0372f
C58813 input3/a_75_212# A[11] 0.23493f
C58814 hold45/a_49_47# _0179_ 0.00813f
C58815 _1059_/a_466_413# acc0.A\[14\] 0.04422f
C58816 _0584_/a_27_297# net157 0.0661f
C58817 net102 clknet_1_1__leaf__0461_ 0.2615f
C58818 _1041_/a_466_413# net7 0.03301f
C58819 _0211_ B[1] 0.01483f
C58820 _0554_/a_68_297# _1035_/a_193_47# 0
C58821 _0195_ clknet_1_0__leaf__0457_ 0
C58822 hold4/a_391_47# _1022_/a_634_159# 0
C58823 hold4/a_49_47# _1022_/a_1059_315# 0
C58824 hold4/a_285_47# _1022_/a_466_413# 0.0041f
C58825 _0094_ clkbuf_0__0459_/a_110_47# 0.01341f
C58826 net16 _0181_ 0.15732f
C58827 _0984_/a_193_47# _0294_ 0
C58828 _0984_/a_27_47# _0218_ 0
C58829 hold31/a_49_47# net58 0
C58830 _0146_ _1047_/a_27_47# 0
C58831 hold97/a_285_47# net94 0
C58832 hold46/a_49_47# _0139_ 0
C58833 _0170_ _1072_/a_381_47# 0.11702f
C58834 control0.count\[3\] _0479_ 0
C58835 output45/a_27_47# pp[18] 0.15722f
C58836 hold29/a_49_47# hold29/a_285_47# 0.22264f
C58837 _0504_/a_27_47# VPWR 0.41126f
C58838 hold20/a_49_47# _0468_ 0.00799f
C58839 hold23/a_285_47# hold23/a_391_47# 0.41909f
C58840 _1047_/a_27_47# _0492_/a_27_47# 0
C58841 _0343_ _0128_ 0.031f
C58842 _1054_/a_466_413# VPWR 0.25407f
C58843 _0357_ net57 0
C58844 acc0.A\[5\] _0987_/a_27_47# 0.0033f
C58845 _1051_/a_1059_315# net73 0.0105f
C58846 _1051_/a_466_413# _0085_ 0
C58847 clknet_1_0__leaf__0462_ _1025_/a_381_47# 0.00918f
C58848 net231 hold84/a_285_47# 0.0101f
C58849 clknet_1_1__leaf__0459_ _0283_ 0.04102f
C58850 _0286_ acc0.A\[11\] 0
C58851 _0770_/a_297_47# _0243_ 0.05417f
C58852 _0770_/a_382_297# _0390_ 0.00188f
C58853 _0512_/a_27_297# net3 0.1887f
C58854 _1038_/a_634_159# VPWR 0.18649f
C58855 _0293_ clknet_1_1__leaf__0465_ 0.01978f
C58856 net233 _0350_ 0.058f
C58857 _0456_ VPWR 0.29727f
C58858 net154 _0524_/a_109_297# 0.0083f
C58859 _1041_/a_634_159# A[15] 0
C58860 _0222_ output51/a_27_47# 0
C58861 VPWR _0655_/a_215_53# 0.13589f
C58862 pp[0] clknet_1_0__leaf__0463_ 0.00872f
C58863 net36 net123 0
C58864 _1018_/a_1059_315# acc0.A\[18\] 0.12589f
C58865 _0183_ _0576_/a_109_47# 0
C58866 _0322_ _0319_ 0.65281f
C58867 net232 _0468_ 0
C58868 hold74/a_285_47# _0219_ 0.01424f
C58869 _1028_/a_381_47# _0365_ 0.00125f
C58870 _0247_ _0460_ 0
C58871 net81 _0668_/a_297_47# 0
C58872 _0996_/a_592_47# _0185_ 0
C58873 _0174_ _0495_/a_68_297# 0
C58874 clknet_0__0458_ _0258_ 0.01111f
C58875 clknet_0_clk _1068_/a_592_47# 0
C58876 _0327_ _0319_ 0
C58877 clkbuf_1_0__f__0457_/a_110_47# _0460_ 0
C58878 net45 _0095_ 0.00226f
C58879 _0627_/a_215_53# _0346_ 0.07041f
C58880 _0755_/a_109_297# _0377_ 0
C58881 hold14/a_49_47# _0557_/a_51_297# 0
C58882 clkbuf_1_1__f__0463_/a_110_47# _0563_/a_51_297# 0.00717f
C58883 hold30/a_49_47# _0121_ 0.29996f
C58884 net44 _0567_/a_27_297# 0
C58885 _0369_ _0988_/a_466_413# 0
C58886 _1019_/a_193_47# clkbuf_1_0__f__0461_/a_110_47# 0
C58887 VPWR _0785_/a_299_297# 0.19426f
C58888 _1001_/a_1059_315# _0195_ 0
C58889 _1019_/a_1059_315# _0350_ 0.0018f
C58890 _1053_/a_27_47# _0519_/a_81_21# 0
C58891 _0781_/a_68_297# net221 0
C58892 net145 _0294_ 0
C58893 _0130_ net203 0
C58894 _1052_/a_1059_315# _0087_ 0
C58895 _1019_/a_592_47# net105 0
C58896 _0315_ _0318_ 0
C58897 net144 net37 0.00609f
C58898 _0817_/a_266_297# _0346_ 0.00252f
C58899 _0857_/a_27_47# _1067_/a_193_47# 0
C58900 net35 _1071_/a_1059_315# 0.00914f
C58901 _0965_/a_285_47# _0483_ 0.04387f
C58902 B[15] B[5] 0.00212f
C58903 input6/a_75_212# _0297_ 0
C58904 net51 _1005_/a_975_413# 0
C58905 clknet_1_1__leaf__0460_ _0697_/a_80_21# 0
C58906 comp0.B\[13\] _1042_/a_634_159# 0
C58907 _0216_ hold8/a_391_47# 0.00183f
C58908 _0108_ acc0.A\[27\] 0.09339f
C58909 _0172_ net18 0.08756f
C58910 _0535_/a_68_297# net31 0
C58911 clknet_1_1__leaf__0460_ net56 0.24217f
C58912 _1038_/a_193_47# _0550_/a_51_297# 0
C58913 _0674_/a_113_47# _0306_ 0.00957f
C58914 _0381_ hold3/a_49_47# 0.00501f
C58915 _0469_ _0161_ 0.03056f
C58916 net66 net143 0.02015f
C58917 _0323_ _0181_ 0
C58918 net173 net174 0.00339f
C58919 _0343_ _0995_/a_1059_315# 0
C58920 _1014_/a_891_413# clknet_1_0__leaf__0461_ 0.00629f
C58921 acc0.A\[4\] net131 0
C58922 _0575_/a_373_47# net50 0
C58923 _0726_/a_512_297# _0109_ 0
C58924 _0668_/a_79_21# net6 0.02144f
C58925 net8 _0177_ 0
C58926 clknet_1_1__leaf__0463_ input25/a_75_212# 0.00268f
C58927 _0673_/a_253_47# acc0.A\[13\] 0
C58928 clknet_0__0461_ _0581_/a_109_297# 0
C58929 _0458_ _0269_ 0.01036f
C58930 _0654_/a_207_413# _0281_ 0.01458f
C58931 comp0.B\[14\] _0139_ 0
C58932 _0180_ _0178_ 0.17648f
C58933 _0292_ _0283_ 0
C58934 _0800_/a_149_47# clknet_1_1__leaf__0459_ 0.0066f
C58935 net34 _1064_/a_891_413# 0.04256f
C58936 control0.state\[1\] _1064_/a_381_47# 0
C58937 _0316_ _0106_ 0
C58938 _0178_ net218 0
C58939 _1033_/a_891_413# clknet_1_1__leaf__0463_ 0
C58940 _1015_/a_634_159# net157 0.00258f
C58941 hold18/a_391_47# _0850_/a_68_297# 0
C58942 _0348_ hold61/a_391_47# 0
C58943 _0286_ hold81/a_391_47# 0
C58944 _1050_/a_1059_315# _0148_ 0
C58945 net68 _0350_ 0
C58946 _0716_/a_27_47# _0304_ 0.05539f
C58947 net40 _0413_ 0
C58948 _1059_/a_193_47# net228 0
C58949 _0750_/a_27_47# _0222_ 0
C58950 _1001_/a_466_413# _0369_ 0
C58951 _0739_/a_297_297# _0365_ 0.00448f
C58952 clkbuf_1_0__f__0457_/a_110_47# _1001_/a_381_47# 0
C58953 clknet_0__0457_ _1001_/a_466_413# 0
C58954 _0467_ _1065_/a_466_413# 0.033f
C58955 _0347_ _0106_ 0.05784f
C58956 control0.state\[0\] _0981_/a_27_297# 0
C58957 net77 _0446_ 0
C58958 _0587_/a_27_47# _0095_ 0
C58959 _0195_ _1047_/a_891_413# 0.01148f
C58960 _0216_ _1047_/a_466_413# 0
C58961 _1014_/a_1059_315# _0265_ 0
C58962 hold12/a_391_47# _0486_ 0
C58963 _1021_/a_27_47# _0369_ 0
C58964 _0465_ _1048_/a_592_47# 0
C58965 pp[28] hold80/a_391_47# 0.00633f
C58966 _0996_/a_27_47# _0996_/a_634_159# 0.14145f
C58967 _0965_/a_285_47# control0.count\[1\] 0
C58968 _0675_/a_68_297# _0308_ 0
C58969 _0294_ net67 0.00547f
C58970 _0552_/a_150_297# comp0.B\[6\] 0
C58971 _0495_/a_68_297# _0208_ 0
C58972 _0990_/a_592_47# _0088_ 0.00188f
C58973 _0244_ _0246_ 0.02889f
C58974 _0388_ _0245_ 0.07433f
C58975 _0174_ net31 0.17871f
C58976 _0982_/a_891_413# _0264_ 0
C58977 _0999_/a_381_47# _0345_ 0
C58978 _0999_/a_634_159# _0219_ 0
C58979 _0793_/a_149_47# _0407_ 0.01702f
C58980 net7 _0953_/a_32_297# 0
C58981 output46/a_27_47# output50/a_27_47# 0
C58982 _0646_/a_47_47# acc0.A\[13\] 0.07313f
C58983 acc0.A\[16\] _1017_/a_1059_315# 0.01202f
C58984 _0949_/a_145_75# _0477_ 0
C58985 _0234_ _0754_/a_512_297# 0.00148f
C58986 _0375_ _0754_/a_51_297# 0
C58987 _0430_ output58/a_27_47# 0.01191f
C58988 _0195_ _0850_/a_68_297# 0
C58989 _0211_ _1035_/a_891_413# 0.00136f
C58990 clknet_1_1__leaf__0463_ net240 0
C58991 net46 net176 0.00475f
C58992 _0230_ _0237_ 0.03248f
C58993 net42 _0301_ 0.07939f
C58994 _0314_ _0324_ 0
C58995 _0313_ _0359_ 0.25789f
C58996 hold57/a_391_47# _0957_/a_32_297# 0
C58997 _1050_/a_1017_47# _0180_ 0
C58998 _0108_ _0110_ 0.00107f
C58999 VPWR _0996_/a_466_413# 0.26934f
C59000 _0191_ acc0.A\[5\] 0
C59001 _0691_/a_68_297# _0219_ 0.00505f
C59002 hold24/a_49_47# _0553_/a_51_297# 0.00134f
C59003 _1065_/a_466_413# comp0.B\[0\] 0.0052f
C59004 net143 _0350_ 0
C59005 _0643_/a_103_199# _0640_/a_109_53# 0
C59006 hold53/a_391_47# acc0.A\[25\] 0
C59007 hold68/a_285_47# net199 0
C59008 net215 _0575_/a_109_47# 0
C59009 _0682_/a_150_297# _0219_ 0
C59010 _0995_/a_381_47# acc0.A\[13\] 0
C59011 _1037_/a_891_413# net28 0.03305f
C59012 clknet_1_0__leaf__0461_ _0771_/a_27_413# 0
C59013 _0480_ _0489_ 0
C59014 _1051_/a_27_47# _0149_ 0.07322f
C59015 _1051_/a_193_47# net137 0.0067f
C59016 _1051_/a_1059_315# _1051_/a_1017_47# 0
C59017 hold65/a_285_47# _0830_/a_79_21# 0.00112f
C59018 _1045_/a_466_413# _1044_/a_466_413# 0.00119f
C59019 _1045_/a_193_47# _1044_/a_891_413# 0
C59020 _1045_/a_891_413# _1044_/a_193_47# 0.0011f
C59021 _0336_ _0704_/a_150_297# 0
C59022 _0227_ _1005_/a_891_413# 0
C59023 _0274_ _0989_/a_27_47# 0
C59024 _0992_/a_27_47# acc0.A\[10\] 0.02f
C59025 _1051_/a_466_413# net131 0
C59026 _1030_/a_27_47# _0353_ 0
C59027 _0837_/a_81_21# _0346_ 0.11897f
C59028 net160 net171 0
C59029 net62 _0986_/a_466_413# 0.02313f
C59030 _0467_ clknet_1_0__leaf__0460_ 0
C59031 net106 _0131_ 0
C59032 _1045_/a_891_413# net131 0
C59033 _1045_/a_1059_315# net184 0
C59034 clkbuf_1_0__f__0464_/a_110_47# _0196_ 0.00731f
C59035 clknet_1_1__leaf__0459_ _0789_/a_75_199# 0.00879f
C59036 hold56/a_49_47# _1032_/a_1059_315# 0
C59037 _0979_/a_109_297# control0.count\[0\] 0
C59038 net23 _1067_/a_891_413# 0.03836f
C59039 _1003_/a_1059_315# net213 0
C59040 _1072_/a_466_413# clknet_1_0__leaf_clk 0
C59041 _0370_ _0352_ 0
C59042 _0643_/a_253_297# _0465_ 0
C59043 _0276_ _0410_ 0
C59044 net63 _0180_ 0
C59045 _1002_/a_27_47# net240 0.08951f
C59046 _0984_/a_634_159# _0158_ 0
C59047 _0733_/a_448_47# _0322_ 0.00751f
C59048 _1043_/a_1059_315# net196 0
C59049 _1043_/a_891_413# net129 0
C59050 net46 _0617_/a_68_297# 0.00168f
C59051 clknet_1_0__leaf__0465_ clknet_0__0465_ 0.00393f
C59052 hold32/a_285_47# _0190_ 0
C59053 _1060_/a_193_47# _0506_/a_299_297# 0
C59054 VPWR _0568_/a_109_47# 0
C59055 VPWR _1015_/a_561_413# 0.00309f
C59056 net133 _0146_ 0
C59057 _0216_ _0782_/a_27_47# 0
C59058 acc0.A\[21\] _0765_/a_215_47# 0.0057f
C59059 clknet_1_0__leaf__0458_ _0982_/a_1059_315# 0
C59060 _0788_/a_68_297# _0346_ 0
C59061 _1016_/a_466_413# hold72/a_49_47# 0
C59062 net160 net24 0.38702f
C59063 _0210_ B[1] 0
C59064 _1072_/a_27_47# _0974_/a_222_93# 0
C59065 net46 hold68/a_49_47# 0.00147f
C59066 _0647_/a_47_47# _0399_ 0
C59067 control0.state\[0\] hold84/a_391_47# 0
C59068 control0.state\[1\] hold84/a_285_47# 0.00194f
C59069 net133 _0492_/a_27_47# 0
C59070 VPWR clkbuf_1_0__f_clk/a_110_47# 1.26702f
C59071 _1032_/a_27_47# _1032_/a_1059_315# 0.04875f
C59072 _1032_/a_193_47# _1032_/a_466_413# 0.08301f
C59073 _0461_ control0.add 0.0024f
C59074 _0748_/a_81_21# _0240_ 0.00111f
C59075 _1021_/a_1059_315# _0100_ 0
C59076 _1054_/a_891_413# _1054_/a_975_413# 0.00851f
C59077 _1054_/a_27_47# net140 0.23169f
C59078 _1054_/a_381_47# _1054_/a_561_413# 0.00123f
C59079 net158 clkbuf_0__0464_/a_110_47# 0.00771f
C59080 hold11/a_391_47# clknet_0__0464_ 0
C59081 _1071_/a_975_413# control0.count\[0\] 0
C59082 _1015_/a_466_413# _1015_/a_561_413# 0.00772f
C59083 _1015_/a_634_159# _1015_/a_975_413# 0
C59084 _0852_/a_35_297# _0850_/a_68_297# 0.001f
C59085 _0748_/a_81_21# _0369_ 0.06509f
C59086 _0983_/a_1017_47# VPWR 0
C59087 _0307_ _0306_ 0.07069f
C59088 _0991_/a_1059_315# _0347_ 0
C59089 clknet_1_1__leaf__0460_ _0345_ 0.40816f
C59090 _0108_ _1010_/a_193_47# 0.19393f
C59091 _0557_/a_149_47# _0173_ 0.01702f
C59092 _0557_/a_51_297# _0208_ 0.16305f
C59093 _0357_ _1010_/a_1059_315# 0
C59094 _0358_ _1010_/a_466_413# 0.00156f
C59095 _0432_ net63 0
C59096 _0369_ _0186_ 0.10593f
C59097 net51 _0360_ 0
C59098 _0352_ _0773_/a_285_47# 0
C59099 clknet_1_1__leaf__0462_ _1027_/a_975_413# 0
C59100 net113 _1027_/a_381_47# 0
C59101 _0335_ hold80/a_285_47# 0.01288f
C59102 clkbuf_1_0__f__0463_/a_110_47# _0206_ 0
C59103 _0792_/a_303_47# _0408_ 0
C59104 _0405_ _0400_ 0.40486f
C59105 _0989_/a_27_47# pp[5] 0
C59106 _0343_ _1031_/a_1059_315# 0
C59107 VPWR _0550_/a_149_47# 0.00187f
C59108 _0096_ clkbuf_1_1__f__0461_/a_110_47# 0.03251f
C59109 net247 _1047_/a_466_413# 0
C59110 _0203_ _0541_/a_150_297# 0
C59111 _1038_/a_634_159# _1038_/a_592_47# 0
C59112 _0211_ _1037_/a_634_159# 0
C59113 clkbuf_0__0460_/a_110_47# _0105_ 0
C59114 _1067_/a_193_47# net107 0
C59115 _1067_/a_466_413# clknet_1_0__leaf__0461_ 0.00594f
C59116 input1/a_27_47# input33/a_75_212# 0
C59117 hold19/a_49_47# _0369_ 0.00344f
C59118 net45 _0777_/a_285_47# 0
C59119 _0655_/a_215_53# _0283_ 0.14529f
C59120 _0290_ _0812_/a_215_47# 0
C59121 _0164_ _0471_ 0.00124f
C59122 net40 _0646_/a_129_47# 0.00435f
C59123 net59 _0220_ 0.06118f
C59124 clknet_1_0__leaf__0465_ _1044_/a_634_159# 0.00144f
C59125 clknet_1_0__leaf__0458_ _0451_ 0.0308f
C59126 _0157_ _0158_ 0
C59127 _0536_/a_51_297# _0498_/a_240_47# 0
C59128 _0536_/a_240_47# _0498_/a_51_297# 0
C59129 _0983_/a_466_413# net69 0
C59130 pp[16] output60/a_27_47# 0.01499f
C59131 _1011_/a_27_47# _0347_ 0
C59132 clkbuf_1_1__f__0465_/a_110_47# _0990_/a_1059_315# 0
C59133 hold86/a_285_47# clkbuf_0__0458_/a_110_47# 0
C59134 _0995_/a_1059_315# A[14] 0
C59135 _0332_ clknet_1_1__leaf__0462_ 0.02782f
C59136 clknet_1_0__leaf__0465_ net184 0.00773f
C59137 _0102_ _0350_ 0.13351f
C59138 _0352_ _0380_ 0.11629f
C59139 _0261_ _0447_ 0.00652f
C59140 net36 _0242_ 0
C59141 _0456_ _0453_ 0
C59142 _0627_/a_109_93# _0258_ 0.06884f
C59143 net40 _0995_/a_975_413# 0
C59144 net245 _0995_/a_381_47# 0.0237f
C59145 _0346_ _0406_ 0
C59146 clknet_1_0__leaf__0460_ _0374_ 0.03229f
C59147 _0286_ _0281_ 0.39127f
C59148 net188 _0511_/a_81_21# 0
C59149 _0659_/a_68_297# _0291_ 0.12615f
C59150 _0659_/a_150_297# acc0.A\[8\] 0
C59151 _0143_ comp0.B\[11\] 0
C59152 pp[28] _0336_ 0
C59153 hold69/a_391_47# VPWR 0.18896f
C59154 _0997_/a_634_159# net42 0.03021f
C59155 _0550_/a_51_297# _0550_/a_512_297# 0.0116f
C59156 _0430_ clkbuf_1_0__f__0465_/a_110_47# 0
C59157 _0116_ hold72/a_285_47# 0
C59158 _0747_/a_215_47# _1006_/a_466_413# 0
C59159 _0236_ _0237_ 0.01682f
C59160 _0368_ acc0.A\[23\] 0.00379f
C59161 acc0.A\[12\] _1058_/a_27_47# 0.01812f
C59162 _1056_/a_891_413# _0154_ 0
C59163 net90 _1007_/a_975_413# 0
C59164 hold21/a_391_47# clknet_1_0__leaf__0465_ 0
C59165 _1048_/a_27_47# _1047_/a_381_47# 0
C59166 _1048_/a_891_413# _1047_/a_193_47# 0
C59167 _1048_/a_466_413# _1047_/a_466_413# 0
C59168 net89 net150 0
C59169 _1054_/a_193_47# acc0.A\[6\] 0.00103f
C59170 _0117_ hold60/a_49_47# 0.38289f
C59171 net55 _0313_ 0
C59172 hold18/a_285_47# net149 0
C59173 _0317_ _0329_ 0.03797f
C59174 _1016_/a_561_413# net166 0
C59175 _1061_/a_466_413# acc0.A\[15\] 0
C59176 acc0.A\[5\] clkbuf_1_0__f__0465_/a_110_47# 0.02685f
C59177 hold25/a_285_47# _0135_ 0
C59178 _0138_ net147 0.12282f
C59179 hold31/a_285_47# _0254_ 0.00138f
C59180 clknet_0__0459_ _0996_/a_592_47# 0
C59181 _0247_ _0614_/a_29_53# 0
C59182 _0534_/a_81_21# hold71/a_285_47# 0
C59183 _0998_/a_381_47# _0398_ 0
C59184 _0998_/a_1059_315# _0096_ 0.00461f
C59185 _0998_/a_891_413# _0399_ 0
C59186 net114 acc0.A\[28\] 0
C59187 _0425_ _0347_ 0
C59188 _0314_ _0347_ 0
C59189 VPWR _0617_/a_150_297# 0.00193f
C59190 hold22/a_49_47# VPWR 0.26954f
C59191 control0.count\[2\] VPWR 0.56245f
C59192 hold11/a_285_47# clknet_1_0__leaf__0464_ 0
C59193 _0780_/a_285_47# _0308_ 0.00149f
C59194 _0535_/a_68_297# _0548_/a_240_47# 0
C59195 _0780_/a_35_297# _0394_ 0.00129f
C59196 _0327_ _0333_ 0.26427f
C59197 clknet_0__0458_ net72 0.00752f
C59198 VPWR _0095_ 0.34107f
C59199 comp0.B\[1\] _0496_/a_27_47# 0
C59200 _0773_/a_35_297# _0773_/a_117_297# 0.00641f
C59201 hold68/a_285_47# VPWR 0.28441f
C59202 _0361_ _0219_ 0.3305f
C59203 _0260_ clknet_1_0__leaf__0464_ 0
C59204 _0179_ _0156_ 0.00776f
C59205 acc0.A\[20\] _0749_/a_81_21# 0
C59206 _1008_/a_193_47# hold50/a_391_47# 0
C59207 _1052_/a_1059_315# net154 0
C59208 _1052_/a_193_47# net11 0.00846f
C59209 _0961_/a_199_47# _0466_ 0
C59210 _0216_ _0585_/a_373_47# 0
C59211 _0984_/a_1059_315# _0451_ 0
C59212 _0157_ acc0.A\[14\] 0.00998f
C59213 _0982_/a_27_47# _1014_/a_634_159# 0.00157f
C59214 _0985_/a_1059_315# _0219_ 0.00143f
C59215 _0201_ _0142_ 0.00247f
C59216 net21 net20 0.53032f
C59217 _0195_ _1017_/a_634_159# 0.01127f
C59218 hold64/a_391_47# _1001_/a_193_47# 0
C59219 hold64/a_285_47# _1001_/a_634_159# 0
C59220 _1057_/a_1017_47# acc0.A\[11\] 0
C59221 clk _0978_/a_27_297# 0.00154f
C59222 hold4/a_285_47# net151 0.01412f
C59223 hold48/a_285_47# net21 0
C59224 net120 _0563_/a_240_47# 0
C59225 _0255_ _0433_ 0.16764f
C59226 _0821_/a_113_47# _0179_ 0
C59227 net242 _0332_ 0
C59228 acc0.A\[0\] _0261_ 0
C59229 hold39/a_285_47# _0213_ 0.06706f
C59230 hold39/a_49_47# _0173_ 0.03367f
C59231 _1016_/a_466_413# clknet_0__0461_ 0
C59232 _0677_/a_47_47# _0308_ 0.0018f
C59233 hold17/a_285_47# clkbuf_1_0__f_clk/a_110_47# 0.0022f
C59234 _0752_/a_300_297# clknet_1_0__leaf__0460_ 0.00204f
C59235 _1057_/a_634_159# VPWR 0.17827f
C59236 comp0.B\[4\] _1034_/a_381_47# 0
C59237 _1048_/a_634_159# _0186_ 0
C59238 _0233_ _0345_ 0.09397f
C59239 _0343_ _0377_ 0.00232f
C59240 _0663_/a_27_413# _0422_ 0
C59241 _0663_/a_207_413# net217 0
C59242 _0647_/a_129_47# _0404_ 0
C59243 net169 VPWR 0.3262f
C59244 net76 clknet_0__0465_ 0.00327f
C59245 _0274_ _0257_ 0.02258f
C59246 net44 _0398_ 0
C59247 clknet_1_0__leaf__0462_ acc0.A\[25\] 0.12003f
C59248 _0315_ _1007_/a_27_47# 0
C59249 _0366_ _1007_/a_193_47# 0.30317f
C59250 _0174_ _0548_/a_240_47# 0.01223f
C59251 clkbuf_1_1__f__0459_/a_110_47# _0300_ 0.00536f
C59252 _0155_ _0511_/a_81_21# 0
C59253 net124 VPWR 0.36388f
C59254 net125 _0138_ 0.00945f
C59255 _0476_ _0949_/a_59_75# 0
C59256 hold5/a_49_47# net152 0
C59257 _0335_ _0220_ 0
C59258 _0992_/a_193_47# _0181_ 0
C59259 pp[7] net63 0.00438f
C59260 net11 net12 0.00255f
C59261 net45 hold59/a_285_47# 0
C59262 pp[6] _0621_/a_35_297# 0
C59263 _0522_/a_27_297# _0522_/a_109_297# 0.17136f
C59264 acc0.A\[7\] net75 0.04063f
C59265 _1050_/a_193_47# clknet_1_1__leaf__0464_ 0
C59266 net35 net164 0
C59267 _0989_/a_1059_315# net75 0
C59268 _1017_/a_193_47# _0240_ 0
C59269 _1067_/a_561_413# _0460_ 0
C59270 _1067_/a_592_47# clknet_1_0__leaf__0457_ 0
C59271 _0967_/a_297_297# _0468_ 0
C59272 _0162_ _0468_ 0
C59273 _0690_/a_150_297# _0321_ 0
C59274 _0815_/a_113_297# net66 0
C59275 _1017_/a_193_47# _0369_ 0.02748f
C59276 _0783_/a_215_47# clkbuf_0__0461_/a_110_47# 0
C59277 _0966_/a_109_297# _0479_ 0
C59278 net188 net181 0
C59279 _0981_/a_27_297# _1068_/a_193_47# 0
C59280 clknet_1_1__leaf__0462_ _0738_/a_68_297# 0
C59281 hold101/a_391_47# net62 0
C59282 net185 hold39/a_391_47# 0
C59283 clknet_1_0__leaf__0460_ _0249_ 0.04157f
C59284 _0672_/a_79_21# _0303_ 0.18249f
C59285 _0327_ _0250_ 0.00839f
C59286 _0607_/a_109_297# _0347_ 0.00276f
C59287 _0443_ clkbuf_1_0__f__0465_/a_110_47# 0
C59288 _1059_/a_1059_315# net41 0
C59289 clknet_1_1__leaf__0460_ net52 0.11146f
C59290 _0965_/a_47_47# _0488_ 0.00552f
C59291 hold100/a_285_47# hold18/a_391_47# 0.00309f
C59292 hold100/a_391_47# hold18/a_285_47# 0.00309f
C59293 _0241_ _0240_ 0
C59294 _1020_/a_891_413# net118 0
C59295 _0760_/a_377_297# _0237_ 0
C59296 _0760_/a_129_47# _0381_ 0.00313f
C59297 net178 _0988_/a_193_47# 0.3158f
C59298 _0427_ _0181_ 0.025f
C59299 _0241_ _0369_ 0
C59300 clknet_0__0457_ _0241_ 0
C59301 _0815_/a_113_297# _0991_/a_27_47# 0
C59302 _0343_ hold16/a_391_47# 0.01349f
C59303 _1012_/a_27_47# _0308_ 0.00176f
C59304 _1031_/a_891_413# _1030_/a_891_413# 0
C59305 _0983_/a_193_47# _0399_ 0.15516f
C59306 net51 _1022_/a_27_47# 0.00248f
C59307 _0981_/a_27_297# _0478_ 0.00116f
C59308 _0181_ hold60/a_285_47# 0
C59309 hold58/a_391_47# _0173_ 0.00925f
C59310 _0328_ _0366_ 0.09204f
C59311 clknet_1_0__leaf__0463_ _1061_/a_634_159# 0.00215f
C59312 hold21/a_49_47# acc0.A\[8\] 0
C59313 net34 _0471_ 0.03712f
C59314 acc0.A\[13\] _0219_ 0.28997f
C59315 net234 acc0.A\[18\] 0
C59316 _1011_/a_27_47# hold95/a_49_47# 0
C59317 _0782_/a_27_47# net100 0.00109f
C59318 _1038_/a_193_47# _0172_ 0
C59319 _1038_/a_466_413# net180 0.0013f
C59320 net160 _1037_/a_466_413# 0
C59321 clknet_1_1__leaf__0463_ _0956_/a_32_297# 0.00179f
C59322 _1025_/a_634_159# _1025_/a_592_47# 0
C59323 _0829_/a_109_297# _0829_/a_27_47# 0
C59324 _0243_ _0462_ 0.00265f
C59325 _0764_/a_299_297# clknet_1_0__leaf__0457_ 0
C59326 _0217_ _0869_/a_27_47# 0
C59327 hold5/a_391_47# _1042_/a_193_47# 0.00773f
C59328 VPWR _0494_/a_27_47# 0.29572f
C59329 _0369_ _0973_/a_109_297# 0.0015f
C59330 net69 _0452_ 0
C59331 _0982_/a_634_159# _0195_ 0
C59332 _0982_/a_27_47# _0216_ 0
C59333 clkbuf_0__0463_/a_110_47# _0463_ 0.3972f
C59334 _1055_/a_561_413# _0181_ 0
C59335 clknet_0__0463_ control0.reset 0.12118f
C59336 acc0.A\[12\] pp[8] 0
C59337 acc0.A\[4\] net170 0
C59338 clkbuf_0_clk/a_110_47# _0972_/a_93_21# 0
C59339 _0118_ _0181_ 0
C59340 acc0.A\[12\] _0664_/a_79_21# 0.01554f
C59341 _0924_/a_27_47# net157 0.00687f
C59342 VPWR clkbuf_1_1__f__0465_/a_110_47# 1.32568f
C59343 clknet_1_1__leaf__0459_ _0808_/a_266_47# 0.00771f
C59344 _1046_/a_1017_47# net10 0
C59345 comp0.B\[6\] _0564_/a_68_297# 0
C59346 comp0.B\[5\] _0564_/a_150_297# 0
C59347 acc0.A\[11\] net79 0
C59348 _0653_/a_113_47# _0417_ 0
C59349 _0982_/a_466_413# _0856_/a_215_47# 0
C59350 hold17/a_285_47# control0.count\[2\] 0.08407f
C59351 _0403_ _0994_/a_1059_315# 0
C59352 _1021_/a_381_47# _1067_/a_1059_315# 0
C59353 _0533_/a_373_47# comp0.B\[15\] 0
C59354 hold86/a_49_47# _0449_ 0
C59355 net31 comp0.B\[9\] 0.28593f
C59356 acc0.A\[14\] _0670_/a_79_21# 0.15641f
C59357 acc0.A\[0\] net47 0.00103f
C59358 _0539_/a_68_297# net195 0
C59359 _0399_ _0526_/a_27_47# 0
C59360 _0996_/a_891_413# _0996_/a_975_413# 0.00851f
C59361 _0996_/a_381_47# _0996_/a_561_413# 0.00123f
C59362 _1055_/a_1059_315# _0517_/a_299_297# 0
C59363 hold59/a_391_47# net104 0.01664f
C59364 _0812_/a_79_21# hold70/a_285_47# 0
C59365 net134 net147 0
C59366 hold57/a_285_47# _0173_ 0.05905f
C59367 _0386_ _0352_ 0.10293f
C59368 _0314_ _1025_/a_27_47# 0
C59369 _0174_ net7 0.36788f
C59370 _0218_ _0771_/a_27_413# 0.00609f
C59371 _0473_ _0138_ 0.0294f
C59372 _0753_/a_465_47# acc0.A\[23\] 0
C59373 _0129_ _0708_/a_150_297# 0
C59374 _0849_/a_297_297# _0350_ 0
C59375 comp0.B\[1\] _0180_ 0
C59376 _0465_ clknet_1_1__leaf__0457_ 0.1843f
C59377 clknet_1_0__leaf__0464_ _1048_/a_975_413# 0
C59378 hold53/a_391_47# net210 0
C59379 _0518_/a_109_47# _0369_ 0
C59380 _0404_ clkbuf_1_1__f__0459_/a_110_47# 0
C59381 input16/a_75_212# A[9] 0.21531f
C59382 _0375_ _0219_ 0.02181f
C59383 _0376_ _0377_ 0.36618f
C59384 net146 _0505_/a_27_297# 0.07124f
C59385 _1052_/a_193_47# clknet_1_1__leaf__0458_ 0
C59386 acc0.A\[16\] _1016_/a_27_47# 0.01465f
C59387 net36 _0209_ 0
C59388 _0714_/a_512_297# _0341_ 0.00264f
C59389 _0698_/a_199_47# _0318_ 0
C59390 hold42/a_391_47# clknet_1_1__leaf__0465_ 0.0083f
C59391 hold70/a_391_47# net228 0.07156f
C59392 clknet_1_0__leaf__0463_ _1039_/a_634_159# 0
C59393 _0701_/a_209_47# clknet_1_1__leaf__0462_ 0
C59394 VPWR _1036_/a_1059_315# 0.40146f
C59395 _1057_/a_891_413# clknet_1_1__leaf__0465_ 0.03553f
C59396 acc0.A\[2\] clknet_1_1__leaf__0457_ 0
C59397 hold27/a_285_47# net8 0
C59398 clknet_0__0457_ _0982_/a_193_47# 0.00127f
C59399 _0536_/a_51_297# net173 0
C59400 _1044_/a_634_159# _1044_/a_466_413# 0.23992f
C59401 _1044_/a_193_47# _1044_/a_1059_315# 0.03405f
C59402 _1044_/a_27_47# _1044_/a_891_413# 0.03224f
C59403 _0596_/a_59_75# acc0.A\[21\] 0.10154f
C59404 _0355_ acc0.A\[29\] 0.05234f
C59405 _0274_ _0640_/a_392_297# 0
C59406 hold46/a_49_47# _0954_/a_32_297# 0.00177f
C59407 hold11/a_391_47# _0536_/a_51_297# 0.01217f
C59408 _0149_ _1044_/a_193_47# 0
C59409 comp0.B\[7\] comp0.B\[10\] 0.00399f
C59410 _0966_/a_27_47# VPWR 0.00611f
C59411 hold52/a_391_47# _0575_/a_27_297# 0
C59412 hold52/a_285_47# _0575_/a_109_297# 0
C59413 _1056_/a_193_47# net16 0
C59414 hold65/a_391_47# _0087_ 0
C59415 net131 _1044_/a_1059_315# 0
C59416 _0217_ _0633_/a_109_297# 0.00388f
C59417 hold59/a_49_47# net234 0
C59418 _0149_ net131 0
C59419 _0244_ _0774_/a_68_297# 0.06053f
C59420 _0580_/a_27_297# clknet_1_0__leaf__0461_ 0.00831f
C59421 VPWR _0777_/a_285_47# 0.00814f
C59422 _0803_/a_150_297# VPWR 0.00351f
C59423 _0357_ clkbuf_1_1__f__0460_/a_110_47# 0.01803f
C59424 _0802_/a_59_75# _0298_ 0
C59425 hold56/a_285_47# net202 0
C59426 clknet_1_1__leaf__0459_ _0345_ 0.50319f
C59427 _1067_/a_27_47# net17 0.03684f
C59428 net46 _1023_/a_466_413# 0.00305f
C59429 net56 _0726_/a_240_47# 0
C59430 clknet_1_1__leaf__0458_ net12 0
C59431 hold56/a_285_47# clknet_1_1__leaf__0463_ 0.00242f
C59432 _1051_/a_1059_315# _0196_ 0
C59433 _0399_ _0793_/a_240_47# 0
C59434 _0789_/a_315_47# VPWR 0.00311f
C59435 _0440_ _0252_ 0.00382f
C59436 net194 clknet_1_1__leaf__0464_ 0.81535f
C59437 _0259_ _0627_/a_215_53# 0.10255f
C59438 VPWR _0754_/a_51_297# 0.5134f
C59439 _0181_ net142 0.02522f
C59440 net245 _0219_ 0.13388f
C59441 net70 _0158_ 0
C59442 hold54/a_49_47# net106 0
C59443 _0359_ _0321_ 0
C59444 _0324_ _0360_ 0.10767f
C59445 _0369_ _0410_ 0.01294f
C59446 net146 _0506_/a_81_21# 0
C59447 _0233_ net52 0
C59448 _0432_ clkbuf_0__0465_/a_110_47# 0.00673f
C59449 clkbuf_0__0460_/a_110_47# _0359_ 0.03327f
C59450 net125 net134 0
C59451 clknet_1_1__leaf__0460_ _0394_ 0.00178f
C59452 _1003_/a_592_47# _0467_ 0
C59453 _0575_/a_109_297# net52 0.00406f
C59454 VPWR _0673_/a_253_47# 0.00278f
C59455 _0464_ VPWR 0.78503f
C59456 VPWR _0672_/a_510_47# 0
C59457 _0369_ net62 0.02695f
C59458 _0627_/a_369_297# clknet_1_1__leaf__0458_ 0
C59459 acc0.A\[4\] _0525_/a_81_21# 0
C59460 _0259_ _0817_/a_266_297# 0
C59461 _0849_/a_215_47# _0849_/a_510_47# 0.00529f
C59462 _0458_ clkbuf_0__0458_/a_110_47# 0.31441f
C59463 clknet_1_0__leaf__0463_ _1040_/a_1017_47# 0
C59464 hold101/a_49_47# _0987_/a_1059_315# 0
C59465 _1032_/a_891_413# _1032_/a_1017_47# 0.00617f
C59466 _1032_/a_193_47# net202 0.23108f
C59467 _0758_/a_79_21# _0103_ 0
C59468 _0568_/a_27_297# _0128_ 0.12484f
C59469 _0568_/a_373_47# net208 0.00122f
C59470 _0429_ pp[5] 0
C59471 _0288_ _0508_/a_384_47# 0
C59472 _0982_/a_27_47# net247 0
C59473 _1032_/a_193_47# clknet_1_1__leaf__0463_ 0.01244f
C59474 _0569_/a_27_297# acc0.A\[29\] 0.13759f
C59475 _0177_ _0492_/a_27_47# 0.00522f
C59476 _0374_ hold94/a_285_47# 0.09824f
C59477 _0578_/a_109_297# _0721_/a_27_47# 0
C59478 _0230_ _0222_ 0.36688f
C59479 _0231_ clknet_1_0__leaf__0460_ 0.06416f
C59480 clknet_0__0460_ _0686_/a_219_297# 0.01206f
C59481 _1051_/a_561_413# _0180_ 0.0015f
C59482 hold46/a_285_47# _0540_/a_51_297# 0
C59483 net27 net28 0
C59484 _0852_/a_285_297# _0446_ 0
C59485 _1014_/a_1017_47# net149 0.00166f
C59486 _1014_/a_891_413# _0112_ 0
C59487 hold39/a_285_47# _0161_ 0
C59488 net247 _0145_ 0.07715f
C59489 _0310_ _0614_/a_111_297# 0
C59490 net33 _1066_/a_975_413# 0
C59491 net211 net46 0.00269f
C59492 hold44/a_285_47# VPWR 0.28638f
C59493 _0328_ _0689_/a_68_297# 0.00118f
C59494 _0765_/a_297_297# _0352_ 0
C59495 net1 clknet_1_0__leaf__0460_ 0.02998f
C59496 _0367_ _0460_ 0
C59497 _0343_ _1055_/a_634_159# 0
C59498 acc0.A\[27\] _1028_/a_193_47# 0.0392f
C59499 comp0.B\[14\] _0954_/a_32_297# 0.13852f
C59500 _0535_/a_68_297# comp0.B\[11\] 0
C59501 _0646_/a_47_47# VPWR 0.32953f
C59502 hold25/a_285_47# _0206_ 0
C59503 hold25/a_391_47# comp0.B\[8\] 0
C59504 _0292_ _0345_ 0.03496f
C59505 _0292_ _0814_/a_27_47# 0.01668f
C59506 clknet_1_0__leaf__0465_ net130 0.01757f
C59507 net45 _0219_ 0.08934f
C59508 hold27/a_285_47# net10 0
C59509 net163 _1030_/a_193_47# 0.0025f
C59510 _0818_/a_193_47# _0181_ 0
C59511 net202 _0721_/a_27_47# 0.00107f
C59512 _0287_ _0295_ 0.50318f
C59513 _0289_ _0304_ 0.00137f
C59514 net168 _1052_/a_466_413# 0
C59515 _0376_ net109 0
C59516 _0234_ acc0.A\[23\] 0
C59517 _0227_ _0369_ 0
C59518 _0140_ hold51/a_285_47# 0
C59519 _0352_ _1006_/a_466_413# 0.00608f
C59520 _0229_ _0103_ 0
C59521 pp[1] _0988_/a_634_159# 0
C59522 _0455_ _0451_ 0
C59523 VPWR _0995_/a_381_47# 0.07676f
C59524 net101 _1015_/a_27_47# 0.22622f
C59525 _0284_ _0993_/a_466_413# 0.00222f
C59526 _0349_ net116 0
C59527 _0216_ _0245_ 0
C59528 net247 _0446_ 0
C59529 net70 acc0.A\[14\] 0
C59530 net192 net4 0.0506f
C59531 _0719_/a_27_47# _0217_ 0
C59532 _1051_/a_634_159# _0525_/a_299_297# 0
C59533 net71 acc0.A\[3\] 0.02123f
C59534 _0216_ _0747_/a_297_297# 0.00247f
C59535 _0183_ clknet_1_0__leaf__0457_ 0.65979f
C59536 _0217_ _0460_ 0.03865f
C59537 _0550_/a_51_297# _0137_ 0.19315f
C59538 _0550_/a_240_47# net180 0.04404f
C59539 _0550_/a_512_297# _0172_ 0
C59540 _0104_ _1006_/a_381_47# 0.13261f
C59541 clknet_1_0__leaf__0458_ _0534_/a_81_21# 0
C59542 _0126_ _1008_/a_466_413# 0
C59543 _0432_ _0824_/a_59_75# 0.11025f
C59544 _0109_ _0725_/a_80_21# 0
C59545 _0951_/a_109_93# _1062_/a_27_47# 0
C59546 acc0.A\[24\] _1007_/a_193_47# 0.00645f
C59547 hold71/a_285_47# hold71/a_391_47# 0.41909f
C59548 _0174_ comp0.B\[11\] 0.02818f
C59549 _0723_/a_27_413# _0334_ 0.11523f
C59550 hold64/a_49_47# _0241_ 0.00103f
C59551 hold14/a_391_47# _0211_ 0.02884f
C59552 B[12] _0542_/a_51_297# 0
C59553 _1000_/a_561_413# _0461_ 0
C59554 hold53/a_49_47# _1024_/a_27_47# 0
C59555 output66/a_27_47# hold34/a_391_47# 0.00122f
C59556 _0762_/a_79_21# hold3/a_49_47# 0.00484f
C59557 _0274_ clknet_1_1__leaf__0458_ 0.17942f
C59558 _0294_ net6 0
C59559 _0136_ net28 0
C59560 net168 _0194_ 0
C59561 clknet_1_0__leaf__0462_ _0103_ 0
C59562 hold33/a_49_47# comp0.B\[10\] 0.00378f
C59563 hold45/a_285_47# acc0.A\[11\] 0.04695f
C59564 clkbuf_1_0__f__0457_/a_110_47# _0373_ 0
C59565 net55 _0707_/a_75_199# 0
C59566 _0216_ hold9/a_285_47# 0
C59567 _0664_/a_79_21# net42 0
C59568 _0346_ clkbuf_1_0__f__0460_/a_110_47# 0
C59569 _0546_/a_149_47# _0546_/a_240_47# 0.06872f
C59570 _0546_/a_51_297# _0205_ 0.1958f
C59571 VPWR _1023_/a_1059_315# 0.41252f
C59572 _1047_/a_634_159# clkbuf_1_1__f__0457_/a_110_47# 0.00655f
C59573 hold100/a_285_47# _0846_/a_149_47# 0
C59574 _1036_/a_592_47# _0175_ 0
C59575 hold59/a_285_47# VPWR 0.28476f
C59576 hold38/a_49_47# net23 0
C59577 _0446_ _0844_/a_382_297# 0.01623f
C59578 _0217_ _0457_ 0
C59579 _0991_/a_634_159# _0991_/a_381_47# 0
C59580 comp0.B\[14\] _0540_/a_245_297# 0.0016f
C59581 _0535_/a_68_297# _0202_ 0.00135f
C59582 _0726_/a_240_47# _0345_ 0
C59583 _0726_/a_51_297# _0219_ 0.16469f
C59584 _0858_/a_27_47# _0195_ 0.00284f
C59585 _0837_/a_266_47# clknet_1_1__leaf__0458_ 0
C59586 _0236_ _0763_/a_193_47# 0
C59587 _0346_ _0250_ 0
C59588 net117 net209 0
C59589 _0587_/a_27_47# _0219_ 0.34182f
C59590 comp0.B\[14\] net173 0
C59591 output66/a_27_47# _0510_/a_27_297# 0
C59592 _1041_/a_891_413# net22 0
C59593 _0747_/a_215_47# _0369_ 0.05048f
C59594 _0461_ _0565_/a_245_297# 0
C59595 _0773_/a_285_47# _0392_ 0.00206f
C59596 _0216_ _1029_/a_193_47# 0.03905f
C59597 hold26/a_285_47# net157 0
C59598 net99 _0218_ 0
C59599 _0210_ _0473_ 0
C59600 net233 hold18/a_391_47# 0
C59601 _0234_ _0602_/a_113_47# 0.00939f
C59602 _0982_/a_27_47# net100 0.00205f
C59603 net68 _1014_/a_27_47# 0
C59604 _0793_/a_512_297# _0345_ 0.00137f
C59605 _0736_/a_56_297# _0462_ 0
C59606 _0328_ acc0.A\[24\] 0.20213f
C59607 _0316_ _0360_ 0
C59608 net55 _0321_ 0
C59609 _0195_ net103 0.0241f
C59610 net7 _1046_/a_193_47# 0
C59611 _1001_/a_1059_315# _0183_ 0
C59612 _1001_/a_381_47# _0217_ 0.00504f
C59613 net169 _0523_/a_81_21# 0
C59614 net123 _1037_/a_27_47# 0.23226f
C59615 clknet_1_0__leaf__0462_ net210 0.04253f
C59616 control0.state\[1\] _0948_/a_109_297# 0
C59617 _0249_ hold94/a_285_47# 0
C59618 _0399_ _0996_/a_891_413# 0.03121f
C59619 output50/a_27_47# net50 0.17648f
C59620 _0574_/a_373_47# acc0.A\[25\] 0.00122f
C59621 net166 clknet_0__0461_ 0
C59622 _0984_/a_27_47# _0268_ 0
C59623 comp0.B\[4\] comp0.B\[2\] 0.03974f
C59624 _0800_/a_51_297# _0300_ 0
C59625 clknet_0__0459_ _0304_ 0
C59626 _0226_ _0762_/a_215_47# 0
C59627 _0598_/a_382_297# _0383_ 0
C59628 _0808_/a_368_297# _0418_ 0.01544f
C59629 net79 _0281_ 0
C59630 _0808_/a_585_47# _0281_ 0.00107f
C59631 input26/a_75_212# control0.sh 0
C59632 _1021_/a_193_47# _0183_ 0.03614f
C59633 _1021_/a_1059_315# net150 0.03061f
C59634 _1021_/a_466_413# _0217_ 0.00345f
C59635 _0548_/a_240_47# comp0.B\[9\] 0.03377f
C59636 _1041_/a_891_413# clknet_1_0__leaf__0463_ 0
C59637 _0347_ _0360_ 0
C59638 _0947_/a_109_297# net35 0.00114f
C59639 _0174_ _0202_ 0.2759f
C59640 clknet_0__0458_ _0642_/a_298_297# 0
C59641 _0222_ _0236_ 0
C59642 _1058_/a_891_413# acc0.A\[10\] 0.03726f
C59643 _0391_ _0771_/a_298_297# 0.03921f
C59644 _0099_ _0771_/a_27_413# 0
C59645 clknet_1_0__leaf__0465_ _0525_/a_299_297# 0.00903f
C59646 _0218_ _0841_/a_510_47# 0
C59647 _0234_ _1003_/a_891_413# 0
C59648 _0546_/a_51_297# _1042_/a_193_47# 0
C59649 _0522_/a_373_47# net13 0
C59650 _0522_/a_109_297# _0193_ 0.00169f
C59651 _0803_/a_68_297# _0286_ 0
C59652 _0800_/a_245_297# _0413_ 0.00109f
C59653 _0461_ _1018_/a_1059_315# 0
C59654 _0456_ _0345_ 0.28988f
C59655 net22 net147 0.00153f
C59656 output66/a_27_47# _0181_ 0.00183f
C59657 _0224_ net109 0.04484f
C59658 _0655_/a_215_53# _0345_ 0.01943f
C59659 net201 _0563_/a_245_297# 0
C59660 _0170_ _1068_/a_193_47# 0
C59661 net167 _1068_/a_1059_315# 0.00143f
C59662 VPWR _0830_/a_79_21# 0.43899f
C59663 hold86/a_49_47# _0260_ 0
C59664 net61 _0628_/a_109_297# 0
C59665 VPWR input33/a_75_212# 0.26739f
C59666 VPWR _1031_/a_381_47# 0.0761f
C59667 _0504_/a_27_47# hold2/a_49_47# 0.005f
C59668 _0304_ _0655_/a_109_93# 0
C59669 _0673_/a_253_47# _0283_ 0
C59670 clknet_0__0465_ _0986_/a_193_47# 0.0104f
C59671 clkbuf_0__0465_/a_110_47# _0986_/a_381_47# 0.00119f
C59672 net126 net31 0
C59673 _0195_ _1019_/a_1059_315# 0
C59674 net46 net241 0
C59675 _0635_/a_27_47# acc0.A\[15\] 0.00368f
C59676 acc0.A\[12\] _0648_/a_109_297# 0
C59677 _0449_ _0823_/a_109_297# 0
C59678 _0289_ _0811_/a_384_47# 0
C59679 _0401_ _0991_/a_891_413# 0
C59680 _0425_ _0991_/a_1059_315# 0
C59681 clknet_1_1__leaf__0459_ _0791_/a_113_297# 0
C59682 _0719_/a_27_47# _0248_ 0.00481f
C59683 _0172_ net29 0
C59684 _0572_/a_27_297# _1025_/a_27_47# 0
C59685 _1043_/a_193_47# hold51/a_391_47# 0
C59686 _0248_ _0460_ 0.04727f
C59687 _0170_ _0478_ 0.00183f
C59688 _1020_/a_27_47# VPWR 0.65029f
C59689 clkbuf_1_1__f__0462_/a_110_47# _0729_/a_68_297# 0
C59690 _0785_/a_299_297# _0345_ 0
C59691 clknet_1_0__leaf__0463_ net147 0.08219f
C59692 _0820_/a_297_297# VPWR 0.00738f
C59693 _0305_ _0459_ 0.02492f
C59694 _0596_/a_145_75# net49 0.00123f
C59695 _0971_/a_299_297# _1063_/a_27_47# 0
C59696 _0971_/a_81_21# _1063_/a_193_47# 0.0015f
C59697 hold41/a_391_47# output67/a_27_47# 0
C59698 _0534_/a_299_297# _0532_/a_81_21# 0
C59699 _0183_ _0850_/a_68_297# 0
C59700 VPWR _0589_/a_113_47# 0
C59701 _0835_/a_78_199# _0255_ 0.07506f
C59702 pp[12] net6 0
C59703 _0238_ _0232_ 0.00415f
C59704 net124 net30 0
C59705 _0829_/a_27_47# _0827_/a_27_47# 0.00289f
C59706 _0264_ _0350_ 0.02916f
C59707 _0150_ _0522_/a_27_297# 0.08687f
C59708 net160 _0135_ 0
C59709 _0251_ hold65/a_285_47# 0.00455f
C59710 _1025_/a_891_413# acc0.A\[25\] 0.0469f
C59711 _0292_ _0819_/a_81_21# 0
C59712 net5 _0301_ 0
C59713 _1020_/a_27_47# _1015_/a_466_413# 0.00151f
C59714 _0984_/a_1017_47# _0347_ 0
C59715 _0971_/a_384_47# clknet_1_0__leaf__0457_ 0
C59716 _0971_/a_81_21# _0460_ 0.00107f
C59717 _0165_ _1067_/a_27_47# 0.12416f
C59718 hold5/a_285_47# net128 0
C59719 net68 _0195_ 0
C59720 clknet_1_0__leaf__0457_ hold40/a_285_47# 0.00393f
C59721 net54 _1008_/a_466_413# 0.0014f
C59722 control0.state\[2\] _0974_/a_79_199# 0.05194f
C59723 control0.state\[0\] net23 0
C59724 _0179_ _0988_/a_1059_315# 0
C59725 clkbuf_0_clk/a_110_47# net231 0
C59726 comp0.B\[7\] _0177_ 0
C59727 hold20/a_49_47# _1072_/a_891_413# 0.01135f
C59728 hold20/a_285_47# _1072_/a_1059_315# 0.00197f
C59729 clknet_0__0457_ _1019_/a_466_413# 0.01532f
C59730 clkbuf_1_0__f__0457_/a_110_47# _1019_/a_381_47# 0
C59731 net16 clknet_1_1__leaf__0465_ 0.1165f
C59732 hold97/a_49_47# _0690_/a_68_297# 0.01354f
C59733 _0244_ hold72/a_391_47# 0
C59734 _0559_/a_149_47# comp0.B\[5\] 0
C59735 _0559_/a_51_297# _0474_ 0.00134f
C59736 _0179_ output37/a_27_47# 0
C59737 hold91/a_49_47# net41 0.32845f
C59738 _0164_ _1063_/a_193_47# 0
C59739 _0080_ _0856_/a_215_47# 0.00299f
C59740 net7 comp0.B\[9\] 0.04791f
C59741 _1021_/a_1059_315# control0.add 0
C59742 hold63/a_391_47# _0572_/a_109_297# 0
C59743 _0800_/a_51_297# _0404_ 0.00852f
C59744 _0190_ _0990_/a_1017_47# 0
C59745 B[13] net32 0.0012f
C59746 net55 _1009_/a_27_47# 0.00395f
C59747 _1045_/a_27_47# clknet_1_1__leaf__0464_ 0
C59748 _0275_ net47 0.02416f
C59749 _1036_/a_27_47# _1036_/a_1059_315# 0.04875f
C59750 _1036_/a_193_47# _1036_/a_466_413# 0.08301f
C59751 _0218_ _0396_ 0.10093f
C59752 net217 net37 0
C59753 _1047_/a_891_413# acc0.A\[15\] 0
C59754 _0769_/a_299_297# _0386_ 0.06185f
C59755 _0769_/a_81_21# _0388_ 0
C59756 _0769_/a_384_47# _0244_ 0.00165f
C59757 clknet_1_1__leaf_clk hold84/a_285_47# 0.0092f
C59758 A[11] net37 0.00544f
C59759 hold90/a_49_47# _0319_ 0
C59760 net170 _0350_ 0
C59761 _0183_ hold19/a_285_47# 0
C59762 _0644_/a_47_47# _0644_/a_129_47# 0.00369f
C59763 _0369_ net219 0
C59764 _0225_ clknet_1_0__leaf__0460_ 0.05949f
C59765 net61 net247 0.0011f
C59766 hold68/a_391_47# net215 0.13417f
C59767 _0488_ clknet_0_clk 0
C59768 net146 _0184_ 0.0378f
C59769 clkload0/a_27_47# VPWR 0.46608f
C59770 hold24/a_49_47# _0555_/a_240_47# 0
C59771 hold59/a_285_47# clknet_1_0__leaf__0459_ 0
C59772 _0111_ _0341_ 0.04627f
C59773 hold31/a_285_47# _0273_ 0
C59774 _0176_ _0546_/a_240_47# 0
C59775 clknet_1_0__leaf__0463_ net125 0.31985f
C59776 control0.state\[0\] net35 0
C59777 _1050_/a_193_47# net148 0
C59778 hold54/a_391_47# net8 0
C59779 _0200_ _0138_ 0
C59780 _0403_ _0787_/a_209_47# 0
C59781 _1059_/a_891_413# clkbuf_0__0459_/a_110_47# 0.00708f
C59782 clknet_1_0__leaf__0463_ _0953_/a_220_297# 0
C59783 net44 _0308_ 0.04285f
C59784 _1065_/a_27_47# _0215_ 0
C59785 _1044_/a_466_413# net130 0
C59786 _1065_/a_634_159# _0175_ 0.01293f
C59787 comp0.B\[13\] comp0.B\[11\] 0
C59788 output36/a_27_47# input29/a_75_212# 0.01143f
C59789 hold11/a_49_47# _0144_ 0.31233f
C59790 _0289_ _0813_/a_109_297# 0
C59791 _0606_/a_392_297# _0383_ 0
C59792 _1041_/a_27_47# hold6/a_285_47# 0
C59793 _1038_/a_1017_47# comp0.B\[6\] 0
C59794 net137 net130 0.01609f
C59795 net188 _1058_/a_634_159# 0
C59796 _0744_/a_27_47# net37 0
C59797 VPWR _0776_/a_27_47# 0.01105f
C59798 _0985_/a_891_413# _0465_ 0.00157f
C59799 _0971_/a_299_297# _1062_/a_1059_315# 0
C59800 _0995_/a_193_47# _0297_ 0
C59801 _0804_/a_215_47# net39 0.01613f
C59802 _0137_ _0913_/a_27_47# 0.01235f
C59803 _0138_ comp0.B\[8\] 0.16818f
C59804 _0117_ clknet_1_0__leaf__0461_ 0.00791f
C59805 _0325_ clkbuf_0__0460_/a_110_47# 0
C59806 clknet_1_1__leaf_clk _1065_/a_561_413# 0
C59807 _0777_/a_47_47# _0777_/a_129_47# 0.00369f
C59808 _0410_ _0409_ 0.00102f
C59809 _1049_/a_634_159# _0465_ 0
C59810 net36 _1038_/a_891_413# 0.01693f
C59811 pp[0] _1038_/a_466_413# 0
C59812 _0231_ hold94/a_285_47# 0
C59813 net61 _0825_/a_68_297# 0.00163f
C59814 hold47/a_49_47# _0142_ 0.32382f
C59815 control0.state\[2\] _1062_/a_193_47# 0
C59816 _0985_/a_891_413# acc0.A\[2\] 0
C59817 _0985_/a_1059_315# net58 0
C59818 _0428_ _0990_/a_27_47# 0.00141f
C59819 _0427_ _0990_/a_193_47# 0
C59820 net61 _0844_/a_382_297# 0.00137f
C59821 hold86/a_285_47# _0447_ 0.00125f
C59822 _0467_ _0974_/a_222_93# 0.00158f
C59823 _0237_ _1005_/a_891_413# 0
C59824 _0722_/a_79_21# _0350_ 0.01125f
C59825 _0675_/a_150_297# _0459_ 0
C59826 _0216_ _1028_/a_381_47# 0
C59827 net46 net177 0.06776f
C59828 _0195_ _1028_/a_975_413# 0.00205f
C59829 _0331_ _0109_ 0
C59830 net57 _0723_/a_297_47# 0
C59831 net49 _0383_ 0
C59832 _1057_/a_634_159# _1057_/a_592_47# 0
C59833 VPWR _0219_ 7.027f
C59834 B[13] _1042_/a_1059_315# 0
C59835 _0984_/a_466_413# _0991_/a_27_47# 0
C59836 net184 _0148_ 0.00124f
C59837 _0111_ _1013_/a_891_413# 0.00605f
C59838 net59 _0347_ 0
C59839 VPWR _1064_/a_561_413# 0.00237f
C59840 _0413_ _0995_/a_27_47# 0.00155f
C59841 _1059_/a_634_159# _1059_/a_592_47# 0
C59842 _0789_/a_75_199# _0789_/a_315_47# 0.02023f
C59843 VPWR _0669_/a_111_297# 0
C59844 VPWR _0728_/a_59_75# 0.20781f
C59845 hold13/a_391_47# net160 0.13101f
C59846 hold13/a_285_47# _0210_ 0.00199f
C59847 hold76/a_49_47# net45 0.02778f
C59848 hold19/a_285_47# acc0.A\[15\] 0
C59849 hold41/a_49_47# _0186_ 0.01939f
C59850 net243 _0123_ 0
C59851 _1015_/a_561_413# _0345_ 0
C59852 hold23/a_49_47# _0195_ 0.00115f
C59853 _0981_/a_27_297# VPWR 0.20855f
C59854 _0433_ _0989_/a_27_47# 0
C59855 _0433_ hold1/a_49_47# 0.00643f
C59856 _0181_ _1047_/a_193_47# 0.00193f
C59857 _0695_/a_80_21# _0462_ 0.02653f
C59858 B[13] net10 0
C59859 net22 _0473_ 0.02494f
C59860 acc0.A\[29\] _0127_ 0.4087f
C59861 _0238_ clkbuf_0__0460_/a_110_47# 0
C59862 _0673_/a_103_199# _0673_/a_337_297# 0.01015f
C59863 clknet_1_0__leaf__0458_ _0849_/a_510_47# 0.00104f
C59864 _0520_/a_27_297# hold83/a_391_47# 0
C59865 _0520_/a_109_297# hold83/a_285_47# 0
C59866 _1056_/a_27_47# _0428_ 0
C59867 comp0.B\[13\] _0202_ 0.00938f
C59868 _0820_/a_215_47# _0088_ 0
C59869 _0386_ _0392_ 0.13371f
C59870 _0672_/a_79_21# _0672_/a_215_47# 0.04584f
C59871 output43/a_27_47# hold98/a_285_47# 0.0185f
C59872 clknet_1_1__leaf__0459_ _0994_/a_27_47# 0.01042f
C59873 _1030_/a_634_159# clknet_1_1__leaf__0462_ 0
C59874 net193 _0138_ 0
C59875 _0984_/a_466_413# _0350_ 0
C59876 _0349_ _0220_ 0
C59877 net233 _0846_/a_149_47# 0.00671f
C59878 _0343_ net141 0.04669f
C59879 _0715_/a_27_47# _0990_/a_27_47# 0
C59880 _1054_/a_27_47# _0087_ 0
C59881 net132 clknet_1_1__leaf__0464_ 0.09677f
C59882 _0138_ _1046_/a_466_413# 0
C59883 VPWR _1008_/a_634_159# 0.18976f
C59884 _0180_ _0528_/a_384_47# 0
C59885 net158 _1046_/a_634_159# 0
C59886 clknet_1_0__leaf__0463_ _0473_ 0.05156f
C59887 net48 _0219_ 0.16421f
C59888 _0459_ _0181_ 0.05191f
C59889 _0467_ _1062_/a_634_159# 0
C59890 _0144_ _0159_ 0
C59891 _0949_/a_145_75# _0469_ 0
C59892 _1021_/a_27_47# _0467_ 0
C59893 _0124_ _0347_ 0
C59894 _1052_/a_975_413# _0186_ 0
C59895 net190 net113 0.00297f
C59896 _0785_/a_81_21# _0819_/a_299_297# 0
C59897 _0785_/a_299_297# _0819_/a_81_21# 0
C59898 _1058_/a_891_413# _0188_ 0
C59899 clknet_1_0__leaf__0458_ hold71/a_391_47# 0.00463f
C59900 _0388_ clknet_0__0461_ 0
C59901 VPWR _0826_/a_301_297# 0.00138f
C59902 clkbuf_1_1__f__0463_/a_110_47# _0173_ 0.12065f
C59903 _0586_/a_27_47# hold40/a_49_47# 0
C59904 _1056_/a_891_413# net181 0
C59905 _0149_ _0525_/a_81_21# 0.11484f
C59906 comp0.B\[11\] comp0.B\[9\] 0
C59907 acc0.A\[31\] _0218_ 0
C59908 _0172_ _0137_ 0.00948f
C59909 _0182_ net8 0
C59910 _0186_ net75 0
C59911 control0.state\[1\] clkbuf_0_clk/a_110_47# 0.03466f
C59912 pp[27] hold95/a_391_47# 0
C59913 comp0.B\[0\] _1062_/a_634_159# 0
C59914 _0180_ net218 0
C59915 clkbuf_1_1__f__0457_/a_110_47# _0208_ 0
C59916 net200 _1026_/a_27_47# 0
C59917 clknet_0__0463_ _0475_ 0.02092f
C59918 pp[18] hold78/a_49_47# 0.00138f
C59919 _0291_ net67 0
C59920 B[8] _0546_/a_51_297# 0
C59921 hold30/a_49_47# hold96/a_285_47# 0
C59922 control0.state\[1\] _1063_/a_634_159# 0.01592f
C59923 clknet_1_1__leaf__0459_ _0156_ 0
C59924 net207 _1014_/a_193_47# 0
C59925 VPWR hold84/a_391_47# 0.17706f
C59926 _0123_ _1024_/a_381_47# 0
C59927 clknet_1_0__leaf__0462_ _1022_/a_381_47# 0.00304f
C59928 _1005_/a_27_47# _1005_/a_891_413# 0.03224f
C59929 _1005_/a_193_47# _1005_/a_1059_315# 0.03405f
C59930 _1005_/a_634_159# _1005_/a_466_413# 0.23992f
C59931 _0240_ _0352_ 0.22152f
C59932 _0195_ _0774_/a_68_297# 0
C59933 _0235_ _0460_ 0.02487f
C59934 net55 _0338_ 0
C59935 _0950_/a_75_212# _0468_ 0
C59936 _0369_ _0352_ 0.2669f
C59937 VPWR _0511_/a_299_297# 0.24313f
C59938 _0519_/a_81_21# _0519_/a_299_297# 0.08213f
C59939 _1047_/a_975_413# clknet_1_1__leaf__0457_ 0.00108f
C59940 _0984_/a_27_47# net222 0
C59941 _0984_/a_891_413# _0849_/a_215_47# 0
C59942 clknet_0__0457_ _0352_ 0.03164f
C59943 _0222_ _0380_ 0
C59944 _1013_/a_27_47# _1013_/a_634_159# 0.14145f
C59945 _0518_/a_27_297# input15/a_75_212# 0
C59946 _0991_/a_634_159# net67 0
C59947 _0991_/a_381_47# net77 0
C59948 _0991_/a_891_413# _0089_ 0
C59949 acc0.A\[12\] A[10] 0
C59950 VPWR _0746_/a_81_21# 0.23934f
C59951 _0356_ net57 0
C59952 _0300_ _0277_ 0.78471f
C59953 net185 hold38/a_285_47# 0.00795f
C59954 _0415_ _0993_/a_466_413# 0
C59955 _0181_ _0265_ 0.0245f
C59956 _0212_ hold38/a_49_47# 0
C59957 hold96/a_285_47# _0352_ 0
C59958 hold96/a_49_47# _0102_ 0.0049f
C59959 _1000_/a_1059_315# clknet_1_0__leaf__0461_ 0.00132f
C59960 _0607_/a_27_297# _0607_/a_109_47# 0.00393f
C59961 _0399_ _0255_ 0.00156f
C59962 _0985_/a_466_413# _0261_ 0.00444f
C59963 _0985_/a_1059_315# _0262_ 0
C59964 clknet_1_1__leaf__0459_ _0997_/a_193_47# 0.02627f
C59965 _0195_ net191 0.00104f
C59966 _0574_/a_27_297# _0216_ 0.26524f
C59967 _0646_/a_47_47# _0995_/a_634_159# 0
C59968 _0499_/a_59_75# acc0.A\[15\] 0
C59969 _0238_ _1009_/a_27_47# 0
C59970 clknet_1_1__leaf__0459_ _0992_/a_891_413# 0.01709f
C59971 acc0.A\[8\] acc0.A\[9\] 0
C59972 _0248_ _0614_/a_29_53# 0
C59973 _0274_ _0642_/a_27_413# 0.00133f
C59974 hold31/a_285_47# _0086_ 0.00231f
C59975 net245 _0997_/a_891_413# 0
C59976 _0095_ _0345_ 0.00433f
C59977 _0982_/a_561_413# acc0.A\[0\] 0
C59978 _1038_/a_27_47# _1040_/a_634_159# 0
C59979 _1038_/a_634_159# _1040_/a_27_47# 0
C59980 _1004_/a_1017_47# acc0.A\[23\] 0
C59981 VPWR _1065_/a_975_413# 0.00439f
C59982 _1012_/a_27_47# hold92/a_391_47# 0
C59983 _1012_/a_193_47# hold92/a_285_47# 0
C59984 _0600_/a_103_199# _0223_ 0.09805f
C59985 _0260_ _0823_/a_109_297# 0.00174f
C59986 _1018_/a_1059_315# _0582_/a_27_297# 0
C59987 comp0.B\[10\] _0203_ 0
C59988 net138 _0186_ 0.02841f
C59989 _1056_/a_193_47# net142 0.00378f
C59990 comp0.B\[9\] _0202_ 0
C59991 _0995_/a_634_159# _0995_/a_381_47# 0
C59992 _0093_ _0297_ 0
C59993 _0119_ _0217_ 0.15911f
C59994 _0211_ net25 0
C59995 net62 _0084_ 0.2221f
C59996 _1060_/a_1017_47# acc0.A\[15\] 0
C59997 _0983_/a_193_47# _0346_ 0
C59998 _1002_/a_891_413# _0382_ 0.00167f
C59999 net59 hold95/a_49_47# 0
C60000 input6/a_75_212# _0668_/a_79_21# 0
C60001 clknet_1_0__leaf__0459_ _0219_ 0.60431f
C60002 _1034_/a_1059_315# _0561_/a_51_297# 0.00139f
C60003 _0436_ _0434_ 0
C60004 _1050_/a_891_413# _0142_ 0
C60005 clknet_0_clk _1065_/a_193_47# 0.01057f
C60006 net32 _1042_/a_634_159# 0.01646f
C60007 net152 _1042_/a_466_413# 0
C60008 net165 _0635_/a_109_297# 0.00113f
C60009 _1018_/a_27_47# _0459_ 0.00335f
C60010 _0123_ _0366_ 0
C60011 hold85/a_49_47# control0.state\[2\] 0
C60012 hold57/a_285_47# net204 0.00983f
C60013 hold45/a_285_47# A[12] 0
C60014 _0287_ _0346_ 0.71239f
C60015 control0.state\[0\] _1062_/a_561_413# 0
C60016 _0412_ _0093_ 0
C60017 _0982_/a_634_159# _0183_ 0.01579f
C60018 _0982_/a_1059_315# _0217_ 0
C60019 _1034_/a_634_159# _0473_ 0
C60020 _0361_ _0328_ 0.0214f
C60021 _0783_/a_79_21# _0219_ 0.00475f
C60022 hold74/a_391_47# _0115_ 0
C60023 pp[28] hold95/a_285_47# 0
C60024 _0401_ hold70/a_391_47# 0
C60025 hold25/a_285_47# A[1] 0
C60026 _0303_ _0301_ 0.12572f
C60027 _0704_/a_68_297# net209 0
C60028 acc0.A\[30\] hold62/a_285_47# 0
C60029 _0182_ net10 0
C60030 _1011_/a_634_159# _1011_/a_592_47# 0
C60031 _1016_/a_975_413# _0369_ 0
C60032 _0133_ _1034_/a_1059_315# 0
C60033 hold96/a_49_47# _0574_/a_109_47# 0
C60034 hold29/a_391_47# acc0.A\[23\] 0.02834f
C60035 _1006_/a_27_47# _1006_/a_193_47# 0.96639f
C60036 net126 net7 0
C60037 clkload2/a_268_47# net170 0
C60038 _0350_ _1006_/a_1017_47# 0.00163f
C60039 _0216_ net105 0.02315f
C60040 net45 _0997_/a_891_413# 0
C60041 _0972_/a_93_21# _0487_ 0.08551f
C60042 _0257_ _0433_ 0.08278f
C60043 _0275_ _0294_ 0.00438f
C60044 _0274_ _0218_ 0
C60045 _0751_/a_29_53# _0751_/a_111_297# 0.005f
C60046 _0216_ _0326_ 0
C60047 _0290_ net67 0.02011f
C60048 hold14/a_391_47# clknet_1_0__leaf__0463_ 0
C60049 _0856_/a_79_21# _0350_ 0.00612f
C60050 _0124_ _1025_/a_27_47# 0
C60051 _1030_/a_193_47# net116 0.01325f
C60052 _1055_/a_1059_315# VPWR 0.40088f
C60053 _1056_/a_592_47# clknet_1_1__leaf__0465_ 0
C60054 net196 hold51/a_49_47# 0
C60055 _1018_/a_193_47# clknet_1_0__leaf__0461_ 0.0415f
C60056 _0102_ net90 0.02419f
C60057 _0350_ _0986_/a_1017_47# 0
C60058 _0453_ _0219_ 0
C60059 _1001_/a_466_413# acc0.A\[19\] 0
C60060 _0577_/a_109_297# net49 0.00156f
C60061 _0352_ _1024_/a_27_47# 0
C60062 _1003_/a_466_413# VPWR 0.27093f
C60063 _0429_ _0828_/a_113_297# 0.15454f
C60064 net9 _0527_/a_109_297# 0.00191f
C60065 hold52/a_391_47# net176 0
C60066 _0346_ net9 0
C60067 net35 _1068_/a_193_47# 0
C60068 _0216_ hold95/a_391_47# 0.00107f
C60069 _0959_/a_80_21# _0163_ 0
C60070 _0986_/a_27_47# _0986_/a_193_47# 0.96469f
C60071 net77 _0082_ 0
C60072 _0585_/a_109_297# _0181_ 0.02261f
C60073 _0404_ _0277_ 0.43287f
C60074 _0298_ _0300_ 0.38896f
C60075 _0311_ _0294_ 0.77296f
C60076 _0150_ _0193_ 0.01697f
C60077 net148 _0987_/a_193_47# 0.0179f
C60078 _0442_ _0186_ 0
C60079 net33 clknet_0_clk 0
C60080 _0225_ hold94/a_285_47# 0.00822f
C60081 clknet_1_1__leaf__0459_ _0411_ 0.01383f
C60082 acc0.A\[7\] _0436_ 0
C60083 _0435_ _0989_/a_891_413# 0.00235f
C60084 net64 acc0.A\[9\] 0
C60085 _0436_ _0989_/a_1059_315# 0
C60086 _1020_/a_27_47# _0113_ 0
C60087 _0118_ _1015_/a_27_47# 0
C60088 _1023_/a_193_47# _1023_/a_466_413# 0.07874f
C60089 _1023_/a_27_47# _1023_/a_1059_315# 0.04875f
C60090 VPWR _0799_/a_209_297# 0.20308f
C60091 clknet_1_0__leaf__0463_ _0497_/a_68_297# 0.00227f
C60092 _1042_/a_634_159# _1042_/a_1059_315# 0
C60093 _1042_/a_27_47# _1042_/a_381_47# 0.05761f
C60094 _1042_/a_193_47# _1042_/a_891_413# 0.19226f
C60095 hold100/a_285_47# acc0.A\[15\] 0.01798f
C60096 _0181_ _1060_/a_381_47# 0.01297f
C60097 net46 _0461_ 0.01256f
C60098 control0.add net223 0
C60099 hold85/a_285_47# _0467_ 0
C60100 _0175_ _0563_/a_240_47# 0
C60101 hold12/a_391_47# clknet_0_clk 0.00169f
C60102 clknet_0__0457_ net207 0.05013f
C60103 _1010_/a_592_47# _0347_ 0.00107f
C60104 _0423_ acc0.A\[9\] 0.29737f
C60105 _0982_/a_634_159# acc0.A\[15\] 0
C60106 _0459_ _0507_/a_373_47# 0
C60107 VPWR hold61/a_49_47# 0.32141f
C60108 _1017_/a_27_47# _0307_ 0
C60109 net9 _1061_/a_193_47# 0
C60110 _0179_ _1050_/a_466_413# 0.01138f
C60111 _0413_ _0299_ 0
C60112 _0800_/a_149_47# _0219_ 0.00951f
C60113 _0347_ _0841_/a_215_47# 0.06279f
C60114 _0825_/a_68_297# _0431_ 0
C60115 clkbuf_1_1__f__0465_/a_110_47# _0345_ 0.00176f
C60116 clkbuf_1_1__f__0465_/a_110_47# _0814_/a_27_47# 0
C60117 _0470_ _0164_ 0
C60118 _0458_ _0447_ 0.27088f
C60119 _0714_/a_240_47# _0339_ 0.00124f
C60120 _1036_/a_891_413# _1036_/a_1017_47# 0.00617f
C60121 _1036_/a_193_47# net161 0.25551f
C60122 net158 _1045_/a_27_47# 0
C60123 hold69/a_391_47# net52 0.05958f
C60124 net10 _1042_/a_634_159# 0.00141f
C60125 _0153_ _0988_/a_193_47# 0
C60126 _0480_ _0162_ 0.00103f
C60127 hold76/a_49_47# VPWR 0.28565f
C60128 _0343_ _0831_/a_35_297# 0
C60129 VPWR _1040_/a_1059_315# 0.40528f
C60130 _0992_/a_193_47# clknet_1_1__leaf__0465_ 0.00129f
C60131 _0218_ _0117_ 0
C60132 hold52/a_285_47# hold68/a_285_47# 0.00214f
C60133 hold27/a_49_47# _0159_ 0
C60134 net163 _0567_/a_27_297# 0
C60135 _0294_ _0583_/a_27_297# 0.02919f
C60136 _1000_/a_27_47# _0241_ 0
C60137 _0997_/a_193_47# _0793_/a_512_297# 0
C60138 _0732_/a_80_21# _1007_/a_381_47# 0
C60139 _0181_ _0267_ 0
C60140 _0094_ net42 0
C60141 _0715_/a_27_47# _0293_ 0
C60142 net43 _0218_ 0.78039f
C60143 _0366_ _0758_/a_510_47# 0
C60144 _0741_/a_109_297# _0347_ 0
C60145 control0.reset _0564_/a_150_297# 0
C60146 _1036_/a_193_47# net26 0
C60147 _1011_/a_466_413# _0334_ 0
C60148 hold88/a_285_47# output47/a_27_47# 0
C60149 _0454_ _0350_ 0
C60150 control0.count\[3\] net167 0
C60151 net188 net144 0.0061f
C60152 hold49/a_285_47# _0141_ 0.06884f
C60153 clknet_1_0__leaf__0458_ _0986_/a_193_47# 0
C60154 _0617_/a_150_297# net52 0
C60155 _0271_ _0444_ 0
C60156 clknet_1_0__leaf__0462_ _1024_/a_592_47# 0
C60157 _0467_ _1063_/a_592_47# 0
C60158 _1058_/a_975_413# net4 0
C60159 _0596_/a_59_75# _0381_ 0
C60160 clknet_0__0458_ clkbuf_1_0__f__0465_/a_110_47# 0.00359f
C60161 _1032_/a_193_47# _1067_/a_466_413# 0
C60162 _1032_/a_27_47# _1067_/a_1059_315# 0
C60163 _0195_ hold71/a_49_47# 0.00106f
C60164 _1032_/a_634_159# _1067_/a_634_159# 0
C60165 _1032_/a_1059_315# _1067_/a_27_47# 0
C60166 _1032_/a_466_413# _1067_/a_193_47# 0
C60167 acc0.A\[25\] _0737_/a_35_297# 0
C60168 pp[0] net172 0
C60169 net135 _0465_ 0
C60170 _0368_ _0105_ 0.07707f
C60171 hold68/a_285_47# net52 0
C60172 comp0.B\[11\] hold5/a_285_47# 0.00205f
C60173 net216 _0366_ 0
C60174 _0999_/a_27_47# _0218_ 0.06809f
C60175 _1054_/a_1059_315# acc0.A\[7\] 0.00631f
C60176 _0562_/a_68_297# _0560_/a_68_297# 0.01958f
C60177 _0216_ acc0.A\[28\] 0.05902f
C60178 _0346_ _0655_/a_297_297# 0
C60179 _0179_ hold100/a_285_47# 0
C60180 net190 hold8/a_285_47# 0
C60181 _0363_ _0107_ 0.1051f
C60182 _0803_/a_150_297# _0345_ 0
C60183 clknet_1_0__leaf__0464_ _1049_/a_193_47# 0.02096f
C60184 _0136_ clknet_0__0463_ 0.00323f
C60185 _1058_/a_27_47# acc0.A\[11\] 0.04547f
C60186 _0984_/a_193_47# net77 0
C60187 net70 _0991_/a_193_47# 0
C60188 _0457_ _0565_/a_512_297# 0
C60189 _0736_/a_311_297# _0219_ 0.00113f
C60190 _0279_ _0788_/a_150_297# 0
C60191 _1053_/a_466_413# _1052_/a_634_159# 0
C60192 _1053_/a_27_47# _1052_/a_891_413# 0
C60193 _1053_/a_891_413# _1052_/a_27_47# 0
C60194 clknet_1_1__leaf__0459_ _0809_/a_299_297# 0
C60195 _0289_ _0421_ 0
C60196 hold64/a_49_47# _0352_ 0
C60197 _0217_ _0758_/a_297_297# 0
C60198 _0550_/a_51_297# _1040_/a_466_413# 0
C60199 _0550_/a_149_47# _1040_/a_27_47# 0
C60200 _0216_ net209 0.0022f
C60201 _0357_ clkbuf_1_1__f__0462_/a_110_47# 0
C60202 _0404_ _0298_ 0.71128f
C60203 _0429_ _0433_ 0
C60204 _0789_/a_75_199# _0219_ 0
C60205 _0754_/a_51_297# _0345_ 0.16341f
C60206 _0754_/a_149_47# _0754_/a_240_47# 0.06872f
C60207 _0643_/a_253_47# _0256_ 0
C60208 _0317_ clknet_0__0462_ 0.10117f
C60209 _0734_/a_47_47# _0250_ 0
C60210 _0549_/a_68_297# input29/a_75_212# 0
C60211 _0230_ _0366_ 0
C60212 _0539_/a_68_297# VPWR 0.17472f
C60213 _0459_ clknet_1_1__leaf__0461_ 0.0182f
C60214 _0673_/a_253_47# _0345_ 0.00235f
C60215 net150 _0487_ 0
C60216 _0170_ VPWR 0.44862f
C60217 _0404_ _0296_ 0
C60218 _1055_/a_561_413# clknet_1_1__leaf__0465_ 0
C60219 net234 _0465_ 0
C60220 _0672_/a_510_47# _0345_ 0
C60221 net15 net12 0
C60222 _0462_ clknet_1_0__leaf__0460_ 0.0524f
C60223 _0590_/a_113_47# _0222_ 0.00952f
C60224 _0508_/a_81_21# acc0.A\[15\] 0.00247f
C60225 clkbuf_0_clk/a_110_47# _1068_/a_634_159# 0.00101f
C60226 _0555_/a_149_47# _0210_ 0.00154f
C60227 _0186_ hold83/a_285_47# 0.00176f
C60228 _1038_/a_193_47# _0207_ 0.00213f
C60229 _1002_/a_1059_315# net187 0
C60230 B[1] control0.sh 0
C60231 _0343_ _0719_/a_27_47# 0.00377f
C60232 _0959_/a_80_21# _1066_/a_27_47# 0
C60233 _1051_/a_466_413# _0524_/a_109_297# 0
C60234 net123 _0208_ 0
C60235 _0343_ _0460_ 0.03675f
C60236 B[12] net198 0.00283f
C60237 _0845_/a_193_297# _0845_/a_109_47# 0.0023f
C60238 _0389_ hold76/a_391_47# 0
C60239 _0243_ hold76/a_285_47# 0.01308f
C60240 _0734_/a_129_47# clknet_1_1__leaf__0460_ 0
C60241 _0362_ _0181_ 0.00679f
C60242 _0200_ net22 0.02734f
C60243 VPWR _0994_/a_1059_315# 0.41434f
C60244 _0343_ _1060_/a_193_47# 0.00147f
C60245 _0974_/a_222_93# _1068_/a_381_47# 0
C60246 net159 _1068_/a_27_47# 0.00104f
C60247 VPWR net94 0.38718f
C60248 net77 clkbuf_0__0458_/a_110_47# 0
C60249 _0490_ clkbuf_1_0__f_clk/a_110_47# 0
C60250 _0476_ net205 0.05391f
C60251 net158 net132 0.01691f
C60252 control0.state\[2\] net17 0
C60253 _0226_ net150 0.00204f
C60254 clkbuf_0__0465_/a_110_47# _0841_/a_215_47# 0
C60255 _0327_ acc0.A\[29\] 0.02972f
C60256 _0461_ _1015_/a_1059_315# 0.00158f
C60257 hold5/a_285_47# _0202_ 0
C60258 _1010_/a_634_159# _0350_ 0.04155f
C60259 pp[27] _1011_/a_634_159# 0
C60260 hold75/a_285_47# _0219_ 0.05942f
C60261 _0557_/a_51_297# clknet_1_1__leaf__0463_ 0.00709f
C60262 _0737_/a_35_297# _0737_/a_117_297# 0.00641f
C60263 hold13/a_49_47# _1034_/a_466_413# 0
C60264 net22 comp0.B\[8\] 0
C60265 clknet_0__0457_ net106 0
C60266 net45 _0582_/a_109_297# 0
C60267 _0222_ _1005_/a_891_413# 0
C60268 _0280_ acc0.A\[15\] 0
C60269 _0216_ _0769_/a_81_21# 0.00392f
C60270 _0289_ _0809_/a_81_21# 0.16744f
C60271 _0129_ net208 0
C60272 net144 _0155_ 0.00122f
C60273 net157 _1061_/a_634_159# 0.00723f
C60274 _0846_/a_51_297# _0350_ 0.10338f
C60275 hold70/a_49_47# hold70/a_391_47# 0.00188f
C60276 clknet_1_0__leaf__0463_ _0200_ 0.00103f
C60277 hold63/a_391_47# _1026_/a_27_47# 0
C60278 hold36/a_285_47# _0538_/a_51_297# 0
C60279 _0369_ _0237_ 0.04006f
C60280 _0995_/a_634_159# _0219_ 0
C60281 _0174_ _0544_/a_149_47# 0.02139f
C60282 _0695_/a_80_21# _0312_ 0.19315f
C60283 _0820_/a_510_47# _0399_ 0
C60284 _1009_/a_466_413# _0350_ 0
C60285 _0670_/a_215_47# clkbuf_0__0459_/a_110_47# 0
C60286 _0180_ _0498_/a_51_297# 0
C60287 _0183_ net103 0.00165f
C60288 _1034_/a_27_47# _1033_/a_27_47# 0.07618f
C60289 _1012_/a_27_47# _0336_ 0
C60290 _0269_ net247 0
C60291 _0467_ _0132_ 0
C60292 _0217_ _1016_/a_27_47# 0
C60293 clknet_1_0__leaf__0462_ acc0.A\[22\] 0.11714f
C60294 _0531_/a_27_297# _1047_/a_193_47# 0
C60295 _0531_/a_109_297# _1047_/a_27_47# 0
C60296 _1031_/a_634_159# _1031_/a_381_47# 0
C60297 pp[14] net6 0.00113f
C60298 _0098_ _0459_ 0
C60299 clknet_1_0__leaf__0463_ comp0.B\[8\] 0.11512f
C60300 _0123_ net112 0.00139f
C60301 _0369_ hold72/a_285_47# 0.00936f
C60302 hold30/a_49_47# _0756_/a_47_47# 0
C60303 net55 _0348_ 0
C60304 net31 net32 0
C60305 _0996_/a_891_413# _0346_ 0
C60306 clknet_1_1__leaf__0465_ net142 0.25567f
C60307 comp0.B\[10\] hold6/a_49_47# 0.00139f
C60308 pp[16] net45 0.03371f
C60309 _0121_ net243 0
C60310 control0.state\[0\] _0161_ 0.03259f
C60311 _1000_/a_1059_315# _0218_ 0
C60312 _0179_ _0508_/a_81_21# 0.06404f
C60313 _0722_/a_79_21# _0722_/a_510_47# 0.00844f
C60314 _0722_/a_297_297# _0722_/a_215_47# 0
C60315 _1005_/a_466_413# net91 0
C60316 _1005_/a_634_159# _0103_ 0.0454f
C60317 _0123_ acc0.A\[24\] 0.04353f
C60318 _1059_/a_381_47# _0288_ 0
C60319 hold33/a_49_47# hold27/a_285_47# 0
C60320 _0502_/a_27_47# net36 0
C60321 _0984_/a_975_413# _0082_ 0
C60322 _1060_/a_27_47# net5 0
C60323 _1013_/a_891_413# _1013_/a_975_413# 0.00851f
C60324 _1013_/a_381_47# _1013_/a_561_413# 0.00123f
C60325 _0191_ input15/a_75_212# 0
C60326 net77 net67 0
C60327 _0251_ _0439_ 0
C60328 net1 _1062_/a_634_159# 0
C60329 _1002_/a_466_413# _1002_/a_381_47# 0.03733f
C60330 _1002_/a_193_47# _1002_/a_975_413# 0
C60331 _1002_/a_1059_315# _1002_/a_891_413# 0.31086f
C60332 _1014_/a_27_47# _0264_ 0
C60333 _0251_ VPWR 1.10028f
C60334 net193 net22 0
C60335 _1021_/a_27_47# net1 0.00169f
C60336 clknet_1_0__leaf__0465_ _0524_/a_109_47# 0
C60337 _0640_/a_109_53# VPWR 0.0995f
C60338 _0758_/a_79_21# _0379_ 0.0642f
C60339 _0594_/a_113_47# VPWR 0
C60340 _0984_/a_891_413# clknet_1_0__leaf__0458_ 0.02269f
C60341 _0858_/a_27_47# acc0.A\[15\] 0
C60342 _0248_ _0373_ 0.00401f
C60343 net22 _1046_/a_466_413# 0.00278f
C60344 _0310_ _0773_/a_285_297# 0
C60345 _0083_ _0261_ 0.02435f
C60346 hold28/a_285_47# _1049_/a_27_47# 0
C60347 hold28/a_49_47# _1049_/a_193_47# 0
C60348 _0965_/a_377_297# clknet_1_0__leaf_clk 0.00281f
C60349 _0154_ _1055_/a_193_47# 0.00175f
C60350 hold35/a_391_47# _1055_/a_1059_315# 0.01554f
C60351 hold87/a_391_47# _0852_/a_35_297# 0
C60352 VPWR _0989_/a_592_47# 0
C60353 VPWR _0997_/a_891_413# 0.19165f
C60354 _0810_/a_113_47# _0283_ 0
C60355 _0421_ _0655_/a_109_93# 0
C60356 _0678_/a_150_297# _0347_ 0
C60357 hold64/a_285_47# net105 0
C60358 _1059_/a_466_413# _0369_ 0
C60359 _0183_ _1019_/a_1059_315# 0.00567f
C60360 _0217_ _1019_/a_381_47# 0
C60361 net55 _0332_ 0.00553f
C60362 _0433_ clknet_1_1__leaf__0458_ 0.09992f
C60363 VPWR _0992_/a_592_47# 0
C60364 _0520_/a_27_297# net9 0
C60365 _1018_/a_1059_315# _0115_ 0
C60366 net104 _0582_/a_109_47# 0
C60367 pp[8] acc0.A\[11\] 0.00689f
C60368 _0355_ clknet_1_1__leaf__0462_ 0
C60369 net103 acc0.A\[15\] 0
C60370 _0765_/a_79_21# _0385_ 0.07573f
C60371 _0664_/a_79_21# acc0.A\[11\] 0
C60372 _1035_/a_1059_315# _0175_ 0
C60373 pp[28] _1011_/a_193_47# 0
C60374 _0749_/a_299_297# _0104_ 0
C60375 VPWR _1061_/a_561_413# 0.00323f
C60376 net55 _0685_/a_68_297# 0.1194f
C60377 net201 clknet_1_0__leaf__0461_ 0
C60378 net67 _0656_/a_59_75# 0.20759f
C60379 net58 _0439_ 0
C60380 net21 _0537_/a_68_297# 0
C60381 clknet_1_0__leaf__0463_ _1046_/a_466_413# 0
C60382 clkbuf_1_0__f__0461_/a_110_47# _0771_/a_27_413# 0.00109f
C60383 _0220_ clknet_1_1__leaf__0461_ 0
C60384 _0244_ _0454_ 0
C60385 _0310_ _0350_ 0
C60386 _1034_/a_561_413# _0173_ 0
C60387 _1034_/a_1059_315# _0208_ 0.0159f
C60388 net58 VPWR 1.47929f
C60389 hold87/a_391_47# _0081_ 0
C60390 _0241_ acc0.A\[19\] 0.99749f
C60391 _1035_/a_891_413# control0.sh 0.01889f
C60392 VPWR hold7/a_49_47# 0.31334f
C60393 _0176_ _0548_/a_51_297# 0.02016f
C60394 _0800_/a_240_47# _0799_/a_80_21# 0
C60395 _0343_ _0796_/a_79_21# 0.00851f
C60396 _0954_/a_32_297# _1044_/a_1059_315# 0.00119f
C60397 net32 net128 0.05078f
C60398 hold31/a_49_47# acc0.A\[8\] 0.32643f
C60399 net233 acc0.A\[15\] 0.00521f
C60400 _1070_/a_891_413# control0.count\[0\] 0
C60401 control0.count\[1\] _1069_/a_891_413# 0.06769f
C60402 _0975_/a_59_75# _0487_ 0.00808f
C60403 VPWR _1069_/a_1017_47# 0
C60404 _0117_ _0099_ 0
C60405 pp[25] hold53/a_49_47# 0.00226f
C60406 net53 hold53/a_391_47# 0.02984f
C60407 _0465_ _0630_/a_109_297# 0
C60408 net68 _0183_ 0
C60409 _0594_/a_113_47# net48 0
C60410 hold18/a_391_47# _0264_ 0.02031f
C60411 _1030_/a_27_47# _0336_ 0.00467f
C60412 _1030_/a_193_47# _0220_ 0
C60413 net185 _1066_/a_634_159# 0
C60414 _1018_/a_193_47# _0218_ 0
C60415 net15 pp[5] 0
C60416 _0323_ _0743_/a_51_297# 0.00406f
C60417 net31 net10 0
C60418 _0369_ _1005_/a_27_47# 0
C60419 _0762_/a_215_47# _1005_/a_1059_315# 0
C60420 _1011_/a_891_413# net57 0.00656f
C60421 _0985_/a_592_47# _0186_ 0
C60422 _0083_ _0509_/a_27_47# 0.00141f
C60423 _1000_/a_193_47# _0245_ 0.02949f
C60424 net50 acc0.A\[23\] 0.14031f
C60425 _0525_/a_299_297# _0525_/a_384_47# 0
C60426 _0216_ clknet_0__0461_ 0
C60427 clknet_0__0458_ _0824_/a_145_75# 0
C60428 acc0.A\[2\] _0630_/a_109_297# 0
C60429 _0182_ _0146_ 0.06599f
C60430 _1006_/a_634_159# _1006_/a_1017_47# 0
C60431 _1006_/a_466_413# _1006_/a_592_47# 0.00553f
C60432 net183 VPWR 0.13784f
C60433 _0993_/a_634_159# net246 0
C60434 _0240_ _0392_ 0.18682f
C60435 net182 _1055_/a_1059_315# 0.00339f
C60436 _0179_ _0858_/a_27_47# 0
C60437 net231 _0487_ 0.17735f
C60438 _0369_ _0392_ 0
C60439 net56 _0219_ 0.03477f
C60440 _1052_/a_891_413# A[5] 0
C60441 clknet_1_0__leaf__0460_ _0754_/a_245_297# 0
C60442 _0695_/a_217_297# _0219_ 0.00636f
C60443 _0984_/a_466_413# _0984_/a_381_47# 0.03733f
C60444 _0984_/a_193_47# _0984_/a_975_413# 0
C60445 _0984_/a_1059_315# _0984_/a_891_413# 0.31086f
C60446 clknet_1_0__leaf__0462_ _0379_ 0.00621f
C60447 _0714_/a_51_297# net42 0
C60448 _0569_/a_27_297# clknet_1_1__leaf__0462_ 0.00118f
C60449 _0808_/a_81_21# _0419_ 0.10384f
C60450 _0808_/a_368_297# _0417_ 0.00284f
C60451 hold100/a_49_47# net165 0
C60452 _0438_ _0988_/a_27_47# 0
C60453 net58 output62/a_27_47# 0.00647f
C60454 _0178_ _0181_ 0.22363f
C60455 acc0.A\[26\] _0687_/a_145_75# 0.00121f
C60456 net213 hold3/a_49_47# 0
C60457 net23 clkbuf_1_1__f_clk/a_110_47# 0
C60458 _0101_ VPWR 0.49685f
C60459 hold97/a_49_47# _0365_ 0
C60460 hold66/a_391_47# _0352_ 0
C60461 clknet_0__0464_ net135 0.02315f
C60462 net56 _0728_/a_59_75# 0
C60463 comp0.B\[5\] hold84/a_49_47# 0
C60464 _1039_/a_561_413# VPWR 0.00225f
C60465 _0195_ _0264_ 0.07658f
C60466 net44 hold92/a_391_47# 0.0079f
C60467 control0.state\[0\] net226 0
C60468 _0986_/a_634_159# _0986_/a_1017_47# 0
C60469 _0986_/a_466_413# _0986_/a_592_47# 0.00553f
C60470 _0589_/a_113_47# _0345_ 0
C60471 _1023_/a_634_159# net109 0
C60472 _1023_/a_193_47# net177 0.28772f
C60473 _1023_/a_891_413# _1023_/a_1017_47# 0.00617f
C60474 _0816_/a_68_297# _0218_ 0.172f
C60475 _1037_/a_193_47# _0175_ 0.00303f
C60476 acc0.A\[10\] net228 0
C60477 net216 acc0.A\[24\] 0
C60478 hold25/a_49_47# _0176_ 0.01695f
C60479 _1044_/a_891_413# _0540_/a_51_297# 0
C60480 net104 net47 0
C60481 clknet_1_0__leaf__0458_ hold18/a_285_47# 0.01482f
C60482 _0662_/a_299_297# VPWR 0.28127f
C60483 net117 pp[30] 0
C60484 net23 _0584_/a_109_297# 0.00625f
C60485 control0.state\[1\] _0946_/a_30_53# 0.12171f
C60486 clknet_1_1__leaf__0464_ _1044_/a_1017_47# 0
C60487 VPWR hold4/a_285_47# 0.27259f
C60488 output36/a_27_47# pp[0] 0.16042f
C60489 _1045_/a_1059_315# _0142_ 0
C60490 _1037_/a_634_159# control0.sh 0.00213f
C60491 net233 _0179_ 0.18736f
C60492 comp0.B\[2\] clknet_1_0__leaf__0461_ 0
C60493 _0718_/a_285_47# hold62/a_49_47# 0.00256f
C60494 _0331_ _1008_/a_27_47# 0
C60495 net243 _0380_ 0.00246f
C60496 _1036_/a_592_47# comp0.B\[4\] 0
C60497 _0466_ _1064_/a_592_47# 0
C60498 _0195_ net170 0.30549f
C60499 _0230_ acc0.A\[24\] 0
C60500 _0129_ _1031_/a_193_47# 0.04017f
C60501 net10 net128 0.01058f
C60502 _0368_ _0359_ 0.12734f
C60503 clkbuf_1_1__f__0460_/a_110_47# _0356_ 0
C60504 _0341_ _0195_ 0.04238f
C60505 _0616_/a_78_199# _0616_/a_493_297# 0
C60506 net208 hold61/a_285_47# 0.00868f
C60507 net64 hold31/a_49_47# 0.03837f
C60508 _1059_/a_193_47# net229 0.06707f
C60509 hold31/a_285_47# _0621_/a_35_297# 0.00232f
C60510 hold22/a_285_47# acc0.A\[7\] 0.08434f
C60511 net165 _0450_ 0.04501f
C60512 _1057_/a_1059_315# net192 0
C60513 _0101_ net48 0.0386f
C60514 _1038_/a_193_47# _1037_/a_1059_315# 0
C60515 _1038_/a_634_159# _1037_/a_466_413# 0.00126f
C60516 _1038_/a_27_47# _1037_/a_891_413# 0
C60517 _1038_/a_466_413# _1037_/a_634_159# 0
C60518 _1038_/a_891_413# _1037_/a_27_47# 0
C60519 _0476_ net160 0.05367f
C60520 _0257_ _0835_/a_78_199# 0.02026f
C60521 clkbuf_1_0__f__0457_/a_110_47# net187 0.02672f
C60522 _0981_/a_109_47# _0466_ 0
C60523 _0294_ _0114_ 0
C60524 _0294_ _0615_/a_109_297# 0.00158f
C60525 _0997_/a_193_47# _0095_ 0.18066f
C60526 _0997_/a_381_47# _0407_ 0
C60527 _0227_ _0374_ 0.34836f
C60528 _0855_/a_299_297# _0265_ 0
C60529 _0852_/a_35_297# _0264_ 0.10161f
C60530 _0343_ _0614_/a_29_53# 0.00101f
C60531 hold19/a_49_47# _0185_ 0
C60532 _0743_/a_51_297# net237 0.24983f
C60533 _0777_/a_285_47# _0394_ 0.06696f
C60534 _0100_ _0765_/a_79_21# 0.0566f
C60535 _1065_/a_27_47# _1065_/a_193_47# 0.96066f
C60536 net150 _0760_/a_47_47# 0.00534f
C60537 net232 _1066_/a_27_47# 0.13935f
C60538 hold30/a_285_47# _0183_ 0.08504f
C60539 hold30/a_391_47# acc0.A\[22\] 0.01082f
C60540 _0571_/a_109_47# acc0.A\[27\] 0
C60541 _0532_/a_299_297# _0532_/a_384_47# 0
C60542 hold85/a_285_47# net1 0
C60543 input11/a_75_212# input15/a_75_212# 0.0849f
C60544 VPWR _0262_ 0.43552f
C60545 _0714_/a_149_47# net162 0
C60546 net48 hold4/a_285_47# 0.00176f
C60547 _0743_/a_149_47# _0219_ 0.00376f
C60548 clknet_1_1__leaf__0463_ _1067_/a_193_47# 0
C60549 _0305_ _0347_ 0.1389f
C60550 _0637_/a_311_297# acc0.A\[15\] 0
C60551 _0349_ _0347_ 0.26675f
C60552 _0216_ _1013_/a_466_413# 0
C60553 _0324_ _0181_ 0
C60554 VPWR _0957_/a_32_297# 0.32584f
C60555 _0081_ _0264_ 0
C60556 net118 net17 0
C60557 VPWR _0582_/a_109_297# 0.17812f
C60558 hold38/a_285_47# net119 0
C60559 VPWR _1007_/a_193_47# 0.3413f
C60560 _0399_ _0989_/a_27_47# 0
C60561 VPWR _1035_/a_1017_47# 0
C60562 net180 _1040_/a_891_413# 0
C60563 _0172_ _1040_/a_466_413# 0.00487f
C60564 _0137_ _1040_/a_193_47# 0
C60565 _0550_/a_51_297# net174 0
C60566 _1001_/a_975_413# net45 0
C60567 _1058_/a_466_413# VPWR 0.25022f
C60568 _0179_ _1051_/a_27_47# 0.02646f
C60569 VPWR net23 0.81921f
C60570 _0345_ _0219_ 2.90714f
C60571 _0982_/a_592_47# _0181_ 0
C60572 _0399_ _0992_/a_27_47# 0
C60573 clknet_1_0__leaf__0465_ _0142_ 0.02318f
C60574 _0311_ _0371_ 0
C60575 _0992_/a_592_47# _0283_ 0
C60576 _0207_ net29 0.23292f
C60577 _0669_/a_111_297# _0345_ 0
C60578 _1055_/a_891_413# _0516_/a_109_297# 0
C60579 _0458_ _0275_ 0
C60580 _1064_/a_193_47# _1064_/a_592_47# 0.00135f
C60581 _1064_/a_466_413# _1064_/a_561_413# 0.00772f
C60582 _1064_/a_634_159# _1064_/a_975_413# 0
C60583 _0235_ _0373_ 0.01436f
C60584 clkbuf_0_clk/a_110_47# clknet_1_1__leaf_clk 0
C60585 _1018_/a_381_47# net149 0
C60586 _0728_/a_59_75# _0345_ 0.0111f
C60587 _0441_ _0270_ 0
C60588 _0440_ _0256_ 0
C60589 _0234_ _0750_/a_181_47# 0
C60590 _0467_ _0477_ 0.12696f
C60591 hold34/a_285_47# _0512_/a_27_297# 0
C60592 _0402_ net38 0
C60593 clknet_1_1__leaf__0465_ _0988_/a_27_47# 0
C60594 clknet_1_1__leaf_clk _1063_/a_634_159# 0
C60595 _0707_/a_544_297# _0334_ 0
C60596 net33 _1065_/a_27_47# 0
C60597 _0440_ _0987_/a_1059_315# 0.00829f
C60598 _0672_/a_215_47# _0301_ 0.0058f
C60599 _0244_ _0771_/a_382_47# 0
C60600 hold97/a_391_47# _0350_ 0
C60601 _0786_/a_217_297# VPWR 0.19792f
C60602 hold78/a_49_47# _0712_/a_297_297# 0
C60603 hold78/a_285_47# _0712_/a_79_21# 0
C60604 _0770_/a_79_21# _1001_/a_891_413# 0
C60605 _1004_/a_27_47# net93 0
C60606 clkbuf_1_0__f__0459_/a_110_47# _1060_/a_193_47# 0.00789f
C60607 _0244_ _0310_ 0
C60608 pp[16] VPWR 0.29575f
C60609 net137 _0524_/a_109_47# 0
C60610 _1051_/a_381_47# net12 0.00131f
C60611 _0316_ _0701_/a_209_297# 0
C60612 _1002_/a_634_159# _0369_ 0
C60613 _0752_/a_300_297# _0227_ 0.03479f
C60614 _0343_ _1017_/a_1059_315# 0.00439f
C60615 net40 _0218_ 0
C60616 _1056_/a_193_47# _1056_/a_975_413# 0
C60617 _0123_ net111 0
C60618 hold41/a_391_47# _0512_/a_27_297# 0
C60619 _0179_ net143 0
C60620 net117 _0339_ 0.00376f
C60621 _0183_ _0774_/a_68_297# 0.00469f
C60622 net168 VPWR 0.40261f
C60623 control0.state\[1\] _0967_/a_109_93# 0.12629f
C60624 control0.state\[0\] _0967_/a_215_297# 0.14407f
C60625 _0399_ hold60/a_49_47# 0.08718f
C60626 net34 _0485_ 0.02684f
C60627 control0.state\[1\] _0487_ 0.90231f
C60628 VPWR _0328_ 0.34527f
C60629 net35 VPWR 1.11407f
C60630 net49 _0486_ 0
C60631 _0701_/a_209_297# _0347_ 0.00101f
C60632 _0664_/a_79_21# _0281_ 0.02032f
C60633 _0285_ _0806_/a_113_297# 0.00177f
C60634 clknet_0__0465_ _0445_ 0.00554f
C60635 _1017_/a_466_413# acc0.A\[17\] 0
C60636 _0174_ _0209_ 0.07033f
C60637 net124 net24 0
C60638 net96 _0350_ 0.08021f
C60639 clknet_1_0__leaf__0462_ net53 0.23218f
C60640 _0477_ comp0.B\[0\] 0.0272f
C60641 output55/a_27_47# _0195_ 0.01313f
C60642 _0737_/a_285_47# _0364_ 0.00206f
C60643 _1008_/a_634_159# _0345_ 0
C60644 net58 _0453_ 0
C60645 _0118_ _0579_/a_27_297# 0.10962f
C60646 _0963_/a_35_297# _1070_/a_1059_315# 0
C60647 clknet_1_1__leaf__0464_ _1042_/a_891_413# 0
C60648 net125 control0.sh 0
C60649 _0836_/a_68_297# _0830_/a_79_21# 0
C60650 hold74/a_391_47# _1016_/a_193_47# 0
C60651 net157 net147 0.00362f
C60652 clkbuf_1_1__f_clk/a_110_47# _1063_/a_466_413# 0
C60653 _0204_ _0543_/a_150_297# 0
C60654 _0412_ _0997_/a_27_47# 0
C60655 _0712_/a_297_297# _0129_ 0.00877f
C60656 _0830_/a_79_21# net212 0.12785f
C60657 _0255_ _0346_ 0.03741f
C60658 hold6/a_285_47# net153 0.00997f
C60659 _0227_ _0249_ 0
C60660 _0787_/a_209_47# VPWR 0.00393f
C60661 _1015_/a_193_47# clknet_1_0__leaf__0461_ 0.00175f
C60662 net1 _0958_/a_27_47# 0.03977f
C60663 net8 net7 0
C60664 clknet_1_0__leaf__0465_ _1052_/a_891_413# 0.00315f
C60665 _0272_ clkbuf_0__0465_/a_110_47# 0.00257f
C60666 _0643_/a_253_47# clknet_0__0465_ 0.00102f
C60667 _1038_/a_193_47# _0553_/a_245_297# 0
C60668 init net33 0.0072f
C60669 _0812_/a_79_21# _0181_ 0
C60670 _0195_ _0532_/a_81_21# 0.01931f
C60671 _1037_/a_561_413# VPWR 0.00309f
C60672 _0557_/a_51_297# _0557_/a_512_297# 0.0116f
C60673 net9 _1047_/a_466_413# 0
C60674 _0255_ net65 0
C60675 _0175_ _1062_/a_193_47# 0
C60676 net7 net32 0
C60677 _0465_ _0913_/a_27_47# 0
C60678 _0402_ hold81/a_285_47# 0.00179f
C60679 _0315_ _0350_ 0
C60680 _0366_ _0380_ 0
C60681 hold23/a_49_47# _0179_ 0
C60682 net43 _0792_/a_80_21# 0
C60683 _0489_ _0976_/a_218_374# 0
C60684 pp[15] _0995_/a_592_47# 0
C60685 _0800_/a_51_297# _0668_/a_297_47# 0
C60686 _1034_/a_634_159# _0477_ 0
C60687 net91 _0103_ 0.00349f
C60688 hold43/a_49_47# hold44/a_391_47# 0
C60689 _0648_/a_27_297# clknet_1_1__leaf__0459_ 0.00141f
C60690 _0835_/a_215_47# _0465_ 0
C60691 clknet_1_1__leaf_clk _1062_/a_381_47# 0.0213f
C60692 _1018_/a_466_413# _0581_/a_27_297# 0
C60693 _1018_/a_634_159# _0581_/a_109_297# 0
C60694 VPWR _0831_/a_285_297# 0.24638f
C60695 _1060_/a_592_47# _0185_ 0
C60696 _0488_ _1069_/a_634_159# 0
C60697 _0976_/a_76_199# clknet_1_0__leaf_clk 0.00868f
C60698 _0466_ _1069_/a_193_47# 0.0019f
C60699 pp[27] _0707_/a_201_297# 0.00327f
C60700 hold91/a_285_47# hold91/a_391_47# 0.41909f
C60701 _1020_/a_27_47# _1020_/a_561_413# 0.0027f
C60702 _1020_/a_634_159# _1020_/a_891_413# 0.03684f
C60703 _1020_/a_193_47# _1020_/a_381_47# 0.09799f
C60704 _1002_/a_381_47# _0100_ 0.12468f
C60705 hold18/a_49_47# hold18/a_285_47# 0.22264f
C60706 _0405_ net42 0.00199f
C60707 _0408_ _0790_/a_285_297# 0.00293f
C60708 _0792_/a_303_47# _0406_ 0.00112f
C60709 hold12/a_285_47# hold12/a_391_47# 0.41909f
C60710 net24 _0494_/a_27_47# 0
C60711 clkbuf_1_0__f__0464_/a_110_47# _1049_/a_193_47# 0.01152f
C60712 _0820_/a_215_47# net214 0.08542f
C60713 _0107_ _0746_/a_384_47# 0
C60714 input18/a_75_212# net10 0.00316f
C60715 _0983_/a_891_413# net47 0.04803f
C60716 _1016_/a_1059_315# net43 0
C60717 _0684_/a_59_75# clknet_1_1__leaf__0460_ 0
C60718 _0209_ _0208_ 0
C60719 _1028_/a_27_47# hold50/a_391_47# 0
C60720 _1028_/a_193_47# hold50/a_285_47# 0
C60721 _1058_/a_381_47# clknet_1_1__leaf__0465_ 0.00708f
C60722 net125 net157 0.07665f
C60723 _0157_ _0369_ 0
C60724 _0747_/a_297_297# _0250_ 0
C60725 _0180_ _1048_/a_891_413# 0.0093f
C60726 _0199_ _1048_/a_634_159# 0
C60727 _0998_/a_27_47# _1017_/a_891_413# 0
C60728 _0998_/a_193_47# _1017_/a_1059_315# 0
C60729 _1013_/a_27_47# net99 0.22685f
C60730 net141 acc0.A\[6\] 0
C60731 _0782_/a_27_47# _0526_/a_27_47# 0.00151f
C60732 _0683_/a_113_47# _0366_ 0
C60733 _1041_/a_27_47# net180 0
C60734 _0457_ _0584_/a_373_47# 0
C60735 clknet_1_1__leaf__0459_ output39/a_27_47# 0
C60736 _0222_ _0369_ 0.00426f
C60737 _1003_/a_891_413# _0466_ 0
C60738 _0244_ _0768_/a_27_47# 0
C60739 _0349_ hold95/a_49_47# 0.04696f
C60740 _0337_ hold95/a_391_47# 0
C60741 _0181_ _0347_ 0.4904f
C60742 output56/a_27_47# net57 0
C60743 _0389_ clknet_1_0__leaf__0461_ 0
C60744 _0459_ clknet_1_1__leaf__0465_ 0
C60745 _0473_ control0.sh 0.02697f
C60746 hold94/a_391_47# _0754_/a_51_297# 0
C60747 _0352_ hold40/a_391_47# 0.04745f
C60748 _0176_ _0540_/a_149_47# 0
C60749 _1039_/a_381_47# _0913_/a_27_47# 0
C60750 net44 _0336_ 0.02702f
C60751 VPWR clknet_1_0__leaf__0464_ 3.08218f
C60752 _0622_/a_193_47# _0253_ 0
C60753 _0992_/a_27_47# _0295_ 0
C60754 _0536_/a_51_297# net135 0
C60755 _0144_ _1049_/a_27_47# 0
C60756 _1036_/a_1059_315# net24 0
C60757 clkload1/a_110_47# clkload1/Y 0.00568f
C60758 _0272_ _0824_/a_59_75# 0.00109f
C60759 _0172_ net154 0.02219f
C60760 _0098_ _0775_/a_510_47# 0
C60761 _1058_/a_27_47# _1057_/a_193_47# 0.00106f
C60762 _1058_/a_193_47# _1057_/a_27_47# 0.00106f
C60763 _0580_/a_373_47# _0350_ 0
C60764 comp0.B\[12\] _1044_/a_975_413# 0
C60765 _0534_/a_299_297# clknet_1_1__leaf__0457_ 0.05444f
C60766 _0219_ net52 0.07031f
C60767 _0642_/a_27_413# _0433_ 0
C60768 net226 _0478_ 0.01173f
C60769 net7 net10 0
C60770 net35 hold17/a_285_47# 0.00114f
C60771 _1000_/a_466_413# _0347_ 0.02091f
C60772 _1000_/a_27_47# _0352_ 0.03552f
C60773 _0257_ _0399_ 0
C60774 _0414_ _0994_/a_975_413# 0
C60775 VPWR _1063_/a_466_413# 0.2471f
C60776 _0664_/a_297_47# _0654_/a_207_413# 0
C60777 _0243_ net47 0
C60778 _0402_ _0282_ 0
C60779 _1052_/a_975_413# net73 0
C60780 hold66/a_391_47# _0237_ 0.01965f
C60781 hold66/a_49_47# _0382_ 0
C60782 _0216_ net97 0.00433f
C60783 _0572_/a_27_297# _0124_ 0.11012f
C60784 _0572_/a_373_47# net155 0.00276f
C60785 acc0.A\[14\] acc0.A\[13\] 0.584f
C60786 _0179_ _0085_ 0
C60787 hold47/a_285_47# net135 0
C60788 _0647_/a_285_47# _0218_ 0
C60789 acc0.A\[3\] _0186_ 0.3965f
C60790 acc0.A\[1\] acc0.A\[0\] 0.08158f
C60791 _0266_ _0263_ 0
C60792 acc0.A\[26\] _0739_/a_510_47# 0.0017f
C60793 _0856_/a_79_21# _0195_ 0
C60794 _0443_ _0841_/a_510_47# 0.00136f
C60795 net190 hold9/a_49_47# 0.04309f
C60796 net197 hold9/a_391_47# 0.03999f
C60797 _0172_ _0465_ 0
C60798 net165 net219 0
C60799 _0804_/a_79_21# clknet_1_1__leaf__0459_ 0
C60800 _0274_ _0268_ 0
C60801 _0984_/a_27_47# net229 0
C60802 hold55/a_285_47# net118 0.01823f
C60803 _0127_ clknet_1_1__leaf__0462_ 0
C60804 clkbuf_1_0__f_clk/a_110_47# control0.count\[0\] 0.03432f
C60805 VPWR _1060_/a_466_413# 0.2573f
C60806 _1019_/a_193_47# _0242_ 0
C60807 pp[28] _0707_/a_75_199# 0.01777f
C60808 net220 _0369_ 0.09899f
C60809 _0090_ acc0.A\[10\] 0.00421f
C60810 _0856_/a_79_21# _0856_/a_510_47# 0.00844f
C60811 _0856_/a_297_297# _0856_/a_215_47# 0
C60812 hold75/a_391_47# _0465_ 0.00257f
C60813 _0137_ _0207_ 0.0298f
C60814 VPWR _0988_/a_975_413# 0.00483f
C60815 VPWR _0553_/a_240_47# 0.01585f
C60816 _0499_/a_59_75# _0171_ 0.1733f
C60817 _0108_ VPWR 0.53116f
C60818 pp[8] A[12] 0.16694f
C60819 _1054_/a_1059_315# _0186_ 0
C60820 clkbuf_0__0463_/a_110_47# acc0.A\[15\] 0.01178f
C60821 _0791_/a_113_297# _0219_ 0.00147f
C60822 _0174_ _1043_/a_466_413# 0.00883f
C60823 _0786_/a_217_297# _0283_ 0.0521f
C60824 hold75/a_285_47# net58 0.10017f
C60825 net190 _1029_/a_27_47# 0
C60826 net157 _1047_/a_1059_315# 0.00123f
C60827 _0216_ _0616_/a_215_47# 0.01837f
C60828 _0311_ _0767_/a_59_75# 0
C60829 _0473_ net157 0.00709f
C60830 _1023_/a_592_47# acc0.A\[23\] 0
C60831 _0088_ net47 0.02827f
C60832 net82 _0996_/a_27_47# 0.2249f
C60833 control0.add _0350_ 0.3046f
C60834 _0619_/a_68_297# _0989_/a_27_47# 0
C60835 _1016_/a_891_413# _0181_ 0.00431f
C60836 net219 acc0.A\[19\] 0
C60837 _0369_ acc0.A\[9\] 0.02947f
C60838 net3 acc0.A\[10\] 0
C60839 _0236_ _0603_/a_150_297# 0
C60840 _0231_ _0227_ 0
C60841 _0094_ net5 0.13776f
C60842 _0670_/a_215_47# _0670_/a_510_47# 0.00529f
C60843 _0433_ _0218_ 0.0063f
C60844 _1031_/a_27_47# clknet_1_1__leaf__0462_ 0.00146f
C60845 pp[27] _1010_/a_27_47# 0
C60846 _0732_/a_303_47# _0359_ 0
C60847 output59/a_27_47# _0110_ 0
C60848 _0325_ _0368_ 0
C60849 _0322_ _0686_/a_219_297# 0.01507f
C60850 net137 _0142_ 0
C60851 comp0.B\[11\] net32 0.01731f
C60852 _0183_ hold71/a_49_47# 0
C60853 net155 acc0.A\[27\] 0.00503f
C60854 _0457_ _1015_/a_891_413# 0.00497f
C60855 comp0.B\[1\] _0181_ 0
C60856 _0322_ _1008_/a_1059_315# 0
C60857 _0329_ _1008_/a_466_413# 0
C60858 _0327_ _0686_/a_219_297# 0.01143f
C60859 _0337_ net209 0
C60860 _0380_ _0378_ 0
C60861 net56 net94 0
C60862 comp0.B\[5\] control0.reset 0.00143f
C60863 clkbuf_1_0__f__0463_/a_110_47# net173 0.00131f
C60864 _0234_ _0606_/a_109_53# 0.02458f
C60865 _1001_/a_975_413# VPWR 0.00464f
C60866 net45 _1017_/a_381_47# 0.00278f
C60867 VPWR _1062_/a_561_413# 0.00292f
C60868 _1018_/a_27_47# _0347_ 0.00176f
C60869 _0370_ acc0.A\[24\] 0
C60870 _0849_/a_297_297# acc0.A\[15\] 0
C60871 clkbuf_0__0465_/a_110_47# _0181_ 0.00445f
C60872 _0359_ clknet_0__0460_ 0.05153f
C60873 _1039_/a_381_47# _0172_ 0
C60874 _1039_/a_1059_315# _0137_ 0.04695f
C60875 _1021_/a_891_413# VPWR 0.19996f
C60876 _1038_/a_634_159# _0135_ 0
C60877 hold58/a_285_47# _0557_/a_51_297# 0
C60878 _0343_ _0373_ 0
C60879 acc0.A\[1\] _0580_/a_109_297# 0
C60880 _0762_/a_297_297# _0369_ 0.00174f
C60881 _0279_ _0647_/a_377_297# 0.00468f
C60882 _0343_ hold88/a_49_47# 0.02371f
C60883 _0810_/a_113_47# _0345_ 0
C60884 _0278_ _0647_/a_47_47# 0
C60885 _0365_ _0738_/a_150_297# 0
C60886 clkbuf_0__0458_/a_110_47# _0841_/a_79_21# 0.00298f
C60887 _0531_/a_27_297# _0178_ 0.00104f
C60888 _0266_ clknet_1_0__leaf__0461_ 0.00169f
C60889 comp0.B\[6\] _0207_ 0.0238f
C60890 acc0.A\[17\] _0393_ 0
C60891 _0776_/a_27_47# _0394_ 0.0532f
C60892 hold10/a_391_47# net36 0.05797f
C60893 _0195_ _0454_ 0
C60894 net175 net149 0
C60895 hold14/a_285_47# _0175_ 0.00795f
C60896 _1065_/a_466_413# _1065_/a_592_47# 0.00553f
C60897 _1065_/a_634_159# _1065_/a_1017_47# 0
C60898 _0677_/a_377_297# _0347_ 0
C60899 input27/a_75_212# _0175_ 0
C60900 VPWR _0213_ 0.44372f
C60901 _0592_/a_68_297# _1022_/a_1059_315# 0
C60902 clknet_0_clk _1062_/a_27_47# 0.00934f
C60903 hold69/a_49_47# _0460_ 0
C60904 _0967_/a_215_297# _1066_/a_193_47# 0.00206f
C60905 hold28/a_49_47# VPWR 0.31249f
C60906 _0485_ _1066_/a_466_413# 0
C60907 hold66/a_285_47# _1005_/a_193_47# 0
C60908 _0817_/a_266_47# _0991_/a_1059_315# 0
C60909 _0998_/a_975_413# _0218_ 0
C60910 _0746_/a_81_21# net52 0.0226f
C60911 _0520_/a_109_297# net13 0.00785f
C60912 _1036_/a_27_47# net23 0
C60913 _1036_/a_193_47# B[15] 0
C60914 _1068_/a_27_47# _0162_ 0
C60915 _1068_/a_634_159# _0487_ 0
C60916 _0992_/a_193_47# _0811_/a_81_21# 0
C60917 _0394_ _0219_ 0.02583f
C60918 _0571_/a_27_297# _1027_/a_193_47# 0
C60919 net189 _0992_/a_1059_315# 0
C60920 _1033_/a_891_413# net201 0.00359f
C60921 _0429_ _0399_ 0
C60922 comp0.B\[11\] _1042_/a_1059_315# 0.06616f
C60923 comp0.B\[12\] _1042_/a_466_413# 0
C60924 _0770_/a_297_47# _0241_ 0.00299f
C60925 _1014_/a_634_159# _1014_/a_381_47# 0
C60926 _0452_ _0265_ 0.18361f
C60927 net32 _0202_ 0
C60928 _1071_/a_27_47# _1071_/a_634_159# 0.14145f
C60929 acc0.A\[15\] hold71/a_49_47# 0.03636f
C60930 _0996_/a_193_47# _0796_/a_79_21# 0
C60931 control0.count\[2\] control0.count\[0\] 0.50084f
C60932 VPWR _1047_/a_592_47# 0
C60933 pp[30] _0704_/a_68_297# 0.00172f
C60934 _0183_ hold72/a_391_47# 0
C60935 _1015_/a_634_159# _0173_ 0
C60936 _0130_ _0565_/a_512_297# 0.00102f
C60937 VPWR output51/a_27_47# 0.30029f
C60938 pp[27] pp[30] 0.17017f
C60939 _0985_/a_466_413# _0458_ 0.01322f
C60940 _0352_ _0374_ 0.02762f
C60941 _0476_ _1034_/a_193_47# 0
C60942 _0172_ net174 0.06347f
C60943 _1050_/a_193_47# net9 0.03212f
C60944 _0458_ _1049_/a_27_47# 0
C60945 _1021_/a_891_413# net48 0.00103f
C60946 _0179_ net131 0
C60947 hold87/a_391_47# _0183_ 0
C60948 VPWR _0536_/a_245_297# 0.00558f
C60949 _0541_/a_68_297# hold51/a_391_47# 0.00359f
C60950 comp0.B\[11\] net10 0.30447f
C60951 VPWR _0796_/a_215_47# 0.00779f
C60952 net54 _0690_/a_68_297# 0.00117f
C60953 _1039_/a_1059_315# comp0.B\[6\] 0
C60954 _0717_/a_209_297# _0334_ 0.02685f
C60955 hold13/a_49_47# _0175_ 0
C60956 _0212_ VPWR 0.61331f
C60957 _1055_/a_975_413# net16 0
C60958 net65 _0830_/a_215_47# 0.06738f
C60959 _0305_ _1059_/a_27_47# 0.02507f
C60960 _0113_ net23 0.18698f
C60961 A[10] acc0.A\[11\] 0.00317f
C60962 clkbuf_1_0__f__0459_/a_110_47# _1017_/a_1059_315# 0
C60963 hold98/a_49_47# output41/a_27_47# 0.00616f
C60964 net45 _0581_/a_27_297# 0.05343f
C60965 hold63/a_49_47# net111 0.00121f
C60966 _0669_/a_29_53# _0301_ 0.10157f
C60967 net188 A[11] 0
C60968 _0664_/a_297_47# _0286_ 0.02307f
C60969 _0441_ _0085_ 0
C60970 VPWR _0547_/a_68_297# 0.16687f
C60971 _0454_ _0852_/a_35_297# 0.17016f
C60972 net2 _0510_/a_27_297# 0.01498f
C60973 _1026_/a_1059_315# acc0.A\[25\] 0
C60974 hold18/a_391_47# _0846_/a_51_297# 0
C60975 hold78/a_49_47# _0344_ 0
C60976 _1012_/a_193_47# _0347_ 0.03915f
C60977 hold67/a_285_47# net66 0.06952f
C60978 _0275_ _0291_ 0.04042f
C60979 hold67/a_49_47# acc0.A\[8\] 0
C60980 _0317_ _0352_ 0
C60981 hold13/a_285_47# control0.sh 0
C60982 net88 _0369_ 0
C60983 hold21/a_285_47# _0179_ 0.00219f
C60984 _0343_ _1016_/a_27_47# 0.01208f
C60985 hold47/a_391_47# VPWR 0.18376f
C60986 acc0.A\[28\] _0319_ 0
C60987 clknet_1_0__leaf__0462_ _0575_/a_27_297# 0.00958f
C60988 hold75/a_49_47# _0261_ 0.00143f
C60989 _0831_/a_35_297# acc0.A\[6\] 0.03624f
C60990 _1013_/a_1017_47# _0339_ 0
C60991 _0216_ _1010_/a_27_47# 0
C60992 _0981_/a_27_297# _0490_ 0.12605f
C60993 net48 output51/a_27_47# 0
C60994 output48/a_27_47# net51 0.00128f
C60995 _0195_ acc0.A\[30\] 0.31195f
C60996 clknet_1_0__leaf__0459_ _1060_/a_466_413# 0
C60997 _1052_/a_27_47# _0180_ 0.02024f
C60998 _1033_/a_634_159# clknet_1_1__leaf_clk 0
C60999 net94 _0345_ 0.02951f
C61000 _0590_/a_113_47# net151 0
C61001 _0222_ _1022_/a_975_413# 0.00148f
C61002 _0402_ _0654_/a_297_47# 0
C61003 _0855_/a_384_47# _0112_ 0
C61004 _0454_ _0081_ 0.00318f
C61005 _0963_/a_285_47# VPWR 0
C61006 _0500_/a_27_47# acc0.A\[1\] 0
C61007 _1037_/a_466_413# _1036_/a_1059_315# 0
C61008 _1037_/a_634_159# _1036_/a_891_413# 0
C61009 _0566_/a_27_47# _0208_ 0.03722f
C61010 _0179_ hold71/a_49_47# 0
C61011 _0750_/a_27_47# VPWR 0.26265f
C61012 _0571_/a_27_297# _1026_/a_1059_315# 0
C61013 _0553_/a_245_297# net29 0.00187f
C61014 _0463_ clknet_1_1__leaf__0457_ 0.00322f
C61015 _0817_/a_266_47# _0425_ 0.04058f
C61016 hold23/a_285_47# _0530_/a_299_297# 0
C61017 hold23/a_391_47# _0530_/a_81_21# 0
C61018 _0352_ acc0.A\[19\] 0.01761f
C61019 _0680_/a_80_21# _0731_/a_81_21# 0
C61020 clkbuf_1_1__f_clk/a_110_47# _0161_ 0.07674f
C61021 _0999_/a_561_413# _0352_ 0.00107f
C61022 _1013_/a_1059_315# pp[31] 0.00256f
C61023 _0344_ _0129_ 0.25235f
C61024 _0457_ net87 0
C61025 net22 _0546_/a_245_297# 0.00251f
C61026 _0498_/a_512_297# net247 0
C61027 _0220_ _0567_/a_27_297# 0
C61028 _0752_/a_300_297# _0352_ 0.00134f
C61029 _0437_ _0087_ 0.00262f
C61030 _0445_ _0986_/a_27_47# 0.10709f
C61031 _0444_ _0986_/a_193_47# 0
C61032 hold87/a_391_47# acc0.A\[15\] 0
C61033 net10 _0202_ 0
C61034 hold29/a_285_47# net51 0
C61035 net1 _0477_ 0.14397f
C61036 _0713_/a_27_47# clknet_1_0__leaf__0461_ 0
C61037 comp0.B\[2\] _1033_/a_891_413# 0.00206f
C61038 _1038_/a_891_413# _0174_ 0
C61039 _1038_/a_27_47# _0136_ 0.00865f
C61040 _0557_/a_51_297# _0134_ 0.12144f
C61041 _0183_ _1005_/a_193_47# 0
C61042 _0126_ _1028_/a_634_159# 0
C61043 _0570_/a_27_297# net114 0
C61044 net190 _1028_/a_891_413# 0.0664f
C61045 net2 _0181_ 0.46466f
C61046 _0949_/a_59_75# net231 0.00148f
C61047 hold46/a_285_47# VPWR 0.29112f
C61048 _0216_ _1014_/a_381_47# 0
C61049 net55 clknet_0__0460_ 0.25999f
C61050 hold42/a_391_47# output67/a_27_47# 0.00561f
C61051 net157 _0497_/a_68_297# 0
C61052 pp[9] _1057_/a_27_47# 0
C61053 _0992_/a_1059_315# _0417_ 0
C61054 hold67/a_285_47# _0350_ 0.06425f
C61055 acc0.A\[31\] _1013_/a_27_47# 0
C61056 _0576_/a_27_297# acc0.A\[23\] 0.10794f
C61057 net151 _1005_/a_891_413# 0
C61058 _1003_/a_1059_315# clknet_1_0__leaf__0460_ 0.00249f
C61059 _0686_/a_27_53# _0686_/a_301_297# 0
C61060 _1021_/a_27_47# _0462_ 0
C61061 _1059_/a_1059_315# acc0.A\[15\] 0.0083f
C61062 _0717_/a_80_21# pp[27] 0.00995f
C61063 VPWR _0775_/a_79_21# 0.49712f
C61064 _0280_ clknet_1_1__leaf__0459_ 0.35776f
C61065 _0279_ _0802_/a_59_75# 0
C61066 _0643_/a_253_47# _0986_/a_27_47# 0
C61067 _0643_/a_337_297# _0986_/a_193_47# 0
C61068 _0663_/a_207_413# _0179_ 0.01694f
C61069 clknet_1_1__leaf__0461_ _0347_ 0.21223f
C61070 clknet_1_0__leaf__0461_ _0612_/a_59_75# 0.00771f
C61071 _0579_/a_27_297# _1001_/a_27_47# 0.01623f
C61072 _1018_/a_466_413# _0116_ 0.03479f
C61073 _1018_/a_381_47# net206 0
C61074 _0339_ _0704_/a_68_297# 0.0039f
C61075 net106 hold40/a_391_47# 0
C61076 _1008_/a_634_159# _1008_/a_592_47# 0
C61077 _1055_/a_27_47# _1055_/a_1059_315# 0.04875f
C61078 _1055_/a_193_47# _1055_/a_466_413# 0.07911f
C61079 input21/a_75_212# net19 0
C61080 B[13] _0203_ 0
C61081 _0488_ clknet_1_0__leaf_clk 0.43404f
C61082 _0505_/a_27_297# _0505_/a_373_47# 0.01338f
C61083 _0172_ clknet_0__0464_ 0.44541f
C61084 _0349_ _1011_/a_27_47# 0
C61085 pp[27] _0339_ 0.04133f
C61086 pp[16] _0995_/a_634_159# 0
C61087 net53 _1025_/a_891_413# 0.01957f
C61088 _1020_/a_1059_315# _0118_ 0.05991f
C61089 _0249_ _0352_ 0
C61090 _0559_/a_51_297# _0173_ 0.15448f
C61091 _1003_/a_27_47# _1003_/a_634_159# 0.14145f
C61092 _0399_ clknet_1_1__leaf__0458_ 0.08833f
C61093 net166 _0583_/a_27_297# 0.00368f
C61094 net23 comp0.B\[3\] 0
C61095 _1055_/a_193_47# net181 0
C61096 _0230_ _0375_ 0.01992f
C61097 _0750_/a_27_47# net48 0
C61098 VPWR _0614_/a_183_297# 0
C61099 _0430_ _0274_ 0.04249f
C61100 pp[30] _0216_ 0.18783f
C61101 _0389_ _0218_ 0.00305f
C61102 _0243_ _0294_ 0
C61103 clknet_0__0458_ _0986_/a_561_413# 0
C61104 _0343_ pp[2] 0
C61105 net114 hold50/a_49_47# 0.04531f
C61106 clknet_0__0457_ _1014_/a_561_413# 0
C61107 clknet_0__0463_ _0533_/a_373_47# 0
C61108 control0.sh _0132_ 0
C61109 _0176_ _0542_/a_245_297# 0
C61110 net194 net9 0
C61111 _0188_ net3 0.03783f
C61112 _1054_/a_891_413# _0518_/a_109_297# 0
C61113 net84 _1017_/a_466_413# 0
C61114 net46 net223 0.58462f
C61115 _0275_ _0290_ 0.03696f
C61116 _1032_/a_891_413# comp0.B\[0\] 0.00346f
C61117 _1041_/a_592_47# _0172_ 0
C61118 _0997_/a_193_47# _0219_ 0.01609f
C61119 _0833_/a_79_21# _0439_ 0.07909f
C61120 clknet_1_0__leaf__0458_ _0445_ 0
C61121 _0452_ _0267_ 0
C61122 clkbuf_1_1__f__0461_/a_110_47# net219 0
C61123 _0217_ acc0.A\[25\] 0.10256f
C61124 _1004_/a_1059_315# _0758_/a_79_21# 0
C61125 _0714_/a_51_297# net60 0
C61126 _0846_/a_240_47# _0449_ 0.0425f
C61127 _0992_/a_592_47# _0345_ 0
C61128 net8 clkbuf_1_1__f__0457_/a_110_47# 0
C61129 VPWR _0833_/a_79_21# 0.42414f
C61130 net190 _0739_/a_79_21# 0
C61131 _0570_/a_27_297# _0365_ 0
C61132 net197 _0739_/a_215_47# 0
C61133 _0216_ _0771_/a_215_297# 0.00365f
C61134 net188 net66 0
C61135 hold94/a_391_47# _0219_ 0.0148f
C61136 net203 _1034_/a_27_47# 0.00353f
C61137 net197 _0352_ 0
C61138 _0227_ _0225_ 0.19584f
C61139 _0991_/a_975_413# acc0.A\[15\] 0
C61140 _0307_ hold72/a_49_47# 0.08434f
C61141 _0837_/a_266_47# acc0.A\[5\] 0
C61142 _0984_/a_381_47# _0184_ 0
C61143 clknet_0__0459_ _0410_ 0
C61144 _0183_ _0264_ 0.03644f
C61145 _1054_/a_27_47# _1053_/a_193_47# 0
C61146 _1054_/a_193_47# _1053_/a_27_47# 0
C61147 _0472_ net29 0
C61148 _0982_/a_634_159# _0456_ 0
C61149 _0982_/a_891_413# net234 0
C61150 _0559_/a_245_297# _0212_ 0
C61151 _0222_ _0756_/a_47_47# 0
C61152 _0123_ net199 0
C61153 net26 _0207_ 0
C61154 net187 _0217_ 0.47085f
C61155 _0399_ _0263_ 0.00525f
C61156 _0298_ _0668_/a_297_47# 0.04825f
C61157 _0299_ _0668_/a_382_297# 0
C61158 _0557_/a_51_297# _0554_/a_68_297# 0
C61159 net58 _0345_ 0.07117f
C61160 net62 acc0.A\[3\] 0
C61161 hold22/a_285_47# _0186_ 0
C61162 clknet_1_0__leaf__0459_ _0796_/a_215_47# 0
C61163 _0674_/a_113_47# clknet_0__0461_ 0
C61164 _0179_ _1059_/a_1059_315# 0
C61165 _0098_ _0347_ 0.28909f
C61166 VPWR _0161_ 1.31654f
C61167 _1059_/a_27_47# _0181_ 0
C61168 _0748_/a_81_21# _0462_ 0.00545f
C61169 _0367_ _0737_/a_117_297# 0
C61170 hold2/a_285_47# _0465_ 0.01483f
C61171 _1016_/a_891_413# clknet_1_1__leaf__0461_ 0.04193f
C61172 clknet_1_0__leaf_clk _1064_/a_27_47# 0.23461f
C61173 VPWR _1017_/a_381_47# 0.07064f
C61174 _1015_/a_27_47# _0178_ 0
C61175 _0259_ _0255_ 0.00108f
C61176 _0365_ hold50/a_49_47# 0.03078f
C61177 _1037_/a_891_413# comp0.B\[5\] 0.00299f
C61178 _1037_/a_1059_315# comp0.B\[6\] 0
C61179 _0415_ _0802_/a_145_75# 0
C61180 VPWR net127 0.33056f
C61181 _0563_/a_245_297# _0563_/a_240_47# 0
C61182 _0548_/a_245_297# net173 0
C61183 net207 acc0.A\[19\] 0
C61184 VPWR _0158_ 0.52114f
C61185 _0506_/a_299_297# _0506_/a_384_47# 0
C61186 VPWR _0543_/a_150_297# 0.0014f
C61187 pp[28] _0338_ 0.00523f
C61188 hold11/a_49_47# clknet_1_1__leaf__0464_ 0
C61189 _0398_ _0459_ 0.00186f
C61190 acc0.A\[20\] _0228_ 0.01067f
C61191 VPWR _1033_/a_466_413# 0.24281f
C61192 clknet_1_1__leaf__0460_ net191 0
C61193 _1038_/a_466_413# comp0.B\[8\] 0
C61194 _1044_/a_193_47# _0141_ 0.00339f
C61195 _1044_/a_1059_315# net19 0
C61196 _1044_/a_891_413# net195 0
C61197 clknet_1_0__leaf__0465_ _1049_/a_466_413# 0.00114f
C61198 net106 comp0.B\[0\] 0
C61199 _0343_ hold62/a_49_47# 0.02762f
C61200 _0732_/a_80_21# _0326_ 0
C61201 _0429_ _0619_/a_68_297# 0.06064f
C61202 _0252_ _0826_/a_27_53# 0
C61203 _0174_ net196 0.13351f
C61204 hold86/a_49_47# VPWR 0.24888f
C61205 _0264_ acc0.A\[15\] 0.01155f
C61206 VPWR _1050_/a_561_413# 0.00302f
C61207 net248 _0825_/a_68_297# 0
C61208 net230 _1054_/a_27_47# 0
C61209 acc0.A\[14\] _0998_/a_1017_47# 0
C61210 _0274_ _0443_ 0.03105f
C61211 _0272_ _0432_ 0.02461f
C61212 _0579_/a_109_297# clknet_1_0__leaf__0461_ 0
C61213 _1010_/a_193_47# _1010_/a_381_47# 0.09503f
C61214 _1010_/a_634_159# _1010_/a_891_413# 0.03684f
C61215 _1010_/a_27_47# _1010_/a_561_413# 0.0027f
C61216 clknet_1_0__leaf__0462_ _1004_/a_1059_315# 0.01751f
C61217 _0327_ clknet_1_1__leaf__0462_ 0.01888f
C61218 net165 _0849_/a_79_21# 0
C61219 _0991_/a_1059_315# _0181_ 0
C61220 _1040_/a_193_47# _1040_/a_466_413# 0.07482f
C61221 _1040_/a_27_47# _1040_/a_1059_315# 0.04672f
C61222 _0670_/a_79_21# _0409_ 0
C61223 _0290_ _0657_/a_109_297# 0.00283f
C61224 _0462_ clknet_0__0462_ 0.00592f
C61225 _0411_ _0219_ 0
C61226 _0305_ _0607_/a_109_297# 0.00694f
C61227 _0645_/a_47_47# clkbuf_0__0459_/a_110_47# 0
C61228 _0697_/a_80_21# _0328_ 0.11287f
C61229 _0146_ _1048_/a_1059_315# 0.02805f
C61230 _0216_ _0339_ 0.04907f
C61231 net71 _0261_ 0.00164f
C61232 _0200_ net157 0
C61233 _0399_ clknet_1_0__leaf__0461_ 0.15897f
C61234 _0266_ _0218_ 0
C61235 _0195_ _1027_/a_27_47# 0
C61236 _0662_/a_299_297# _0345_ 0.00177f
C61237 _1002_/a_466_413# _0183_ 0
C61238 _1002_/a_891_413# _0217_ 0
C61239 control0.state\[1\] _0949_/a_59_75# 0.02154f
C61240 control0.state\[0\] _0949_/a_145_75# 0
C61241 hold88/a_49_47# _0990_/a_381_47# 0
C61242 net63 _0438_ 0.00148f
C61243 _0326_ _0250_ 1.10291f
C61244 VPWR _0391_ 0.49403f
C61245 _0372_ _1006_/a_27_47# 0
C61246 _0248_ _1006_/a_193_47# 0
C61247 _0234_ _0238_ 0.0276f
C61248 _0148_ _0142_ 0.00183f
C61249 _1020_/a_975_413# _0461_ 0
C61250 clkbuf_1_1__f__0463_/a_110_47# _0562_/a_68_297# 0
C61251 _0623_/a_109_297# VPWR 0.00748f
C61252 _0846_/a_51_297# _0846_/a_149_47# 0.02487f
C61253 net45 _1016_/a_634_159# 0.00109f
C61254 _1067_/a_27_47# _1067_/a_1059_315# 0.04875f
C61255 _1067_/a_193_47# _1067_/a_466_413# 0.07495f
C61256 net9 _0987_/a_193_47# 0.03639f
C61257 _0346_ hold1/a_49_47# 0
C61258 clknet_1_0__leaf__0459_ _0775_/a_79_21# 0.00205f
C61259 net124 _0135_ 0
C61260 _1019_/a_27_47# _1015_/a_27_47# 0.00179f
C61261 hold31/a_49_47# _0369_ 0
C61262 _0231_ _0352_ 0.10525f
C61263 _0346_ _0992_/a_27_47# 0
C61264 net84 _0094_ 0
C61265 _1000_/a_27_47# _0392_ 0
C61266 _1072_/a_193_47# _1071_/a_466_413# 0
C61267 _1072_/a_27_47# _1071_/a_1059_315# 0
C61268 _0845_/a_109_297# acc0.A\[15\] 0
C61269 VPWR _0581_/a_27_297# 0.193f
C61270 _1009_/a_1059_315# _1009_/a_891_413# 0.31086f
C61271 _1009_/a_193_47# _1009_/a_975_413# 0
C61272 _1009_/a_466_413# _1009_/a_381_47# 0.03733f
C61273 _0620_/a_113_47# net65 0
C61274 net65 _0989_/a_27_47# 0.03709f
C61275 _0833_/a_510_47# clknet_1_1__leaf__0465_ 0
C61276 net65 hold1/a_49_47# 0
C61277 _0989_/a_27_47# _0989_/a_466_413# 0.27314f
C61278 _0989_/a_193_47# _0989_/a_634_159# 0.11072f
C61279 hold1/a_285_47# hold1/a_391_47# 0.41909f
C61280 acc0.A\[14\] VPWR 1.56788f
C61281 _0237_ _0374_ 0.12108f
C61282 VPWR clkbuf_1_0__f__0464_/a_110_47# 1.35455f
C61283 net1 _0352_ 0.36569f
C61284 _0238_ clknet_0__0460_ 0
C61285 _0956_/a_32_297# net201 0.05455f
C61286 comp0.B\[15\] _0565_/a_149_47# 0.00224f
C61287 hold65/a_285_47# acc0.A\[8\] 0
C61288 _1065_/a_381_47# control0.reset 0
C61289 hold5/a_391_47# _0140_ 0.00381f
C61290 hold18/a_285_47# _0448_ 0
C61291 _0982_/a_381_47# VPWR 0.07591f
C61292 _0476_ _1066_/a_891_413# 0.00188f
C61293 _0967_/a_109_93# clknet_1_1__leaf_clk 0
C61294 _0487_ clknet_1_1__leaf_clk 0.07158f
C61295 hold66/a_49_47# net91 0
C61296 _0992_/a_27_47# _0992_/a_466_413# 0.27314f
C61297 _0992_/a_193_47# _0992_/a_634_159# 0.12729f
C61298 _0817_/a_585_47# _0089_ 0
C61299 _1036_/a_975_413# net121 0
C61300 comp0.B\[4\] _1035_/a_1059_315# 0
C61301 _0307_ clknet_0__0461_ 0.31566f
C61302 _0186_ net13 0.81548f
C61303 _0607_/a_27_297# net43 0.16781f
C61304 clkbuf_1_1__f__0461_/a_110_47# _0352_ 0
C61305 VPWR _1053_/a_634_159# 0.18289f
C61306 _0125_ _1027_/a_193_47# 0.03765f
C61307 acc0.A\[27\] _1027_/a_1059_315# 0.10343f
C61308 _0718_/a_47_47# pp[27] 0.013f
C61309 _0280_ _0655_/a_215_53# 0.27697f
C61310 _1032_/a_1059_315# net118 0
C61311 hold79/a_391_47# control0.count\[1\] 0.00211f
C61312 _0557_/a_240_47# _0211_ 0.04252f
C61313 net226 VPWR 0.19497f
C61314 _1014_/a_634_159# acc0.A\[0\] 0.00216f
C61315 _1014_/a_381_47# net100 0.01524f
C61316 _0361_ _0370_ 0
C61317 _1071_/a_891_413# _1071_/a_975_413# 0.00851f
C61318 _1071_/a_381_47# _1071_/a_561_413# 0.00123f
C61319 net71 _0509_/a_27_47# 0.04363f
C61320 _0996_/a_1059_315# _0410_ 0
C61321 _0996_/a_891_413# net238 0.04385f
C61322 _0311_ _0388_ 0
C61323 _1045_/a_193_47# _1043_/a_193_47# 0.00123f
C61324 _0835_/a_78_199# _0218_ 0.012f
C61325 clkbuf_1_0__f__0458_/a_110_47# _0846_/a_51_297# 0.01717f
C61326 _1000_/a_193_47# clknet_0__0461_ 0.00464f
C61327 _1000_/a_1059_315# clkbuf_1_0__f__0461_/a_110_47# 0.01616f
C61328 _0768_/a_109_297# _0240_ 0
C61329 _0212_ _1036_/a_27_47# 0
C61330 hold96/a_285_47# net243 0.0102f
C61331 clkload4/a_110_47# _0219_ 0
C61332 _0346_ hold60/a_49_47# 0.00249f
C61333 _0327_ net242 0
C61334 _0251_ _0836_/a_68_297# 0
C61335 _0083_ _0458_ 0.11641f
C61336 net45 _0714_/a_149_47# 0
C61337 acc0.A\[16\] net42 0
C61338 _0343_ _0400_ 0.04514f
C61339 _0123_ VPWR 0.65608f
C61340 _0251_ net212 0.00146f
C61341 clknet_1_1__leaf__0459_ net143 0.00181f
C61342 _0425_ _0181_ 0.00385f
C61343 _0216_ _1026_/a_193_47# 0.02334f
C61344 net157 _1046_/a_466_413# 0
C61345 _0553_/a_245_297# comp0.B\[6\] 0.00242f
C61346 _0483_ _0481_ 0
C61347 _0363_ _0734_/a_47_47# 0.00106f
C61348 _0350_ hold50/a_391_47# 0
C61349 _0176_ input19/a_75_212# 0.00901f
C61350 _0216_ _1024_/a_891_413# 0
C61351 _0252_ _0087_ 0.20499f
C61352 _0817_/a_81_21# acc0.A\[9\] 0.01261f
C61353 _0087_ _0989_/a_381_47# 0.11472f
C61354 input6/a_75_212# pp[14] 0.00154f
C61355 _0285_ _0399_ 0
C61356 hold2/a_49_47# _0262_ 0
C61357 _0179_ net170 0
C61358 net16 _0988_/a_193_47# 0
C61359 net45 _0116_ 0.09452f
C61360 acc0.A\[10\] hold70/a_49_47# 0
C61361 _0650_/a_150_297# net37 0
C61362 _0479_ _0487_ 0
C61363 _0517_/a_81_21# _0290_ 0
C61364 clkbuf_1_0__f__0459_/a_110_47# _1016_/a_27_47# 0
C61365 net2 _0187_ 0
C61366 _1020_/a_466_413# acc0.A\[20\] 0
C61367 B[2] _0175_ 0.00394f
C61368 _0390_ _0391_ 0.06075f
C61369 _0389_ _0099_ 0
C61370 _1042_/a_634_159# _0203_ 0
C61371 _1012_/a_592_47# _0352_ 0
C61372 _0427_ _0428_ 0.02367f
C61373 _0619_/a_68_297# clknet_1_1__leaf__0458_ 0
C61374 _0296_ _0420_ 0
C61375 hold89/a_49_47# net1 0
C61376 _0660_/a_113_47# _0427_ 0
C61377 _0530_/a_81_21# hold71/a_391_47# 0
C61378 _0530_/a_299_297# hold71/a_285_47# 0
C61379 net119 _0564_/a_68_297# 0.00992f
C61380 _0786_/a_217_297# _0345_ 0.00183f
C61381 _0780_/a_117_297# _0392_ 0
C61382 _0984_/a_466_413# acc0.A\[15\] 0.00548f
C61383 _0137_ _0472_ 0.02229f
C61384 clknet_1_0__leaf__0459_ _1017_/a_381_47# 0.00146f
C61385 pp[16] _0345_ 0
C61386 _0241_ _0462_ 0.00252f
C61387 _0752_/a_300_297# _0237_ 0
C61388 hold87/a_285_47# net165 0
C61389 net25 control0.sh 0.0216f
C61390 VPWR _1028_/a_193_47# 0.28805f
C61391 _1069_/a_634_159# _1069_/a_466_413# 0.23992f
C61392 _1069_/a_193_47# _1069_/a_1059_315# 0.03405f
C61393 _1069_/a_27_47# _1069_/a_891_413# 0.02974f
C61394 net162 _0342_ 0
C61395 _0226_ net46 0
C61396 _0490_ _0170_ 0.03289f
C61397 _0786_/a_300_47# _0295_ 0.0013f
C61398 _0343_ _0773_/a_117_297# 0.00133f
C61399 hold60/a_285_47# hold60/a_391_47# 0.41909f
C61400 _1059_/a_466_413# _0507_/a_27_297# 0
C61401 _0501_/a_27_47# acc0.A\[15\] 0
C61402 acc0.A\[4\] net135 0
C61403 _0328_ _0345_ 0.02418f
C61404 _0954_/a_32_297# _0954_/a_304_297# 0.00167f
C61405 net119 clknet_1_1__leaf_clk 0
C61406 _1037_/a_193_47# comp0.B\[4\] 0
C61407 _0135_ _1036_/a_1059_315# 0
C61408 _0481_ control0.count\[1\] 0.15354f
C61409 _0536_/a_51_297# _0172_ 0.14778f
C61410 _0343_ net76 0
C61411 hold66/a_285_47# _0762_/a_215_47# 0
C61412 _0253_ _0827_/a_109_297# 0
C61413 hold10/a_285_47# _1039_/a_193_47# 0
C61414 hold10/a_391_47# _1039_/a_27_47# 0
C61415 _0180_ _0181_ 0.55042f
C61416 _0255_ _0253_ 0
C61417 net123 clknet_1_1__leaf__0463_ 0.00278f
C61418 _1059_/a_193_47# hold82/a_285_47# 0.00171f
C61419 _1059_/a_27_47# hold82/a_391_47# 0
C61420 comp0.B\[2\] _0956_/a_32_297# 0.14206f
C61421 _0181_ net218 0
C61422 hold37/a_285_47# VPWR 0.3003f
C61423 net62 pp[4] 0.02217f
C61424 _0405_ net5 0.18365f
C61425 hold58/a_391_47# net186 0
C61426 _0985_/a_891_413# _0350_ 0
C61427 control0.state\[2\] _0468_ 0.32144f
C61428 clkbuf_1_1__f__0459_/a_110_47# _0347_ 0
C61429 net247 _0159_ 0
C61430 B[14] _0139_ 0
C61431 _1018_/a_193_47# clkbuf_1_0__f__0461_/a_110_47# 0
C61432 _0084_ _0986_/a_592_47# 0.00124f
C61433 _0218_ _0612_/a_59_75# 0
C61434 _0592_/a_150_297# _0378_ 0
C61435 _0743_/a_51_297# clkbuf_1_0__f__0462_/a_110_47# 0.00803f
C61436 _0217_ _0103_ 0
C61437 _0163_ _0950_/a_75_212# 0
C61438 _0607_/a_109_297# _0181_ 0
C61439 clknet_1_0__leaf__0462_ pp[19] 0
C61440 _0126_ net114 0.08019f
C61441 _0538_/a_51_297# _0538_/a_149_47# 0.02487f
C61442 _0260_ _0846_/a_240_47# 0
C61443 _1037_/a_1059_315# net26 0.00412f
C61444 comp0.B\[3\] _0213_ 0
C61445 clknet_1_1__leaf__0462_ _1008_/a_561_413# 0
C61446 _0715_/a_27_47# _0427_ 0.00919f
C61447 _0532_/a_81_21# acc0.A\[15\] 0
C61448 _0955_/a_32_297# _0132_ 0.00255f
C61449 comp0.B\[6\] _0561_/a_240_47# 0
C61450 _1032_/a_193_47# net201 0
C61451 hold47/a_285_47# _0172_ 0
C61452 comp0.B\[7\] net7 0
C61453 VPWR _1046_/a_975_413# 0.00418f
C61454 VPWR _0798_/a_199_47# 0
C61455 A[10] A[12] 0.18615f
C61456 comp0.B\[13\] net196 0
C61457 _1022_/a_634_159# _1022_/a_592_47# 0
C61458 net123 net8 0
C61459 clkbuf_1_0__f__0463_/a_110_47# clknet_1_1__leaf__0457_ 0.0012f
C61460 _0994_/a_27_47# _0994_/a_1059_315# 0.04875f
C61461 _0994_/a_193_47# _0994_/a_466_413# 0.0802f
C61462 net234 clkbuf_0__0457_/a_110_47# 0
C61463 net207 net1 0
C61464 _1020_/a_27_47# clknet_1_0__leaf__0457_ 0.0438f
C61465 _0108_ net56 0
C61466 _0275_ _0986_/a_1059_315# 0.06357f
C61467 _0272_ _0986_/a_381_47# 0
C61468 _0285_ _0808_/a_266_297# 0.00513f
C61469 _0284_ _0808_/a_81_21# 0.02019f
C61470 _0779_/a_79_21# _0779_/a_510_47# 0.00844f
C61471 _0779_/a_297_297# _0779_/a_215_47# 0
C61472 comp0.B\[10\] _0545_/a_68_297# 0
C61473 net211 _1001_/a_891_413# 0.00251f
C61474 _0473_ _0474_ 0.06335f
C61475 _0472_ comp0.B\[6\] 0.05414f
C61476 _0475_ comp0.B\[5\] 0
C61477 _0289_ _0812_/a_510_47# 0
C61478 input32/a_75_212# net32 0.10849f
C61479 clk _0466_ 0.02224f
C61480 _0179_ _0525_/a_81_21# 0.00234f
C61481 _1055_/a_891_413# _1055_/a_1017_47# 0.00617f
C61482 _1055_/a_193_47# net179 0.31476f
C61483 _1055_/a_634_159# net141 0
C61484 hold88/a_391_47# _0439_ 0
C61485 net247 _0447_ 0
C61486 _0505_/a_373_47# _0184_ 0
C61487 _1023_/a_27_47# output51/a_27_47# 0.00977f
C61488 _0718_/a_47_47# _0216_ 0
C61489 _0995_/a_27_47# _0218_ 0.03618f
C61490 hold88/a_391_47# VPWR 0.17032f
C61491 VPWR _0758_/a_510_47# 0
C61492 _0984_/a_466_413# _0179_ 0
C61493 _0466_ _1063_/a_891_413# 0
C61494 _1003_/a_381_47# _1003_/a_561_413# 0.00123f
C61495 _1003_/a_27_47# net89 0.23152f
C61496 _1003_/a_891_413# _1003_/a_975_413# 0.00851f
C61497 net36 _1047_/a_193_47# 0.14693f
C61498 net166 _0114_ 0.24138f
C61499 _1036_/a_634_159# net27 0
C61500 _1036_/a_381_47# input27/a_75_212# 0
C61501 _0693_/a_68_297# _0324_ 0.05614f
C61502 _0954_/a_32_297# _0540_/a_240_47# 0
C61503 clknet_1_0__leaf__0459_ _0581_/a_27_297# 0
C61504 _0207_ _1040_/a_466_413# 0.0045f
C61505 net171 _1040_/a_1059_315# 0
C61506 hold26/a_49_47# comp0.B\[10\] 0
C61507 _0967_/a_215_297# VPWR 0.36519f
C61508 _0257_ _0346_ 0.02771f
C61509 acc0.A\[14\] clknet_1_0__leaf__0459_ 0.00177f
C61510 _0168_ _0485_ 0
C61511 clknet_1_0__leaf__0460_ hold4/a_391_47# 0
C61512 _0469_ _0467_ 0.00903f
C61513 _0212_ comp0.B\[3\] 0.17727f
C61514 hold46/a_49_47# _0172_ 0.00152f
C61515 VPWR net216 0.66239f
C61516 _0183_ _0856_/a_79_21# 0.01803f
C61517 _0217_ _0856_/a_215_47# 0
C61518 _0257_ net65 0
C61519 _0504_/a_27_47# net68 0
C61520 _0428_ net142 0
C61521 _1004_/a_891_413# _0102_ 0.00561f
C61522 _1004_/a_381_47# _0352_ 0.00745f
C61523 _1004_/a_592_47# _0347_ 0
C61524 net225 net60 0.00455f
C61525 _0852_/a_285_297# acc0.A\[0\] 0
C61526 _0126_ _0365_ 0.002f
C61527 _0983_/a_466_413# _0347_ 0.00368f
C61528 net36 _0459_ 0
C61529 hold56/a_285_47# comp0.B\[2\] 0.01469f
C61530 _0642_/a_27_413# _0399_ 0
C61531 hold91/a_285_47# net42 0
C61532 hold15/a_49_47# acc0.A\[30\] 0
C61533 net23 _1065_/a_1059_315# 0.02348f
C61534 _0330_ _1011_/a_193_47# 0
C61535 net236 clk 0.04126f
C61536 _0799_/a_209_297# _0411_ 0.06201f
C61537 _0626_/a_68_297# _0465_ 0.0015f
C61538 _0765_/a_215_47# hold73/a_391_47# 0
C61539 net68 _0456_ 0
C61540 _1012_/a_891_413# _0350_ 0
C61541 _0195_ _0580_/a_373_47# 0
C61542 _0469_ comp0.B\[0\] 0
C61543 _0500_/a_27_47# _0198_ 0
C61544 _0230_ VPWR 0.14645f
C61545 VPWR _0987_/a_561_413# 0.00342f
C61546 hold23/a_285_47# net175 0.00134f
C61547 hold30/a_49_47# _0225_ 0.00131f
C61548 _1024_/a_634_159# _1024_/a_1059_315# 0
C61549 _1024_/a_27_47# _1024_/a_381_47# 0.06222f
C61550 _1024_/a_193_47# _1024_/a_891_413# 0.19685f
C61551 _1058_/a_592_47# net189 0.0011f
C61552 _0276_ _0403_ 0
C61553 _0811_/a_81_21# _0420_ 0.00222f
C61554 VPWR _0823_/a_109_297# 0.00653f
C61555 hold41/a_285_47# net67 0.01706f
C61556 _0337_ _0707_/a_201_297# 0
C61557 B[9] _1042_/a_193_47# 0.0011f
C61558 _0285_ _0295_ 0
C61559 _1011_/a_634_159# _0333_ 0
C61560 VPWR _0727_/a_277_47# 0
C61561 _0985_/a_193_47# _0180_ 0
C61562 _0284_ _0296_ 0.00141f
C61563 acc0.A\[14\] _0453_ 0
C61564 _0812_/a_79_21# clknet_1_1__leaf__0465_ 0
C61565 _1000_/a_891_413# _0388_ 0.00344f
C61566 VPWR _1029_/a_561_413# 0.00354f
C61567 _0097_ _0240_ 0.0015f
C61568 comp0.B\[2\] _1032_/a_193_47# 0
C61569 _0540_/a_245_297# _0540_/a_240_47# 0
C61570 _0982_/a_381_47# _0453_ 0
C61571 acc0.A\[0\] net247 0
C61572 clk _1064_/a_193_47# 0.00935f
C61573 net9 net132 0
C61574 clkbuf_1_1__f__0460_/a_110_47# _1010_/a_466_413# 0
C61575 _1048_/a_466_413# _1048_/a_561_413# 0.00772f
C61576 _1048_/a_634_159# _1048_/a_975_413# 0
C61577 net53 _0737_/a_35_297# 0
C61578 _1034_/a_1059_315# clknet_1_1__leaf__0463_ 0.01763f
C61579 _0225_ _0352_ 0.02434f
C61580 clknet_1_1__leaf__0464_ net20 0.42127f
C61581 net63 _0522_/a_109_297# 0
C61582 _0348_ pp[28] 0.01299f
C61583 hold48/a_285_47# clknet_1_1__leaf__0464_ 0
C61584 input32/a_75_212# net10 0.00129f
C61585 VPWR _1016_/a_634_159# 0.17807f
C61586 _1068_/a_27_47# _0969_/a_109_297# 0
C61587 net211 _0586_/a_27_47# 0
C61588 net176 _0758_/a_79_21# 0
C61589 _0502_/a_27_47# _0174_ 0
C61590 _0856_/a_79_21# acc0.A\[15\] 0
C61591 _0600_/a_103_199# clkbuf_1_0__f__0460_/a_110_47# 0
C61592 net189 _0186_ 0
C61593 hold11/a_49_47# net158 0.00134f
C61594 _0179_ net37 0.02234f
C61595 _0387_ acc0.A\[17\] 0.00842f
C61596 _0313_ _0330_ 0
C61597 VPWR _0131_ 0.36662f
C61598 net124 _0206_ 0
C61599 net172 comp0.B\[8\] 0
C61600 _1016_/a_27_47# clkbuf_0__0461_/a_110_47# 0.00125f
C61601 clknet_1_0__leaf__0465_ _0147_ 0.00191f
C61602 comp0.B\[14\] _0172_ 0.07052f
C61603 _0670_/a_297_297# acc0.A\[15\] 0.00535f
C61604 _0670_/a_215_47# net42 0.05432f
C61605 _0232_ _0618_/a_79_21# 0.07224f
C61606 _0399_ _0218_ 1.3216f
C61607 net36 _0265_ 0.02235f
C61608 _0230_ net48 0
C61609 _0183_ _0454_ 0
C61610 _0328_ net52 0
C61611 hold33/a_49_47# net7 0.03549f
C61612 _0139_ _0544_/a_51_297# 0.00106f
C61613 net152 _0544_/a_240_47# 0.06744f
C61614 net32 _0544_/a_149_47# 0.00361f
C61615 comp0.B\[1\] _1015_/a_27_47# 0
C61616 pp[30] hold15/a_391_47# 0.01093f
C61617 _1010_/a_891_413# net96 0
C61618 _0130_ _1015_/a_891_413# 0
C61619 net149 acc0.A\[18\] 0
C61620 _1056_/a_193_47# net2 0
C61621 net54 net114 0
C61622 _0315_ net90 0.00405f
C61623 _0599_/a_113_47# net52 0
C61624 _1040_/a_193_47# net174 0.55986f
C61625 _1040_/a_891_413# _1040_/a_1017_47# 0.00617f
C61626 _1053_/a_27_47# acc0.A\[6\] 0
C61627 clknet_1_0__leaf__0465_ _1054_/a_193_47# 0
C61628 hold28/a_285_47# net71 0
C61629 net1 net106 0
C61630 _0748_/a_81_21# _0312_ 0
C61631 _1017_/a_466_413# acc0.A\[18\] 0
C61632 _0979_/a_373_47# _0480_ 0
C61633 _1031_/a_27_47# _0218_ 0
C61634 clknet_1_1__leaf__0465_ _0347_ 0.02405f
C61635 _0527_/a_109_297# net11 0.00922f
C61636 _1072_/a_634_159# _1072_/a_1059_315# 0
C61637 _1072_/a_27_47# _1072_/a_381_47# 0.05761f
C61638 _1072_/a_193_47# _1072_/a_891_413# 0.19421f
C61639 _0216_ _1027_/a_592_47# 0.00188f
C61640 _0830_/a_297_297# _0186_ 0.00462f
C61641 _0279_ _0414_ 0.09365f
C61642 _0513_/a_81_21# net37 0
C61643 _0346_ net11 0
C61644 _0183_ _0505_/a_27_297# 0.09453f
C61645 net30 net127 0
C61646 _0100_ _0183_ 0.02082f
C61647 VPWR _1019_/a_975_413# 0.00416f
C61648 _0714_/a_149_47# VPWR 0
C61649 _0313_ _0732_/a_209_297# 0.03624f
C61650 _0172_ _0543_/a_68_297# 0
C61651 net1 _0237_ 0
C61652 hold68/a_49_47# _0758_/a_79_21# 0
C61653 _0195_ _0309_ 0
C61654 acc0.A\[14\] _0996_/a_1017_47# 0.0011f
C61655 comp0.B\[5\] net27 0
C61656 _1067_/a_891_413# _1067_/a_1017_47# 0.00617f
C61657 _0244_ _1018_/a_1059_315# 0
C61658 net44 hold95/a_285_47# 0
C61659 _0429_ net65 0.23695f
C61660 _0251_ _0989_/a_891_413# 0.03698f
C61661 _0429_ _0989_/a_466_413# 0
C61662 _0412_ _0410_ 0.00234f
C61663 _0343_ clkbuf_0__0459_/a_110_47# 0.00286f
C61664 _0154_ A[10] 0.09411f
C61665 _0538_/a_51_297# clkbuf_0__0464_/a_110_47# 0.00781f
C61666 _1071_/a_381_47# _0169_ 0.11472f
C61667 _0985_/a_27_47# net10 0
C61668 _0702_/a_113_47# _0333_ 0
C61669 hold90/a_391_47# _0219_ 0.00289f
C61670 _1004_/a_193_47# _0380_ 0
C61671 _1004_/a_634_159# _0350_ 0
C61672 VPWR _0116_ 0.7072f
C61673 _0693_/a_68_297# _0347_ 0
C61674 control0.state\[1\] _1002_/a_381_47# 0
C61675 _0252_ _0989_/a_975_413# 0
C61676 _0989_/a_1059_315# _0989_/a_1017_47# 0
C61677 _0502_/a_27_47# _0208_ 0
C61678 VPWR _0807_/a_150_297# 0.00195f
C61679 hold75/a_49_47# hold86/a_285_47# 0
C61680 _0997_/a_634_159# _0997_/a_1059_315# 0
C61681 _0997_/a_27_47# _0997_/a_381_47# 0.05761f
C61682 _0997_/a_193_47# _0997_/a_891_413# 0.19226f
C61683 _1037_/a_27_47# input24/a_75_212# 0
C61684 clknet_1_0__leaf__0462_ net176 0.06869f
C61685 _0454_ acc0.A\[15\] 0
C61686 _0544_/a_149_47# _1042_/a_1059_315# 0
C61687 _0181_ _0986_/a_381_47# 0
C61688 _0372_ _0247_ 0
C61689 _0992_/a_1059_315# _0992_/a_1017_47# 0
C61690 VPWR _1051_/a_1059_315# 0.40948f
C61691 _0498_/a_240_47# acc0.A\[15\] 0
C61692 net26 _0561_/a_240_47# 0
C61693 _0312_ clknet_0__0462_ 0.002f
C61694 net78 hold81/a_391_47# 0
C61695 _0183_ _0506_/a_81_21# 0
C61696 _0236_ VPWR 0.59696f
C61697 hold6/a_285_47# _1042_/a_193_47# 0
C61698 hold6/a_391_47# _1042_/a_27_47# 0
C61699 VPWR _1045_/a_381_47# 0.07545f
C61700 net158 _0159_ 0
C61701 VPWR net139 0.37455f
C61702 net54 _0365_ 0.02892f
C61703 net89 hold93/a_285_47# 0
C61704 clknet_0__0458_ _0841_/a_510_47# 0
C61705 _0109_ _1029_/a_891_413# 0
C61706 control0.reset _1061_/a_891_413# 0
C61707 net100 acc0.A\[0\] 0.00384f
C61708 hold13/a_285_47# _0474_ 0.00139f
C61709 hold63/a_49_47# VPWR 0.32862f
C61710 _0192_ acc0.A\[6\] 0
C61711 clkbuf_0__0463_/a_110_47# _0171_ 0.02118f
C61712 _1045_/a_27_47# net129 0
C61713 _0793_/a_51_297# _0400_ 0.00108f
C61714 net243 _0756_/a_47_47# 0
C61715 _0743_/a_245_297# _0105_ 0
C61716 _1027_/a_27_47# _1027_/a_466_413# 0.27314f
C61717 _1027_/a_193_47# _1027_/a_634_159# 0.11897f
C61718 _0558_/a_150_297# comp0.B\[4\] 0
C61719 _0253_ _0830_/a_215_47# 0
C61720 hold46/a_285_47# hold26/a_391_47# 0.01305f
C61721 hold46/a_391_47# hold26/a_285_47# 0.00232f
C61722 _0285_ _0811_/a_299_297# 0
C61723 acc0.A\[15\] _0505_/a_27_297# 0.0147f
C61724 _0996_/a_27_47# net41 0.00849f
C61725 _0465_ _1061_/a_1059_315# 0.00966f
C61726 hold54/a_391_47# net201 0.13136f
C61727 _1061_/a_193_47# _1061_/a_592_47# 0.00135f
C61728 _1061_/a_634_159# _1061_/a_975_413# 0
C61729 _1061_/a_466_413# _1061_/a_561_413# 0.00772f
C61730 A[13] _0300_ 0
C61731 _0955_/a_32_297# net25 0
C61732 net51 _0754_/a_240_47# 0.00129f
C61733 hold98/a_49_47# _0341_ 0
C61734 net66 _0990_/a_891_413# 0.03749f
C61735 acc0.A\[8\] _0990_/a_1059_315# 0.0098f
C61736 _0291_ _0990_/a_466_413# 0
C61737 net160 B[5] 0
C61738 clkbuf_1_0__f__0457_/a_110_47# hold40/a_49_47# 0.01705f
C61739 net155 net112 0
C61740 _1007_/a_975_413# _0219_ 0
C61741 _1054_/a_466_413# A[4] 0
C61742 _0136_ comp0.B\[5\] 0
C61743 _0313_ net190 0
C61744 _0399_ _0833_/a_215_47# 0.00223f
C61745 _1035_/a_634_159# _1035_/a_466_413# 0.23992f
C61746 _1035_/a_193_47# _1035_/a_1059_315# 0.03384f
C61747 _1035_/a_27_47# _1035_/a_891_413# 0.03224f
C61748 _0734_/a_129_47# _0219_ 0
C61749 net105 _0526_/a_27_47# 0
C61750 _0279_ _0300_ 0
C61751 _0959_/a_472_297# _1065_/a_193_47# 0
C61752 clknet_1_0__leaf__0462_ hold68/a_49_47# 0.00918f
C61753 _0416_ _0414_ 0
C61754 hold75/a_285_47# acc0.A\[14\] 0
C61755 _0118_ acc0.A\[20\] 0.06981f
C61756 _0477_ _0955_/a_32_297# 0.01206f
C61757 _0217_ _1014_/a_1017_47# 0
C61758 _0489_ _1069_/a_891_413# 0.02725f
C61759 _0983_/a_27_47# _0849_/a_79_21# 0
C61760 output60/a_27_47# pp[31] 0.15785f
C61761 _1013_/a_193_47# clknet_1_1__leaf__0461_ 0
C61762 net113 _0320_ 0
C61763 net101 _0208_ 0.08342f
C61764 comp0.B\[1\] _0215_ 0
C61765 net211 net149 0.0044f
C61766 net48 _0236_ 0.0049f
C61767 _0222_ _0374_ 0.46918f
C61768 _0195_ clknet_1_1__leaf__0457_ 0.7743f
C61769 hold11/a_285_47# net134 0
C61770 net76 _0990_/a_381_47# 0
C61771 _0299_ _0218_ 0.03478f
C61772 hold20/a_285_47# _0466_ 0
C61773 acc0.A\[15\] _0506_/a_81_21# 0.00448f
C61774 acc0.A\[29\] _1029_/a_193_47# 0.0039f
C61775 _0268_ _0636_/a_145_75# 0.00134f
C61776 clknet_1_0__leaf__0459_ _1016_/a_634_159# 0
C61777 _1069_/a_634_159# _0167_ 0.00178f
C61778 _1069_/a_466_413# clknet_1_0__leaf_clk 0.00176f
C61779 _1056_/a_891_413# net66 0.00264f
C61780 hold98/a_285_47# _1013_/a_1059_315# 0
C61781 _0343_ output65/a_27_47# 0
C61782 VPWR _0422_ 0.36875f
C61783 _0854_/a_510_47# _0181_ 0.00447f
C61784 _0349_ net59 0
C61785 _0337_ pp[30] 0.0104f
C61786 _0384_ hold73/a_285_47# 0
C61787 VPWR B[7] 0.26523f
C61788 _0500_/a_27_47# net247 0.04509f
C61789 hold74/a_49_47# _0781_/a_68_297# 0.01017f
C61790 _1059_/a_975_413# acc0.A\[13\] 0
C61791 _1059_/a_466_413# _0185_ 0.00175f
C61792 VPWR _0534_/a_384_47# 0
C61793 pp[8] _1055_/a_466_413# 0
C61794 _0399_ _0112_ 0
C61795 _0233_ _0600_/a_337_297# 0.00312f
C61796 _0231_ _0600_/a_253_297# 0
C61797 VPWR hold62/a_391_47# 0.1742f
C61798 _0181_ _0498_/a_51_297# 0
C61799 net36 _0267_ 0
C61800 _1041_/a_891_413# _1040_/a_891_413# 0
C61801 _1015_/a_193_47# _0721_/a_27_47# 0.00125f
C61802 _1031_/a_1017_47# _0220_ 0.00207f
C61803 _0997_/a_891_413# _0411_ 0
C61804 hold10/a_49_47# net125 0
C61805 pp[8] net181 0.04263f
C61806 _0990_/a_891_413# _0350_ 0
C61807 clknet_1_0__leaf__0460_ _1063_/a_1059_315# 0
C61808 _0346_ clknet_1_1__leaf__0458_ 0.02583f
C61809 hold19/a_285_47# _0219_ 0
C61810 _1027_/a_381_47# _1026_/a_27_47# 0
C61811 _0846_/a_51_297# acc0.A\[15\] 0.00317f
C61812 _0179_ _0505_/a_27_297# 0
C61813 _0533_/a_109_297# _0171_ 0
C61814 _0176_ net18 0.02795f
C61815 _1002_/a_1017_47# _0181_ 0
C61816 _0490_ net35 0
C61817 _0183_ _1022_/a_1059_315# 0
C61818 acc0.A\[22\] _1022_/a_891_413# 0.02141f
C61819 net65 clknet_1_1__leaf__0458_ 0.01994f
C61820 hold57/a_391_47# _0210_ 0.00281f
C61821 _0343_ _1006_/a_193_47# 0
C61822 clknet_1_1__leaf__0458_ _0989_/a_466_413# 0
C61823 _0538_/a_240_47# net21 0.0646f
C61824 VPWR _0760_/a_377_297# 0.00595f
C61825 clknet_1_0__leaf__0463_ _0498_/a_149_47# 0.00227f
C61826 _0121_ VPWR 0.36269f
C61827 _0474_ _0132_ 0.02244f
C61828 hold20/a_285_47# net236 0
C61829 _0271_ acc0.A\[6\] 0
C61830 pp[25] _0572_/a_373_47# 0
C61831 output53/a_27_47# net155 0
C61832 net23 hold93/a_49_47# 0
C61833 _0482_ clkbuf_1_0__f_clk/a_110_47# 0
C61834 _0343_ _0986_/a_193_47# 0
C61835 _0325_ _0693_/a_150_297# 0
C61836 _0987_/a_891_413# acc0.A\[6\] 0
C61837 _0987_/a_27_47# _0193_ 0
C61838 hold64/a_285_47# _0580_/a_109_297# 0
C61839 hold64/a_391_47# _0580_/a_27_297# 0
C61840 _0579_/a_27_297# _1019_/a_27_47# 0
C61841 net199 _1025_/a_975_413# 0
C61842 _0994_/a_891_413# _0994_/a_1017_47# 0.00617f
C61843 _0285_ _0091_ 0.20206f
C61844 _0579_/a_109_297# _0099_ 0
C61845 _0500_/a_27_47# _1048_/a_466_413# 0
C61846 _0891_/a_27_47# clknet_1_0__leaf__0461_ 0
C61847 _0311_ _0216_ 0
C61848 _0972_/a_93_21# _0972_/a_346_47# 0.01191f
C61849 hold56/a_391_47# _0215_ 0
C61850 _1023_/a_381_47# pp[23] 0
C61851 _1023_/a_975_413# net51 0
C61852 _0423_ _0990_/a_1059_315# 0
C61853 _0401_ _0990_/a_634_159# 0
C61854 _0346_ _0263_ 0
C61855 _0781_/a_150_297# net43 0
C61856 net234 _0350_ 0.07435f
C61857 _0966_/a_109_297# _0484_ 0
C61858 _0415_ _0277_ 0
C61859 _1003_/a_1017_47# _0101_ 0.00109f
C61860 _0752_/a_300_297# _0222_ 0.06239f
C61861 _0179_ _0506_/a_81_21# 0.06615f
C61862 A[5] acc0.A\[6\] 0
C61863 hold37/a_49_47# _0172_ 0
C61864 _0279_ _0404_ 0.0731f
C61865 _0399_ _0099_ 0
C61866 _0993_/a_634_159# _0993_/a_1059_315# 0
C61867 _0993_/a_27_47# _0993_/a_381_47# 0.06222f
C61868 _0993_/a_193_47# _0993_/a_891_413# 0.19685f
C61869 _0816_/a_150_297# _0656_/a_59_75# 0
C61870 _1058_/a_466_413# _0156_ 0
C61871 _0182_ net201 0
C61872 clknet_1_0__leaf__0459_ _0116_ 0
C61873 hold45/a_285_47# net144 0.07653f
C61874 _0207_ net174 0
C61875 _0149_ net135 0
C61876 _1039_/a_466_413# _1039_/a_561_413# 0.00772f
C61877 _1039_/a_634_159# _1039_/a_975_413# 0
C61878 _0180_ _0531_/a_27_297# 0.10217f
C61879 _0182_ _0531_/a_109_297# 0.04351f
C61880 hold67/a_49_47# _0369_ 0.04831f
C61881 hold33/a_391_47# _0138_ 0.03576f
C61882 _0197_ net10 0.01752f
C61883 _1020_/a_592_47# _0457_ 0
C61884 hold32/a_49_47# acc0.A\[9\] 0.01974f
C61885 _0785_/a_81_21# clknet_0__0465_ 0.0272f
C61886 net46 _0350_ 0.17216f
C61887 net175 hold71/a_285_47# 0.00137f
C61888 _0578_/a_373_47# net1 0.00174f
C61889 _0663_/a_27_413# _0289_ 0.04046f
C61890 output55/a_27_47# clknet_1_1__leaf__0460_ 0
C61891 _0996_/a_193_47# _0400_ 0.00223f
C61892 _0736_/a_56_297# _0371_ 0
C61893 _0172_ _1046_/a_561_413# 0.00127f
C61894 _0179_ _0846_/a_51_297# 0.03412f
C61895 _1049_/a_466_413# _0148_ 0
C61896 _0465_ _0631_/a_109_297# 0
C61897 _0393_ acc0.A\[18\] 0
C61898 net26 B[4] 0.02368f
C61899 _1026_/a_1059_315# _1026_/a_891_413# 0.31086f
C61900 _1026_/a_193_47# _1026_/a_975_413# 0
C61901 _1026_/a_466_413# _1026_/a_381_47# 0.03733f
C61902 hold74/a_285_47# _0369_ 0
C61903 net33 _1062_/a_1017_47# 0
C61904 net39 acc0.A\[12\] 0.44513f
C61905 _0551_/a_27_47# control0.sh 0.08846f
C61906 _0286_ _0807_/a_68_297# 0
C61907 net140 _1053_/a_1017_47# 0
C61908 net88 _0467_ 0
C61909 _0222_ _0249_ 0.04477f
C61910 _0629_/a_145_75# _0261_ 0.00124f
C61911 _0629_/a_59_75# _0263_ 0.03476f
C61912 acc0.A\[2\] _0631_/a_109_297# 0.00285f
C61913 _0720_/a_68_297# _0720_/a_150_297# 0.00477f
C61914 _0337_ _0717_/a_80_21# 0
C61915 _0430_ _0433_ 0.00737f
C61916 _1024_/a_1059_315# net110 0
C61917 _1024_/a_466_413# _0122_ 0.00473f
C61918 _0225_ _0237_ 0
C61919 _1024_/a_27_47# acc0.A\[24\] 0
C61920 VPWR _0370_ 1.22043f
C61921 _0337_ _0339_ 0.00128f
C61922 _1014_/a_1059_315# _0181_ 0
C61923 net97 _0333_ 0
C61924 _0278_ _0646_/a_129_47# 0
C61925 _0083_ acc0.A\[1\] 0
C61926 net67 net4 0.02373f
C61927 net61 _0255_ 0.04132f
C61928 _0821_/a_113_47# net168 0
C61929 _1057_/a_634_159# net143 0
C61930 _0439_ acc0.A\[8\] 0.05999f
C61931 acc0.A\[5\] _0433_ 0.47966f
C61932 net104 acc0.A\[1\] 0
C61933 pp[16] _0997_/a_193_47# 0
C61934 net45 _0386_ 0
C61935 _0949_/a_59_75# clknet_1_1__leaf_clk 0.00474f
C61936 hold89/a_49_47# control0.count\[1\] 0
C61937 net2 clknet_1_1__leaf__0465_ 0.29608f
C61938 VPWR acc0.A\[8\] 0.99648f
C61939 _0276_ acc0.A\[13\] 0.22861f
C61940 _0469_ net1 0.12231f
C61941 _0209_ net8 0
C61942 _0356_ _0568_/a_109_297# 0
C61943 _0957_/a_32_297# net24 0.04178f
C61944 _0831_/a_285_47# _0434_ 0.00159f
C61945 _0346_ clknet_1_0__leaf__0461_ 0.08101f
C61946 _0533_/a_27_297# control0.sh 0
C61947 _1020_/a_466_413# _0208_ 0
C61948 _1041_/a_634_159# _1041_/a_466_413# 0.23992f
C61949 _1041_/a_193_47# _1041_/a_1059_315# 0.03324f
C61950 _1041_/a_27_47# _1041_/a_891_413# 0.02996f
C61951 _0624_/a_145_75# _0256_ 0
C61952 VPWR _0991_/a_193_47# 0.32825f
C61953 hold99/a_391_47# _0993_/a_193_47# 0
C61954 net167 clkbuf_0_clk/a_110_47# 0
C61955 clknet_1_0__leaf__0460_ net93 0.00731f
C61956 _1059_/a_466_413# _0289_ 0
C61957 _0504_/a_27_47# hold71/a_49_47# 0.0861f
C61958 VPWR _0773_/a_285_47# 0
C61959 acc0.A\[27\] _0317_ 0.15353f
C61960 _0217_ _0764_/a_81_21# 0.00136f
C61961 _0340_ net60 0.15518f
C61962 _1015_/a_381_47# comp0.B\[15\] 0
C61963 init B[0] 0.128f
C61964 _0682_/a_68_297# _0216_ 0
C61965 _1002_/a_634_159# net1 0
C61966 _0416_ _0404_ 0.27885f
C61967 _0274_ _0825_/a_150_297# 0
C61968 net31 hold6/a_49_47# 0
C61969 hold54/a_49_47# VPWR 0.26396f
C61970 _0551_/a_27_47# net157 0
C61971 acc0.A\[16\] acc0.A\[17\] 0.17804f
C61972 clknet_0__0464_ _1061_/a_1059_315# 0
C61973 pp[2] acc0.A\[6\] 0.00276f
C61974 hold86/a_49_47# _0345_ 0
C61975 net163 _0336_ 0.21395f
C61976 clknet_0__0460_ _1006_/a_891_413# 0.00168f
C61977 _0707_/a_201_297# _0333_ 0.01124f
C61978 _0369_ _0610_/a_59_75# 0.04544f
C61979 hold44/a_391_47# _1029_/a_634_159# 0
C61980 hold44/a_49_47# _1029_/a_1059_315# 0
C61981 hold44/a_285_47# _1029_/a_466_413# 0.0041f
C61982 clknet_0__0458_ _0627_/a_369_297# 0
C61983 _0422_ _0283_ 0.076f
C61984 _0752_/a_27_413# _0762_/a_215_47# 0
C61985 net63 _0150_ 0
C61986 VPWR _0380_ 0.67122f
C61987 output58/a_27_47# _0827_/a_27_47# 0
C61988 _0444_ _0445_ 0.1568f
C61989 _0183_ _0184_ 0
C61990 _0284_ _0652_/a_109_297# 0.01263f
C61991 net186 clkbuf_1_1__f__0463_/a_110_47# 0.00487f
C61992 _0317_ _0364_ 0
C61993 _0330_ _0321_ 0
C61994 clkbuf_1_0__f__0459_/a_110_47# clkbuf_0__0459_/a_110_47# 0
C61995 _0399_ net228 0
C61996 _0081_ _0583_/a_109_47# 0
C61997 _1013_/a_381_47# net60 0
C61998 VPWR _1025_/a_975_413# 0.0052f
C61999 _0293_ _0991_/a_891_413# 0
C62000 _0661_/a_205_297# _0089_ 0
C62001 _0573_/a_27_47# clknet_1_1__leaf__0457_ 0.00168f
C62002 _0391_ _0345_ 0
C62003 _0462_ _0352_ 0.04392f
C62004 _0254_ _0252_ 0.16698f
C62005 _0743_/a_51_297# _0324_ 0
C62006 _0743_/a_245_297# _0359_ 0.00394f
C62007 _0533_/a_27_297# net157 0
C62008 _0625_/a_59_75# _0836_/a_150_297# 0
C62009 net105 _1015_/a_592_47# 0
C62010 _1012_/a_27_47# _0351_ 0.00194f
C62011 net64 _0439_ 0
C62012 acc0.A\[4\] _0172_ 0.03356f
C62013 net22 _0540_/a_51_297# 0
C62014 clknet_1_1__leaf__0460_ _1006_/a_1017_47# 0
C62015 _0225_ _1005_/a_27_47# 0
C62016 net64 VPWR 0.96107f
C62017 _0643_/a_103_199# _0084_ 0
C62018 _0275_ _0841_/a_79_21# 0
C62019 _1051_/a_1059_315# _0523_/a_81_21# 0
C62020 net155 net111 0
C62021 VPWR _0621_/a_117_297# 0.00729f
C62022 _0190_ _0833_/a_215_47# 0
C62023 _1059_/a_27_47# clknet_1_1__leaf__0465_ 0
C62024 _0195_ _0570_/a_109_47# 0.00179f
C62025 _0216_ _0570_/a_27_297# 0.17659f
C62026 _0107_ _0359_ 0
C62027 _0595_/a_109_297# clknet_1_0__leaf__0460_ 0
C62028 acc0.A\[3\] _0529_/a_27_297# 0.02428f
C62029 _1053_/a_891_413# _0150_ 0
C62030 hold11/a_285_47# net22 0
C62031 _0285_ _0346_ 0.20855f
C62032 _0460_ hold93/a_391_47# 0.02109f
C62033 _0140_ _1042_/a_891_413# 0
C62034 net198 _1042_/a_592_47# 0.00105f
C62035 net18 _1042_/a_975_413# 0
C62036 VPWR _1044_/a_891_413# 0.18445f
C62037 _0198_ _1049_/a_27_47# 0
C62038 clknet_1_0__leaf__0462_ _0605_/a_109_297# 0
C62039 acc0.A\[14\] _0345_ 0.03417f
C62040 hold100/a_285_47# _0219_ 0
C62041 VPWR _0423_ 0.44371f
C62042 _0349_ _1010_/a_592_47# 0.00143f
C62043 _0683_/a_113_47# VPWR 0
C62044 clkbuf_1_0__f__0459_/a_110_47# _1059_/a_381_47# 0
C62045 _0732_/a_209_47# _0360_ 0.00201f
C62046 _0608_/a_27_47# net43 0
C62047 _0470_ hold84/a_49_47# 0.00106f
C62048 _0398_ _0347_ 0.00342f
C62049 _0960_/a_27_47# _0979_/a_27_297# 0.01248f
C62050 _0218_ _0091_ 0.00545f
C62051 _0756_/a_47_47# _0378_ 0.37469f
C62052 _0407_ _0408_ 0.18126f
C62053 _1001_/a_891_413# _0461_ 0.00741f
C62054 _0786_/a_472_297# _0421_ 0
C62055 net36 _0178_ 0.0196f
C62056 _1027_/a_27_47# net156 0.10162f
C62057 _1027_/a_1059_315# _1027_/a_1017_47# 0
C62058 _0643_/a_337_297# _0643_/a_253_47# 0.00219f
C62059 output44/a_27_47# _0341_ 0
C62060 net44 _0710_/a_381_47# 0
C62061 _0764_/a_299_297# control0.add 0
C62062 clknet_1_1__leaf__0459_ _0341_ 0
C62063 hold8/a_391_47# clknet_1_1__leaf__0462_ 0.00372f
C62064 _0547_/a_68_297# _1040_/a_27_47# 0.01172f
C62065 acc0.A\[15\] _0184_ 0.01124f
C62066 hold11/a_285_47# clknet_1_0__leaf__0463_ 0
C62067 hold89/a_285_47# control0.count\[2\] 0
C62068 VPWR _1032_/a_1017_47# 0
C62069 _0464_ _1051_/a_27_47# 0
C62070 _0362_ _0308_ 0
C62071 _0231_ _0222_ 0.2774f
C62072 clknet_1_0__leaf__0465_ acc0.A\[6\] 0.00835f
C62073 net101 _1019_/a_193_47# 0
C62074 _0749_/a_81_21# _0749_/a_384_47# 0.00138f
C62075 clknet_1_0__leaf__0462_ _1023_/a_466_413# 0.00239f
C62076 net46 _0244_ 0.00214f
C62077 net206 acc0.A\[18\] 0.1238f
C62078 net64 output62/a_27_47# 0.01391f
C62079 net169 A[4] 0
C62080 _0195_ hold50/a_391_47# 0
C62081 _0216_ hold50/a_49_47# 0
C62082 net133 _1061_/a_193_47# 0
C62083 clknet_1_0__leaf__0464_ _1061_/a_466_413# 0
C62084 net70 net165 0
C62085 clkload2/a_268_47# net135 0
C62086 clknet_0__0458_ _0274_ 0.12637f
C62087 hold20/a_391_47# hold12/a_391_47# 0
C62088 control0.reset _1063_/a_193_47# 0
C62089 _0991_/a_1059_315# clknet_1_1__leaf__0465_ 0.00445f
C62090 _1035_/a_634_159# _0133_ 0.06295f
C62091 _1035_/a_466_413# net121 0.00141f
C62092 acc0.A\[27\] net197 0.04552f
C62093 _0389_ clkbuf_1_0__f__0461_/a_110_47# 0.00194f
C62094 _0248_ _0764_/a_81_21# 0
C62095 _0358_ _0729_/a_150_297# 0
C62096 hold39/a_49_47# _1034_/a_466_413# 0.01477f
C62097 hold39/a_391_47# _1034_/a_193_47# 0.00108f
C62098 hold39/a_285_47# _1034_/a_634_159# 0.0021f
C62099 _1058_/a_27_47# _1058_/a_634_159# 0.14145f
C62100 _0446_ _0843_/a_68_297# 0.04579f
C62101 _0218_ _0306_ 0
C62102 _0329_ _0690_/a_68_297# 0.03327f
C62103 _0322_ _0690_/a_150_297# 0.00105f
C62104 input23/a_75_212# net23 0.11037f
C62105 _0946_/a_30_53# _1064_/a_1059_315# 0.01627f
C62106 _0277_ _0347_ 0
C62107 _0312_ _0747_/a_215_47# 0
C62108 _0477_ _0474_ 0
C62109 _1051_/a_466_413# _0172_ 0.03398f
C62110 net124 A[1] 0.00137f
C62111 _0410_ _0669_/a_183_297# 0
C62112 _0172_ _1045_/a_891_413# 0
C62113 _0983_/a_193_47# _0082_ 0
C62114 _0343_ _0103_ 0
C62115 _1030_/a_1059_315# _0334_ 0
C62116 clknet_1_1__leaf__0459_ _1013_/a_891_413# 0
C62117 _0680_/a_80_21# _0680_/a_217_297# 0.12661f
C62118 _0310_ _0780_/a_35_297# 0.04742f
C62119 _0718_/a_47_47# _0337_ 0.06437f
C62120 _1054_/a_1017_47# acc0.A\[8\] 0
C62121 _1011_/a_27_47# _0354_ 0.0295f
C62122 _0343_ hold91/a_391_47# 0.00286f
C62123 _0243_ _0632_/a_113_47# 0
C62124 _1069_/a_1017_47# control0.count\[0\] 0
C62125 clknet_1_0__leaf_clk _0167_ 0.28752f
C62126 clknet_1_0__leaf__0465_ _0523_/a_384_47# 0
C62127 _1033_/a_634_159# _1065_/a_891_413# 0
C62128 net32 _1043_/a_466_413# 0
C62129 _1030_/a_27_47# _0351_ 0
C62130 _0182_ _1015_/a_193_47# 0
C62131 _0157_ _0185_ 0.25552f
C62132 _0966_/a_27_47# _0482_ 0.04087f
C62133 _1052_/a_634_159# net148 0
C62134 _0316_ hold77/a_49_47# 0
C62135 net55 hold77/a_285_47# 0.08595f
C62136 pp[8] net179 0.02685f
C62137 _0160_ hold84/a_391_47# 0.01031f
C62138 net190 _0321_ 0
C62139 net197 _0364_ 0
C62140 _0432_ _0438_ 0.00235f
C62141 _0457_ control0.reset 0
C62142 _0179_ _0524_/a_109_297# 0.00462f
C62143 net45 _0342_ 0.001f
C62144 net125 _1061_/a_975_413# 0
C62145 _0734_/a_285_47# _0318_ 0.05235f
C62146 _0398_ _1016_/a_891_413# 0
C62147 net150 _0183_ 0.31399f
C62148 _0217_ acc0.A\[22\] 0.25811f
C62149 comp0.B\[10\] _1061_/a_193_47# 0
C62150 net156 _1026_/a_466_413# 0
C62151 _1027_/a_27_47# acc0.A\[26\] 0.08673f
C62152 hold65/a_285_47# _0369_ 0.02164f
C62153 _0195_ _1018_/a_1059_315# 0.04537f
C62154 _0553_/a_240_47# net171 0.05177f
C62155 net58 _0988_/a_1059_315# 0
C62156 _0179_ _0184_ 0.17055f
C62157 hold77/a_49_47# _0347_ 0.00132f
C62158 net1 net220 0
C62159 _0467_ _1067_/a_891_413# 0
C62160 _0128_ hold62/a_49_47# 0.31186f
C62161 hold97/a_49_47# _0319_ 0
C62162 hold20/a_285_47# clkload0/X 0
C62163 hold15/a_285_47# net162 0.00972f
C62164 _1038_/a_193_47# _0176_ 0.03713f
C62165 _0343_ net57 0.03008f
C62166 _0563_/a_512_297# _0208_ 0.00334f
C62167 _0461_ _0586_/a_27_47# 0.00365f
C62168 _0530_/a_81_21# _1048_/a_27_47# 0
C62169 net202 _0566_/a_27_47# 0
C62170 hold59/a_49_47# net206 0.04248f
C62171 hold58/a_285_47# _1034_/a_1059_315# 0.00341f
C62172 _0996_/a_193_47# clkbuf_0__0459_/a_110_47# 0.00398f
C62173 _0295_ net228 0.11844f
C62174 net59 _1012_/a_193_47# 0.00325f
C62175 output66/a_27_47# output67/a_27_47# 0
C62176 B[10] B[11] 0.18036f
C62177 _1065_/a_975_413# _0160_ 0
C62178 net49 _0228_ 0.02471f
C62179 _0403_ _0993_/a_27_47# 0
C62180 _0801_/a_113_47# net80 0
C62181 _1037_/a_27_47# net121 0
C62182 comp0.B\[11\] _0203_ 0.01753f
C62183 _0954_/a_32_297# _0141_ 0
C62184 net89 _0974_/a_448_47# 0
C62185 net211 _1019_/a_891_413# 0.01233f
C62186 _0995_/a_193_47# pp[14] 0.00552f
C62187 _0183_ _0580_/a_373_47# 0.00127f
C62188 net30 B[7] 0.00981f
C62189 _0137_ input30/a_75_212# 0
C62190 _0982_/a_592_47# net36 0.00253f
C62191 _0520_/a_109_47# net168 0
C62192 net55 _0107_ 0
C62193 _0538_/a_245_297# _0174_ 0
C62194 _0343_ _0670_/a_510_47# 0
C62195 VPWR _1042_/a_27_47# 0.40119f
C62196 _0425_ clknet_1_1__leaf__0465_ 0
C62197 net61 _0830_/a_215_47# 0
C62198 clknet_1_0__leaf__0465_ _0624_/a_59_75# 0
C62199 net58 _0635_/a_27_47# 0.00103f
C62200 net45 _1013_/a_592_47# 0
C62201 hold91/a_285_47# net5 0.04434f
C62202 _0179_ _1048_/a_592_47# 0.00107f
C62203 _0684_/a_59_75# _0219_ 0.00286f
C62204 pp[30] _0333_ 0
C62205 _0518_/a_27_297# hold1/a_285_47# 0
C62206 _1043_/a_891_413# _1042_/a_634_159# 0
C62207 _1043_/a_1059_315# _1042_/a_466_413# 0
C62208 _1043_/a_634_159# _1042_/a_891_413# 0
C62209 _1043_/a_466_413# _1042_/a_1059_315# 0
C62210 _0290_ _0088_ 0.00492f
C62211 _0458_ net71 0.03377f
C62212 net116 hold92/a_391_47# 0
C62213 _1055_/a_381_47# net74 0
C62214 _0386_ VPWR 0.24898f
C62215 _0642_/a_27_413# net65 0.0444f
C62216 _0642_/a_298_297# _0989_/a_193_47# 0
C62217 _0426_ acc0.A\[9\] 0.24585f
C62218 _0988_/a_27_47# _0988_/a_193_47# 0.9705f
C62219 net178 acc0.A\[10\] 0
C62220 pp[27] _1030_/a_466_413# 0
C62221 _0269_ _0840_/a_68_297# 0
C62222 _0342_ _0587_/a_27_47# 0
C62223 hold6/a_285_47# clknet_1_1__leaf__0464_ 0
C62224 _0352_ _0754_/a_245_297# 0.00234f
C62225 _0437_ pp[3] 0
C62226 _0255_ _0431_ 0.37042f
C62227 _0984_/a_193_47# _0983_/a_193_47# 0
C62228 output45/a_27_47# _1013_/a_1059_315# 0
C62229 _0751_/a_183_297# net46 0
C62230 _0730_/a_215_47# _0730_/a_510_47# 0.00529f
C62231 clknet_1_1__leaf__0460_ _1010_/a_634_159# 0
C62232 acc0.A\[29\] hold95/a_391_47# 0.03137f
C62233 comp0.B\[2\] _0495_/a_68_297# 0
C62234 _0146_ _0197_ 0.00419f
C62235 net10 _1043_/a_466_413# 0
C62236 _0456_ _0264_ 0.11375f
C62237 hold21/a_285_47# hold22/a_49_47# 0.01404f
C62238 _0296_ _0347_ 0.02224f
C62239 _0501_/a_27_47# _0171_ 0.01646f
C62240 _0266_ clkbuf_1_0__f__0461_/a_110_47# 0
C62241 _0475_ control0.reset 0.00606f
C62242 _0542_/a_51_297# _0542_/a_245_297# 0.01218f
C62243 _0147_ _0148_ 0
C62244 _0162_ _1064_/a_634_159# 0.00226f
C62245 _0485_ _1064_/a_891_413# 0.00583f
C62246 _0487_ _1064_/a_1059_315# 0
C62247 hold92/a_285_47# hold92/a_391_47# 0.41909f
C62248 pp[9] net141 0
C62249 hold52/a_285_47# _0123_ 0.00557f
C62250 _0747_/a_510_47# _0219_ 0
C62251 _1026_/a_466_413# acc0.A\[26\] 0.0012f
C62252 _1059_/a_975_413# VPWR 0.00493f
C62253 _0465_ _1047_/a_381_47# 0.00187f
C62254 _0480_ control0.state\[2\] 0
C62255 _0472_ _0465_ 0
C62256 _0376_ _0103_ 0.01594f
C62257 _0322_ _0359_ 0
C62258 _0472_ _1061_/a_381_47# 0
C62259 net76 acc0.A\[6\] 0.00195f
C62260 clknet_1_1__leaf__0460_ _1009_/a_466_413# 0.01294f
C62261 _0590_/a_113_47# VPWR 0
C62262 acc0.A\[19\] _0771_/a_298_297# 0
C62263 _1020_/a_891_413# _0099_ 0
C62264 hold65/a_49_47# _0825_/a_68_297# 0.01354f
C62265 _0327_ _0359_ 0.03359f
C62266 _0203_ _0202_ 0.00253f
C62267 _0542_/a_240_47# net20 0.0461f
C62268 _0183_ control0.add 0.02552f
C62269 net122 control0.sh 0
C62270 _0346_ _0218_ 0.10968f
C62271 _0423_ _0283_ 0.00273f
C62272 _0982_/a_27_47# hold60/a_49_47# 0
C62273 pp[26] _0571_/a_109_297# 0.04911f
C62274 net59 clknet_1_1__leaf__0461_ 0
C62275 _0966_/a_27_47# hold89/a_285_47# 0
C62276 hold76/a_285_47# _0241_ 0.03194f
C62277 net24 _0213_ 0.02638f
C62278 _0789_/a_208_47# _0405_ 0.00108f
C62279 _0850_/a_150_297# _0465_ 0
C62280 _0230_ _0345_ 0.13489f
C62281 _0273_ _0437_ 0.00194f
C62282 _0736_/a_311_297# _0370_ 0
C62283 clknet_1_1__leaf__0459_ net37 0.06474f
C62284 _0680_/a_80_21# _0372_ 0
C62285 _0174_ _1040_/a_561_413# 0
C62286 _0136_ _1040_/a_634_159# 0
C62287 net65 _0218_ 0
C62288 _1037_/a_466_413# _1037_/a_561_413# 0.00772f
C62289 _1037_/a_634_159# _1037_/a_975_413# 0
C62290 input15/a_75_212# net12 0
C62291 _0345_ _0823_/a_109_297# 0
C62292 _0123_ net52 0.00942f
C62293 net186 _0163_ 0
C62294 _0199_ acc0.A\[3\] 0
C62295 _0195_ _0998_/a_27_47# 0.4218f
C62296 _0217_ _0379_ 0
C62297 _0606_/a_215_297# clknet_1_0__leaf__0460_ 0
C62298 net58 _0850_/a_68_297# 0
C62299 _0369_ acc0.A\[13\] 0.14656f
C62300 _0259_ clknet_1_1__leaf__0458_ 0
C62301 net59 _1030_/a_193_47# 0.00176f
C62302 _0184_ VGND 0.28208f
C62303 net6 VGND 0.48242f
C62304 _0505_/a_373_47# VGND 0.00233f 
C62305 _0505_/a_109_47# VGND 0.00618f 
C62306 _0505_/a_109_297# VGND 0.00396f 
C62307 _0505_/a_27_297# VGND 0.4303f 
C62308 pp[5] VGND 0.69989f
C62309 output63/a_27_47# VGND 0.72343f 
C62310 pp[14] VGND 0.66508f
C62311 net41 VGND 1.26745f
C62312 output41/a_27_47# VGND 0.46752f 
C62313 pp[24] VGND 1.03933f
C62314 net52 VGND 1.52166f
C62315 output52/a_27_47# VGND 0.45056f 
C62316 _0103_ VGND 0.93818f
C62317 net91 VGND 0.49112f
C62318 _1005_/a_1017_47# VGND 0.00538f 
C62319 _1005_/a_592_47# VGND 0.00748f 
C62320 _1005_/a_975_413# VGND 0 
C62321 _1005_/a_381_47# VGND 0.06688f 
C62322 _1005_/a_891_413# VGND 0.31218f 
C62323 _1005_/a_1059_315# VGND 0.46643f 
C62324 _1005_/a_466_413# VGND 0.23949f 
C62325 _1005_/a_634_159# VGND 0.28101f 
C62326 _1005_/a_193_47# VGND 0.37718f 
C62327 _1005_/a_27_47# VGND 0.65741f 
C62328 _0193_ VGND 0.74301f
C62329 net13 VGND 0.58443f
C62330 acc0.A\[6\] VGND 1.73282f
C62331 _0522_/a_373_47# VGND 0.00212f 
C62332 _0522_/a_109_47# VGND 0.00618f 
C62333 _0522_/a_109_297# VGND 0.0045f 
C62334 _0522_/a_27_297# VGND 0.43259f 
C62335 hold95/a_391_47# VGND 0.23989f 
C62336 hold95/a_285_47# VGND 0.39167f 
C62337 hold95/a_49_47# VGND 0.43302f 
C62338 hold84/a_391_47# VGND 0.30089f 
C62339 hold84/a_285_47# VGND 0.4469f 
C62340 hold84/a_49_47# VGND 0.48845f 
C62341 hold73/a_391_47# VGND 0.25651f 
C62342 hold73/a_285_47# VGND 0.45238f 
C62343 hold73/a_49_47# VGND 0.47989f 
C62344 net209 VGND 0.36025f
C62345 hold62/a_391_47# VGND 0.27699f 
C62346 hold62/a_285_47# VGND 0.4174f 
C62347 hold62/a_49_47# VGND 0.44916f 
C62348 hold51/a_391_47# VGND 0.23636f 
C62349 hold51/a_285_47# VGND 0.395f 
C62350 hold51/a_49_47# VGND 0.4322f 
C62351 hold40/a_391_47# VGND 0.26447f 
C62352 hold40/a_285_47# VGND 0.45159f 
C62353 hold40/a_49_47# VGND 0.50555f 
C62354 _0599_/a_113_47# VGND 0.00175f 
C62355 _0418_ VGND 0.16435f
C62356 _0281_ VGND 1.87646f
C62357 _0806_/a_199_47# VGND 0.00372f 
C62358 _0806_/a_113_297# VGND 0.03749f 
C62359 _0364_ VGND 0.46834f
C62360 _0321_ VGND 0.76252f
C62361 _0360_ VGND 1.53564f
C62362 _0737_/a_285_47# VGND 0.00505f 
C62363 _0737_/a_285_297# VGND 0.0033f 
C62364 _0737_/a_117_297# VGND 0.00135f 
C62365 _0737_/a_35_297# VGND 0.41895f 
C62366 _0668_/a_297_47# VGND 0.20501f 
C62367 _0668_/a_382_297# VGND 0 
C62368 _0668_/a_79_21# VGND 0.31403f 
C62369 net151 VGND 0.46f
C62370 _1022_/a_1017_47# VGND 0.00416f 
C62371 _1022_/a_592_47# VGND 0.01038f 
C62372 _1022_/a_975_413# VGND 0 
C62373 _1022_/a_561_413# VGND 0.00225f 
C62374 _1022_/a_381_47# VGND 0.07948f 
C62375 _1022_/a_891_413# VGND 0.27884f 
C62376 _1022_/a_1059_315# VGND 0.38979f 
C62377 _1022_/a_466_413# VGND 0.24858f 
C62378 _1022_/a_634_159# VGND 0.27718f 
C62379 _1022_/a_193_47# VGND 0.47813f 
C62380 _1022_/a_27_47# VGND 0.64553f 
C62381 _0685_/a_150_297# VGND 0 
C62382 _0685_/a_68_297# VGND 0.2696f 
C62383 _0431_ VGND 0.90603f
C62384 _0823_/a_109_297# VGND 0 
C62385 _0219_ VGND 8.78613f
C62386 net241 VGND 0.45056f
C62387 _0377_ VGND 0.20722f
C62388 _0345_ VGND 8.87126f
C62389 _0754_/a_240_47# VGND 0.16489f 
C62390 _0754_/a_149_47# VGND 0.12844f 
C62391 _0754_/a_512_297# VGND 0 
C62392 _0754_/a_245_297# VGND 0 
C62393 _0754_/a_51_297# VGND 0.28536f 
C62394 _0468_ VGND 1.43269f
C62395 _0969_/a_109_297# VGND 0 
C62396 _0840_/a_150_297# VGND 0 
C62397 _0840_/a_68_297# VGND 0.26457f 
C62398 _0771_/a_382_47# VGND 0.00573f 
C62399 _0771_/a_298_297# VGND 0.00487f 
C62400 _0771_/a_215_297# VGND 0.41854f 
C62401 _0771_/a_27_413# VGND 0.26798f 
C62402 _0986_/a_1017_47# VGND 0.00404f 
C62403 _0986_/a_592_47# VGND 0.00662f 
C62404 _0986_/a_381_47# VGND 0.06058f 
C62405 _0986_/a_891_413# VGND 0.27437f 
C62406 _0986_/a_1059_315# VGND 0.38405f 
C62407 _0986_/a_466_413# VGND 0.21103f 
C62408 _0986_/a_634_159# VGND 0.25514f 
C62409 _0986_/a_193_47# VGND 0.34412f 
C62410 _0986_/a_27_47# VGND 0.55526f 
C62411 net229 VGND 0.99612f
C62412 _0506_/a_384_47# VGND 0.00449f 
C62413 _0506_/a_299_297# VGND 0.05298f 
C62414 _0506_/a_81_21# VGND 0.33083f 
C62415 pp[4] VGND 0.6728f
C62416 output62/a_27_47# VGND 0.69998f 
C62417 pp[13] VGND 0.63369f
C62418 output40/a_27_47# VGND 0.44281f 
C62419 pp[23] VGND 0.95614f
C62420 net51 VGND 3.65958f
C62421 output51/a_27_47# VGND 0.45219f 
C62422 net92 VGND 0.58201f
C62423 _1006_/a_1017_47# VGND 0.00404f 
C62424 _1006_/a_592_47# VGND 0.00662f 
C62425 _1006_/a_381_47# VGND 0.06019f 
C62426 _1006_/a_891_413# VGND 0.27462f 
C62427 _1006_/a_1059_315# VGND 0.38308f 
C62428 _1006_/a_466_413# VGND 0.21067f 
C62429 _1006_/a_634_159# VGND 0.25177f 
C62430 _1006_/a_193_47# VGND 0.34999f 
C62431 _1006_/a_27_47# VGND 0.57763f 
C62432 _0150_ VGND 0.3217f
C62433 _0523_/a_384_47# VGND 0.00325f 
C62434 _0523_/a_299_297# VGND 0.04097f 
C62435 _0523_/a_81_21# VGND 0.30997f 
C62436 hold94/a_391_47# VGND 0.23875f 
C62437 hold94/a_285_47# VGND 0.40864f 
C62438 hold94/a_49_47# VGND 0.45054f 
C62439 hold83/a_391_47# VGND 0.24151f 
C62440 hold83/a_285_47# VGND 0.39909f 
C62441 hold83/a_49_47# VGND 0.43471f 
C62442 hold72/a_391_47# VGND 0.2609f 
C62443 hold72/a_285_47# VGND 0.44005f 
C62444 hold72/a_49_47# VGND 0.46715f 
C62445 hold61/a_391_47# VGND 0.24139f 
C62446 hold61/a_285_47# VGND 0.3966f 
C62447 hold61/a_49_47# VGND 0.46739f 
C62448 hold50/a_391_47# VGND 0.24283f 
C62449 hold50/a_285_47# VGND 0.39598f 
C62450 hold50/a_49_47# VGND 0.46318f 
C62451 _0301_ VGND 0.61014f
C62452 _0669_/a_183_297# VGND 0 
C62453 _0669_/a_111_297# VGND 0 
C62454 _0669_/a_29_53# VGND 0.4468f 
C62455 net244 VGND 0.3443f
C62456 _0738_/a_150_297# VGND 0 
C62457 _0738_/a_68_297# VGND 0.27171f 
C62458 net246 VGND 0.86085f
C62459 _0807_/a_150_297# VGND 0.00202f 
C62460 _0807_/a_68_297# VGND 0.32138f 
C62461 acc0.A\[23\] VGND 2.29102f
C62462 net177 VGND 0.51672f
C62463 net109 VGND 0.89768f
C62464 _1023_/a_1017_47# VGND 0.00463f 
C62465 _1023_/a_592_47# VGND 0.00778f 
C62466 _1023_/a_975_413# VGND 0 
C62467 _1023_/a_561_413# VGND 0 
C62468 _1023_/a_381_47# VGND 0.06747f 
C62469 _1023_/a_891_413# VGND 0.29613f 
C62470 _1023_/a_1059_315# VGND 0.41731f 
C62471 _1023_/a_466_413# VGND 0.22242f 
C62472 _1023_/a_634_159# VGND 0.27f 
C62473 _1023_/a_193_47# VGND 0.45377f 
C62474 _1023_/a_27_47# VGND 0.64654f 
C62475 _0142_ VGND 0.55687f
C62476 net20 VGND 2.03586f
C62477 _0202_ VGND 0.68234f
C62478 _0540_/a_240_47# VGND 0.1914f 
C62479 _0540_/a_149_47# VGND 0.13364f 
C62480 _0540_/a_512_297# VGND 0.00312f 
C62481 _0540_/a_245_297# VGND 0.00101f 
C62482 _0540_/a_51_297# VGND 0.33661f 
C62483 net142 VGND 0.59934f
C62484 _0318_ VGND 0.89262f
C62485 _0686_/a_301_297# VGND 0 
C62486 _0686_/a_27_53# VGND 0.32171f 
C62487 _0686_/a_219_297# VGND 0.26418f 
C62488 _0374_ VGND 0.56613f
C62489 _0755_/a_109_297# VGND 0 
C62490 _0824_/a_145_75# VGND 0.00486f 
C62491 _0824_/a_59_75# VGND 0.32499f 
C62492 net174 VGND 0.30776f
C62493 _1040_/a_1017_47# VGND 0.00404f 
C62494 _1040_/a_592_47# VGND 0.00662f 
C62495 _1040_/a_975_413# VGND 0 
C62496 _1040_/a_561_413# VGND 0 
C62497 _1040_/a_381_47# VGND 0.06105f 
C62498 _1040_/a_891_413# VGND 0.27674f 
C62499 _1040_/a_1059_315# VGND 0.39188f 
C62500 _1040_/a_466_413# VGND 0.21056f 
C62501 _1040_/a_634_159# VGND 0.25258f 
C62502 _1040_/a_193_47# VGND 0.34472f 
C62503 _1040_/a_27_47# VGND 0.5682f 
C62504 _0084_ VGND 0.47725f
C62505 _0445_ VGND 0.4609f
C62506 _0444_ VGND 0.4469f
C62507 _0841_/a_510_47# VGND 0.00785f 
C62508 _0841_/a_215_47# VGND 0.23529f 
C62509 _0841_/a_79_21# VGND 0.39324f 
C62510 _0099_ VGND 0.4906f
C62511 _0391_ VGND 0.19916f
C62512 net223 VGND 0.3221f
C62513 _0772_/a_510_47# VGND 0.00683f 
C62514 _0772_/a_215_47# VGND 0.22873f 
C62515 _0772_/a_297_297# VGND 0 
C62516 _0772_/a_79_21# VGND 0.3513f 
C62517 net75 VGND 0.32956f
C62518 _0085_ VGND 0.7164f
C62519 net73 VGND 0.33571f
C62520 _0987_/a_1017_47# VGND 0.00447f 
C62521 _0987_/a_592_47# VGND 0.00748f 
C62522 _0987_/a_975_413# VGND 0 
C62523 _0987_/a_381_47# VGND 0.06538f 
C62524 _0987_/a_891_413# VGND 0.28669f 
C62525 _0987_/a_1059_315# VGND 0.39475f 
C62526 _0987_/a_466_413# VGND 0.21748f 
C62527 _0987_/a_634_159# VGND 0.25846f 
C62528 _0987_/a_193_47# VGND 0.36503f 
C62529 _0987_/a_27_47# VGND 0.59589f 
C62530 _0185_ VGND 0.70691f
C62531 net5 VGND 1.40079f
C62532 acc0.A\[13\] VGND 3.37823f
C62533 _0507_/a_373_47# VGND 0.003f 
C62534 _0507_/a_109_47# VGND 0.00767f 
C62535 _0507_/a_109_297# VGND 0.00274f 
C62536 _0507_/a_27_297# VGND 0.43819f 
C62537 pp[3] VGND 0.62777f
C62538 output61/a_27_47# VGND 0.70873f 
C62539 pp[22] VGND 0.95063f
C62540 net50 VGND 2.70399f
C62541 output50/a_27_47# VGND 0.47758f 
C62542 _0105_ VGND 0.44428f
C62543 net93 VGND 0.6303f
C62544 _1007_/a_1017_47# VGND 0.00525f 
C62545 _1007_/a_592_47# VGND 0.00786f 
C62546 _1007_/a_975_413# VGND 0 
C62547 _1007_/a_561_413# VGND 0 
C62548 _1007_/a_381_47# VGND 0.06233f 
C62549 _1007_/a_891_413# VGND 0.31367f 
C62550 _1007_/a_1059_315# VGND 0.44273f 
C62551 _1007_/a_466_413# VGND 0.23107f 
C62552 _1007_/a_634_159# VGND 0.28155f 
C62553 _1007_/a_193_47# VGND 0.37358f 
C62554 _1007_/a_27_47# VGND 0.627f 
C62555 _0194_ VGND 0.24603f
C62556 net12 VGND 0.5414f
C62557 net148 VGND 0.54515f
C62558 _0524_/a_373_47# VGND 0.00288f 
C62559 _0524_/a_109_47# VGND 0.00753f 
C62560 _0524_/a_109_297# VGND 0.00274f 
C62561 _0524_/a_27_297# VGND 0.43632f 
C62562 hold93/a_391_47# VGND 0.23718f 
C62563 hold93/a_285_47# VGND 0.39241f 
C62564 hold93/a_49_47# VGND 0.43149f 
C62565 hold82/a_391_47# VGND 0.25613f 
C62566 hold82/a_285_47# VGND 0.45967f 
C62567 hold82/a_49_47# VGND 0.5291f 
C62568 net218 VGND 0.50327f
C62569 hold71/a_391_47# VGND 0.25196f 
C62570 hold71/a_285_47# VGND 0.40948f 
C62571 hold71/a_49_47# VGND 0.44755f 
C62572 hold60/a_391_47# VGND 0.24213f 
C62573 hold60/a_285_47# VGND 0.40217f 
C62574 hold60/a_49_47# VGND 0.43284f 
C62575 _0106_ VGND 0.58453f
C62576 _0365_ VGND 0.44927f
C62577 _0739_/a_510_47# VGND 0.00585f 
C62578 _0739_/a_215_47# VGND 0.22445f 
C62579 _0739_/a_79_21# VGND 0.37479f 
C62580 _0091_ VGND 0.49038f
C62581 _0419_ VGND 0.41644f
C62582 _0417_ VGND 0.3741f
C62583 _0808_/a_585_47# VGND 0 
C62584 _0808_/a_266_47# VGND 0.19308f 
C62585 _0808_/a_266_297# VGND 0 
C62586 _0808_/a_81_21# VGND 0.34618f 
C62587 acc0.A\[24\] VGND 1.12405f
C62588 _0122_ VGND 0.447f
C62589 net110 VGND 0.4592f
C62590 _1024_/a_1017_47# VGND 0.00447f 
C62591 _1024_/a_592_47# VGND 0.00748f 
C62592 _1024_/a_975_413# VGND 0 
C62593 _1024_/a_381_47# VGND 0.06714f 
C62594 _1024_/a_891_413# VGND 0.29277f 
C62595 _1024_/a_1059_315# VGND 0.42771f 
C62596 _1024_/a_466_413# VGND 0.22436f 
C62597 _1024_/a_634_159# VGND 0.27599f 
C62598 _1024_/a_193_47# VGND 0.47803f 
C62599 _1024_/a_27_47# VGND 0.64962f 
C62600 _0541_/a_150_297# VGND 0 
C62601 _0541_/a_68_297# VGND 0.27856f 
C62602 _0242_ VGND 2.03551f
C62603 acc0.A\[19\] VGND 1.19012f
C62604 _0610_/a_145_75# VGND 0.00334f 
C62605 _0610_/a_59_75# VGND 0.31556f 
C62606 _0379_ VGND 0.20513f
C62607 _0378_ VGND 0.78748f
C62608 _0756_/a_285_47# VGND 0.21282f 
C62609 _0756_/a_129_47# VGND 0.0043f 
C62610 _0756_/a_377_297# VGND 0 
C62611 _0756_/a_47_47# VGND 0.31372f 
C62612 _0687_/a_145_75# VGND 0.00514f 
C62613 _0687_/a_59_75# VGND 0.31339f 
C62614 _0825_/a_150_297# VGND 0 
C62615 _0825_/a_68_297# VGND 0.27267f 
C62616 comp0.B\[9\] VGND 1.76356f
C62617 net153 VGND 0.41793f
C62618 net127 VGND 0.62327f
C62619 _1041_/a_1017_47# VGND 0.00482f 
C62620 _1041_/a_592_47# VGND 0.007f 
C62621 _1041_/a_975_413# VGND 0 
C62622 _1041_/a_561_413# VGND 0 
C62623 _1041_/a_381_47# VGND 0.06301f 
C62624 _1041_/a_891_413# VGND 0.28656f 
C62625 _1041_/a_1059_315# VGND 0.4001f 
C62626 _1041_/a_466_413# VGND 0.21593f 
C62627 _1041_/a_634_159# VGND 0.2584f 
C62628 _1041_/a_193_47# VGND 0.3675f 
C62629 _1041_/a_27_47# VGND 0.57489f 
C62630 _0392_ VGND 0.41106f
C62631 _0773_/a_285_47# VGND 0.00475f 
C62632 _0773_/a_285_297# VGND 0.01008f 
C62633 _0773_/a_117_297# VGND 0 
C62634 _0773_/a_35_297# VGND 0.44665f 
C62635 _0842_/a_145_75# VGND 0.00487f 
C62636 _0842_/a_59_75# VGND 0.32252f 
C62637 net90 VGND 0.43517f
C62638 net74 VGND 0.32269f
C62639 _0988_/a_1017_47# VGND 0.00422f 
C62640 _0988_/a_592_47# VGND 0.00688f 
C62641 _0988_/a_975_413# VGND 0 
C62642 _0988_/a_561_413# VGND 0 
C62643 _0988_/a_381_47# VGND 0.06195f 
C62644 _0988_/a_891_413# VGND 0.29635f 
C62645 _0988_/a_1059_315# VGND 0.40975f 
C62646 _0988_/a_466_413# VGND 0.23313f 
C62647 _0988_/a_634_159# VGND 0.26988f 
C62648 _0988_/a_193_47# VGND 0.37656f 
C62649 _0988_/a_27_47# VGND 0.59118f 
C62650 _0406_ VGND 0.44575f
C62651 acc0.A\[15\] VGND 5.07806f
C62652 net42 VGND 1.67696f
C62653 _0790_/a_285_47# VGND 0.00424f 
C62654 _0790_/a_285_297# VGND 0.00153f 
C62655 _0790_/a_35_297# VGND 0.4329f 
C62656 net228 VGND 1.40008f
C62657 _0508_/a_384_47# VGND 0.00397f 
C62658 _0508_/a_299_297# VGND 0.0492f 
C62659 _0508_/a_81_21# VGND 0.33866f 
C62660 pp[31] VGND 0.52283f
C62661 output60/a_27_47# VGND 0.43544f 
C62662 net94 VGND 0.60791f
C62663 _1008_/a_1017_47# VGND 0.00494f 
C62664 _1008_/a_592_47# VGND 0.00815f 
C62665 _1008_/a_975_413# VGND 0 
C62666 _1008_/a_561_413# VGND 0 
C62667 _1008_/a_381_47# VGND 0.06918f 
C62668 _1008_/a_891_413# VGND 0.29523f 
C62669 _1008_/a_1059_315# VGND 0.40949f 
C62670 _1008_/a_466_413# VGND 0.22395f 
C62671 _1008_/a_634_159# VGND 0.27089f 
C62672 _1008_/a_193_47# VGND 0.38014f 
C62673 _1008_/a_27_47# VGND 0.64529f 
C62674 _0525_/a_384_47# VGND 0.00368f 
C62675 _0525_/a_299_297# VGND 0.04009f 
C62676 _0525_/a_81_21# VGND 0.32639f 
C62677 hold92/a_391_47# VGND 0.25571f 
C62678 hold92/a_285_47# VGND 0.41914f 
C62679 hold92/a_49_47# VGND 0.46139f 
C62680 hold81/a_391_47# VGND 0.2558f 
C62681 hold81/a_285_47# VGND 0.42315f 
C62682 hold81/a_49_47# VGND 0.4852f 
C62683 net37 VGND 1.60265f
C62684 hold70/a_391_47# VGND 0.24533f 
C62685 hold70/a_285_47# VGND 0.40512f 
C62686 hold70/a_49_47# VGND 0.4391f 
C62687 _0420_ VGND 0.57488f
C62688 _0809_/a_384_47# VGND 0.00329f 
C62689 _0809_/a_299_297# VGND 0.04102f 
C62690 _0809_/a_81_21# VGND 0.31848f 
C62691 acc0.A\[25\] VGND 2.9917f
C62692 _1025_/a_1017_47# VGND 0.00415f 
C62693 _1025_/a_592_47# VGND 0.00909f 
C62694 _1025_/a_975_413# VGND 0 
C62695 _1025_/a_561_413# VGND 0.00264f 
C62696 _1025_/a_381_47# VGND 0.06911f 
C62697 _1025_/a_891_413# VGND 0.29792f 
C62698 _1025_/a_1059_315# VGND 0.41681f 
C62699 _1025_/a_466_413# VGND 0.25907f 
C62700 _1025_/a_634_159# VGND 0.28143f 
C62701 _1025_/a_193_47# VGND 0.39608f 
C62702 _1025_/a_27_47# VGND 0.63254f 
C62703 _0611_/a_150_297# VGND 0 
C62704 _0611_/a_68_297# VGND 0.27242f 
C62705 _0141_ VGND 0.28337f
C62706 net19 VGND 0.33244f
C62707 net195 VGND 0.5078f
C62708 _0203_ VGND 0.55296f
C62709 _0542_/a_240_47# VGND 0.16117f 
C62710 _0542_/a_149_47# VGND 0.125f 
C62711 _0542_/a_51_297# VGND 0.27188f 
C62712 _0320_ VGND 0.50268f
C62713 _0688_/a_109_297# VGND 0 
C62714 _0380_ VGND 0.26373f
C62715 _0350_ VGND 8.39509f
C62716 _0757_/a_150_297# VGND 0 
C62717 _0757_/a_68_297# VGND 0.26126f 
C62718 _0434_ VGND 0.78414f
C62719 _0826_/a_301_297# VGND 0 
C62720 _0826_/a_27_53# VGND 0.34202f 
C62721 _0826_/a_219_297# VGND 0.26027f 
C62722 net128 VGND 0.53851f
C62723 _1042_/a_1017_47# VGND 0.00447f 
C62724 _1042_/a_592_47# VGND 0.00748f 
C62725 _1042_/a_975_413# VGND 0 
C62726 _1042_/a_381_47# VGND 0.06538f 
C62727 _1042_/a_891_413# VGND 0.28336f 
C62728 _1042_/a_1059_315# VGND 0.40856f 
C62729 _1042_/a_466_413# VGND 0.2178f 
C62730 _1042_/a_634_159# VGND 0.25851f 
C62731 _1042_/a_193_47# VGND 0.35007f 
C62732 _1042_/a_27_47# VGND 0.56269f 
C62733 _0774_/a_150_297# VGND 0 
C62734 _0774_/a_68_297# VGND 0.27032f 
C62735 _0843_/a_150_297# VGND 0 
C62736 _0843_/a_68_297# VGND 0.26878f 
C62737 clkbuf_0__0457_/a_110_47# VGND 2.29179f 
C62738 _0989_/a_1017_47# VGND 0.00447f 
C62739 _0989_/a_592_47# VGND 0.00863f 
C62740 _0989_/a_975_413# VGND 0 
C62741 _0989_/a_561_413# VGND 0.00108f 
C62742 _0989_/a_381_47# VGND 0.06441f 
C62743 _0989_/a_891_413# VGND 0.28476f 
C62744 _0989_/a_1059_315# VGND 0.39386f 
C62745 _0989_/a_466_413# VGND 0.22629f 
C62746 _0989_/a_634_159# VGND 0.27611f 
C62747 _0989_/a_193_47# VGND 0.36687f 
C62748 _0989_/a_27_47# VGND 0.61027f 
C62749 _0791_/a_199_47# VGND 0.00382f 
C62750 _0791_/a_113_297# VGND 0.03855f 
C62751 _0186_ VGND 4.18527f
C62752 _0509_/a_27_47# VGND 0.43529f 
C62753 _1009_/a_1017_47# VGND 0.00415f 
C62754 _1009_/a_592_47# VGND 0.00772f 
C62755 _1009_/a_975_413# VGND 0 
C62756 _1009_/a_561_413# VGND 0 
C62757 _1009_/a_381_47# VGND 0.07155f 
C62758 _1009_/a_891_413# VGND 0.28969f 
C62759 _1009_/a_1059_315# VGND 0.42255f 
C62760 _1009_/a_466_413# VGND 0.24318f 
C62761 _1009_/a_634_159# VGND 0.26992f 
C62762 _1009_/a_193_47# VGND 0.44618f 
C62763 _1009_/a_27_47# VGND 0.65508f 
C62764 _0526_/a_27_47# VGND 0.72837f 
C62765 hold91/a_391_47# VGND 0.25285f 
C62766 hold91/a_285_47# VGND 0.44319f 
C62767 hold91/a_49_47# VGND 0.46962f 
C62768 hold80/a_391_47# VGND 0.26117f 
C62769 hold80/a_285_47# VGND 0.42909f 
C62770 hold80/a_49_47# VGND 0.46395f 
C62771 acc0.A\[26\] VGND 1.1428f
C62772 net112 VGND 0.33872f
C62773 _1026_/a_1017_47# VGND 0.00454f 
C62774 _1026_/a_592_47# VGND 0.00773f 
C62775 _1026_/a_975_413# VGND 0 
C62776 _1026_/a_561_413# VGND 0 
C62777 _1026_/a_381_47# VGND 0.06091f 
C62778 _1026_/a_891_413# VGND 0.28395f 
C62779 _1026_/a_1059_315# VGND 0.39266f 
C62780 _1026_/a_466_413# VGND 0.22686f 
C62781 _1026_/a_634_159# VGND 0.27766f 
C62782 _1026_/a_193_47# VGND 0.46159f 
C62783 _1026_/a_27_47# VGND 0.58483f 
C62784 _0543_/a_150_297# VGND 0 
C62785 _0543_/a_68_297# VGND 0.27308f 
C62786 acc0.A\[18\] VGND 1.39142f
C62787 _0612_/a_145_75# VGND 0.0048f 
C62788 _0612_/a_59_75# VGND 0.29914f 
C62789 _0319_ VGND 0.81969f
C62790 _0689_/a_150_297# VGND 0 
C62791 _0689_/a_68_297# VGND 0.27911f 
C62792 _0102_ VGND 0.49288f
C62793 _0352_ VGND 7.32117f
C62794 _0347_ VGND 8.86814f
C62795 _0758_/a_510_47# VGND 0.00955f 
C62796 _0758_/a_215_47# VGND 0.23982f 
C62797 _0758_/a_297_297# VGND 0 
C62798 _0758_/a_79_21# VGND 0.38513f 
C62799 _0827_/a_27_47# VGND 0.17584f 
C62800 _0827_/a_109_297# VGND 0 
C62801 net196 VGND 0.30834f
C62802 net129 VGND 0.3064f
C62803 _1043_/a_1017_47# VGND 0.00447f 
C62804 _1043_/a_592_47# VGND 0.00748f 
C62805 _1043_/a_381_47# VGND 0.06684f 
C62806 _1043_/a_891_413# VGND 0.28795f 
C62807 _1043_/a_1059_315# VGND 0.39712f 
C62808 _1043_/a_466_413# VGND 0.21978f 
C62809 _1043_/a_634_159# VGND 0.26583f 
C62810 _1043_/a_193_47# VGND 0.35524f 
C62811 _1043_/a_27_47# VGND 0.59847f 
C62812 _0560_/a_150_297# VGND 0 
C62813 _0560_/a_68_297# VGND 0.27185f 
C62814 _0393_ VGND 0.41525f
C62815 _0775_/a_510_47# VGND 0.00733f 
C62816 _0775_/a_215_47# VGND 0.2197f 
C62817 _0775_/a_79_21# VGND 0.37455f 
C62818 _0913_/a_27_47# VGND 0.31018f 
C62819 _0448_ VGND 0.52535f
C62820 _0447_ VGND 0.46717f
C62821 _0844_/a_297_47# VGND 0.20882f 
C62822 _0844_/a_382_297# VGND 0 
C62823 _0844_/a_79_21# VGND 0.28792f 
C62824 _0158_ VGND 0.4623f
C62825 net146 VGND 0.43543f
C62826 _1060_/a_1017_47# VGND 0.0048f 
C62827 _1060_/a_592_47# VGND 0.00797f 
C62828 _1060_/a_975_413# VGND 0 
C62829 _1060_/a_561_413# VGND 0 
C62830 _1060_/a_381_47# VGND 0.06673f 
C62831 _1060_/a_891_413# VGND 0.29807f 
C62832 _1060_/a_1059_315# VGND 0.38745f 
C62833 _1060_/a_466_413# VGND 0.23635f 
C62834 _1060_/a_634_159# VGND 0.30211f 
C62835 _1060_/a_193_47# VGND 0.39195f 
C62836 _1060_/a_27_47# VGND 0.636f 
C62837 clkbuf_0__0458_/a_110_47# VGND 2.28002f 
C62838 _0408_ VGND 0.23009f
C62839 _0400_ VGND 1.70001f
C62840 _0405_ VGND 1.0976f
C62841 _0792_/a_303_47# VGND 0.00505f 
C62842 _0792_/a_209_47# VGND 0.00544f 
C62843 _0792_/a_209_297# VGND 0.00621f 
C62844 _0792_/a_80_21# VGND 0.39847f 
C62845 net11 VGND 0.61511f
C62846 net154 VGND 0.62333f
C62847 _0527_/a_373_47# VGND 0.00288f 
C62848 _0527_/a_109_47# VGND 0.00753f 
C62849 _0527_/a_109_297# VGND 0.00274f 
C62850 _0527_/a_27_297# VGND 0.4483f 
C62851 hold90/a_391_47# VGND 0.27953f 
C62852 hold90/a_285_47# VGND 0.41768f 
C62853 hold90/a_49_47# VGND 0.43992f 
C62854 net156 VGND 0.27512f
C62855 _1027_/a_1017_47# VGND 0.00447f 
C62856 _1027_/a_592_47# VGND 0.00748f 
C62857 _1027_/a_381_47# VGND 0.06538f 
C62858 _1027_/a_891_413# VGND 0.28256f 
C62859 _1027_/a_1059_315# VGND 0.40588f 
C62860 _1027_/a_466_413# VGND 0.21743f 
C62861 _1027_/a_634_159# VGND 0.25845f 
C62862 _1027_/a_193_47# VGND 0.35027f 
C62863 _1027_/a_27_47# VGND 0.56258f 
C62864 net113 VGND 0.31316f
C62865 clknet_1_1__leaf__0462_ VGND 4.45105f
C62866 _0140_ VGND 0.35082f
C62867 net18 VGND 1.51038f
C62868 net198 VGND 0.2833f
C62869 _0204_ VGND 0.27091f
C62870 _0544_/a_240_47# VGND 0.16839f 
C62871 _0544_/a_149_47# VGND 0.12594f 
C62872 _0544_/a_512_297# VGND 0 
C62873 _0544_/a_245_297# VGND 0 
C62874 _0544_/a_51_297# VGND 0.28162f 
C62875 _0613_/a_109_297# VGND 0 
C62876 net72 VGND 0.31571f
C62877 clknet_1_1__leaf__0458_ VGND 3.91855f
C62878 _0436_ VGND 0.16827f
C62879 _0435_ VGND 0.44121f
C62880 _0828_/a_199_47# VGND 0.00414f 
C62881 _0828_/a_113_297# VGND 0.04256f 
C62882 _0373_ VGND 1.0534f
C62883 _0759_/a_113_47# VGND 0.00181f 
C62884 net79 VGND 0.42617f
C62885 net130 VGND 0.80853f
C62886 _1044_/a_1017_47# VGND 0.00531f 
C62887 _1044_/a_592_47# VGND 0.00748f 
C62888 _1044_/a_975_413# VGND 0 
C62889 _1044_/a_561_413# VGND 0 
C62890 _1044_/a_381_47# VGND 0.06213f 
C62891 _1044_/a_891_413# VGND 0.29978f 
C62892 _1044_/a_1059_315# VGND 0.43185f 
C62893 _1044_/a_466_413# VGND 0.21271f 
C62894 _1044_/a_634_159# VGND 0.25967f 
C62895 _1044_/a_193_47# VGND 0.35177f 
C62896 _1044_/a_27_47# VGND 0.57585f 
C62897 _0630_/a_109_297# VGND 0.00164f 
C62898 _0492_/a_27_47# VGND 0.40275f 
C62899 _0132_ VGND 0.3387f
C62900 _0208_ VGND 4.51375f
C62901 _0173_ VGND 2.48759f
C62902 _0213_ VGND 0.47788f
C62903 _0561_/a_240_47# VGND 0.16542f 
C62904 _0561_/a_149_47# VGND 0.12909f 
C62905 _0561_/a_245_297# VGND 0 
C62906 _0561_/a_51_297# VGND 0.29706f 
C62907 clknet_1_1__leaf__0465_ VGND 6.06567f
C62908 clknet_1_1__leaf__0464_ VGND 3.90686f
C62909 _0394_ VGND 0.36375f
C62910 _0306_ VGND 0.56658f
C62911 _0308_ VGND 0.99262f
C62912 _0776_/a_27_47# VGND 0.19572f 
C62913 _0776_/a_109_297# VGND 0 
C62914 _0449_ VGND 0.23176f
C62915 _0845_/a_109_47# VGND 0.24277f 
C62916 _0845_/a_193_297# VGND 0 
C62917 _0845_/a_109_297# VGND 0 
C62918 net147 VGND 0.42092f
C62919 _1061_/a_1017_47# VGND 0.00447f 
C62920 _1061_/a_592_47# VGND 0.00769f 
C62921 _1061_/a_975_413# VGND 0 
C62922 _1061_/a_561_413# VGND 0 
C62923 _1061_/a_381_47# VGND 0.06889f 
C62924 _1061_/a_891_413# VGND 0.3046f 
C62925 _1061_/a_1059_315# VGND 0.53293f 
C62926 _1061_/a_466_413# VGND 0.22505f 
C62927 _1061_/a_634_159# VGND 0.27006f 
C62928 _1061_/a_193_47# VGND 0.46803f 
C62929 _1061_/a_27_47# VGND 0.58351f 
C62930 net98 VGND 0.39019f
C62931 clknet_1_1__leaf__0461_ VGND 4.83892f
C62932 clkbuf_0__0459_/a_110_47# VGND 2.25914f 
C62933 _0095_ VGND 0.39315f
C62934 _0407_ VGND 0.17891f
C62935 _0793_/a_240_47# VGND 0.16104f 
C62936 _0793_/a_149_47# VGND 0.125f 
C62937 _0793_/a_51_297# VGND 0.28856f 
C62938 net107 VGND 0.33574f
C62939 clknet_1_0__leaf__0461_ VGND 4.06178f
C62940 clknet_1_1__leaf__0457_ VGND 2.38951f
C62941 clkbuf_1_1__f__0457_/a_110_47# VGND 2.17124f 
C62942 _0148_ VGND 0.31957f
C62943 net170 VGND 1.77305f
C62944 _0196_ VGND 0.27424f
C62945 _0528_/a_384_47# VGND 0.00339f 
C62946 _0528_/a_299_297# VGND 0.04292f 
C62947 _0528_/a_81_21# VGND 0.31329f 
C62948 acc0.A\[28\] VGND 1.22141f
C62949 net114 VGND 0.8497f
C62950 _1028_/a_1017_47# VGND 0.00447f 
C62951 _1028_/a_592_47# VGND 0.00748f 
C62952 _1028_/a_381_47# VGND 0.06538f 
C62953 _1028_/a_891_413# VGND 0.3041f 
C62954 _1028_/a_1059_315# VGND 0.4147f 
C62955 _1028_/a_466_413# VGND 0.23829f 
C62956 _1028_/a_634_159# VGND 0.28273f 
C62957 _1028_/a_193_47# VGND 0.3669f 
C62958 _1028_/a_27_47# VGND 0.58277f 
C62959 _0545_/a_150_297# VGND 0 
C62960 _0545_/a_68_297# VGND 0.26519f 
C62961 _0246_ VGND 1.28181f
C62962 _0245_ VGND 0.64579f
C62963 _0614_/a_29_53# VGND 0.41764f 
C62964 _0829_/a_27_47# VGND 0.17888f 
C62965 _0829_/a_109_297# VGND 0 
C62966 net184 VGND 0.39094f
C62967 net131 VGND 0.35063f
C62968 _1045_/a_1017_47# VGND 0.00408f 
C62969 _1045_/a_592_47# VGND 0.00788f 
C62970 _1045_/a_975_413# VGND 0 
C62971 _1045_/a_561_413# VGND 0 
C62972 _1045_/a_381_47# VGND 0.06928f 
C62973 _1045_/a_891_413# VGND 0.29961f 
C62974 _1045_/a_1059_315# VGND 0.43574f 
C62975 _1045_/a_466_413# VGND 0.22564f 
C62976 _1045_/a_634_159# VGND 0.27245f 
C62977 _1045_/a_193_47# VGND 0.46988f 
C62978 _1045_/a_27_47# VGND 0.57659f 
C62979 _0171_ VGND 1.46663f
C62980 _0493_/a_27_47# VGND 0.3399f 
C62981 _0562_/a_150_297# VGND 0 
C62982 _0562_/a_68_297# VGND 0.28177f 
C62983 _0263_ VGND 1.60498f
C62984 _0261_ VGND 0.96187f
C62985 _0262_ VGND 0.40807f
C62986 _0631_/a_109_297# VGND 0.00122f 
C62987 _0332_ VGND 0.41235f
C62988 _0700_/a_113_47# VGND 0.002f 
C62989 hold9/a_391_47# VGND 0.24555f 
C62990 hold9/a_285_47# VGND 0.40359f 
C62991 hold9/a_49_47# VGND 0.44617f 
C62992 _0395_ VGND 0.9376f
C62993 _0777_/a_285_47# VGND 0.23615f 
C62994 _0777_/a_129_47# VGND 0.00456f 
C62995 _0777_/a_377_297# VGND 0.00181f 
C62996 _0777_/a_47_47# VGND 0.34414f 
C62997 _0846_/a_240_47# VGND 0.16256f 
C62998 _0846_/a_149_47# VGND 0.12645f 
C62999 _0846_/a_512_297# VGND 0 
C63000 _0846_/a_245_297# VGND 0 
C63001 _0846_/a_51_297# VGND 0.29645f 
C63002 _0160_ VGND 0.48199f
C63003 _1062_/a_1017_47# VGND 0.0046f 
C63004 _1062_/a_592_47# VGND 0.00788f 
C63005 _1062_/a_975_413# VGND 0 
C63006 _1062_/a_561_413# VGND 0 
C63007 _1062_/a_381_47# VGND 0.06803f 
C63008 _1062_/a_891_413# VGND 0.28624f 
C63009 _1062_/a_1059_315# VGND 0.39432f 
C63010 _1062_/a_466_413# VGND 0.22217f 
C63011 _1062_/a_634_159# VGND 0.27077f 
C63012 _1062_/a_193_47# VGND 0.41364f 
C63013 _1062_/a_27_47# VGND 0.61387f 
C63014 _0277_ VGND 0.86094f
C63015 _0300_ VGND 0.59297f
C63016 _0297_ VGND 2.07613f
C63017 _0794_/a_326_47# VGND 0.00481f 
C63018 _0794_/a_27_47# VGND 0.23915f 
C63019 _0794_/a_110_297# VGND 0 
C63020 clkbuf_1_1__f__0458_/a_110_47# VGND 2.25396f 
C63021 _0460_ VGND 1.76205f
C63022 clknet_1_0__leaf__0457_ VGND 3.98944f
C63023 _0880_/a_27_47# VGND 0.31527f 
C63024 net10 VGND 1.52427f
C63025 _0529_/a_373_47# VGND 0.00468f 
C63026 _0529_/a_109_47# VGND 0.00842f 
C63027 _0529_/a_109_297# VGND 0.01525f 
C63028 _0529_/a_27_297# VGND 0.4778f 
C63029 net191 VGND 0.31274f
C63030 net115 VGND 0.63571f
C63031 _1029_/a_1017_47# VGND 0.00526f 
C63032 _1029_/a_592_47# VGND 0.01049f 
C63033 _1029_/a_975_413# VGND 0 
C63034 _1029_/a_561_413# VGND 0 
C63035 _1029_/a_381_47# VGND 0.07142f 
C63036 _1029_/a_891_413# VGND 0.32401f 
C63037 _1029_/a_1059_315# VGND 0.45031f 
C63038 _1029_/a_466_413# VGND 0.24689f 
C63039 _1029_/a_634_159# VGND 0.30818f 
C63040 _1029_/a_193_47# VGND 0.50915f 
C63041 _1029_/a_27_47# VGND 0.64769f 
C63042 _0615_/a_109_297# VGND 0 
C63043 _0139_ VGND 0.47574f
C63044 net32 VGND 0.30746f
C63045 net152 VGND 0.8292f
C63046 _0205_ VGND 0.2634f
C63047 _0546_/a_240_47# VGND 0.17083f 
C63048 _0546_/a_149_47# VGND 0.12614f 
C63049 _0546_/a_512_297# VGND 0 
C63050 _0546_/a_245_297# VGND 0 
C63051 _0546_/a_51_297# VGND 0.28302f 
C63052 net132 VGND 0.5401f
C63053 _1046_/a_1017_47# VGND 0.00474f 
C63054 _1046_/a_592_47# VGND 0.008f 
C63055 _1046_/a_975_413# VGND 0 
C63056 _1046_/a_561_413# VGND 0 
C63057 _1046_/a_381_47# VGND 0.06776f 
C63058 _1046_/a_891_413# VGND 0.29844f 
C63059 _1046_/a_1059_315# VGND 0.42252f 
C63060 _1046_/a_466_413# VGND 0.22178f 
C63061 _1046_/a_634_159# VGND 0.26462f 
C63062 _1046_/a_193_47# VGND 0.39479f 
C63063 _1046_/a_27_47# VGND 0.61316f 
C63064 _0494_/a_27_47# VGND 0.44977f 
C63065 _0264_ VGND 0.84874f
C63066 _0632_/a_113_47# VGND 0.002f 
C63067 _0214_ VGND 0.37942f
C63068 _0563_/a_240_47# VGND 0.16239f 
C63069 _0563_/a_149_47# VGND 0.12619f 
C63070 _0563_/a_512_297# VGND 0 
C63071 _0563_/a_245_297# VGND 0 
C63072 _0563_/a_51_297# VGND 0.29169f 
C63073 _0333_ VGND 1.7197f
C63074 _0701_/a_303_47# VGND 0.00505f 
C63075 _0701_/a_209_47# VGND 0.00544f 
C63076 _0701_/a_209_297# VGND 0.00669f 
C63077 _0701_/a_80_21# VGND 0.40144f 
C63078 hold8/a_391_47# VGND 0.25406f 
C63079 hold8/a_285_47# VGND 0.40945f 
C63080 hold8/a_49_47# VGND 0.4853f 
C63081 _0847_/a_109_297# VGND 0 
C63082 _0778_/a_150_297# VGND 0 
C63083 _0778_/a_68_297# VGND 0.28189f 
C63084 _0161_ VGND 0.90461f
C63085 _1063_/a_1017_47# VGND 0.00404f 
C63086 _1063_/a_592_47# VGND 0.00674f 
C63087 _1063_/a_561_413# VGND 0 
C63088 _1063_/a_381_47# VGND 0.06129f 
C63089 _1063_/a_891_413# VGND 0.27452f 
C63090 _1063_/a_1059_315# VGND 0.38454f 
C63091 _1063_/a_466_413# VGND 0.21343f 
C63092 _1063_/a_634_159# VGND 0.25207f 
C63093 _1063_/a_193_47# VGND 0.34703f 
C63094 _1063_/a_27_47# VGND 0.57365f 
C63095 _0117_ VGND 0.19672f
C63096 _0580_/a_373_47# VGND 0.00216f 
C63097 _0580_/a_109_47# VGND 0.00631f 
C63098 _0580_/a_109_297# VGND 0.00376f 
C63099 _0580_/a_27_297# VGND 0.4325f 
C63100 _0409_ VGND 0.49806f
C63101 _0795_/a_384_47# VGND 0.00329f 
C63102 _0795_/a_299_297# VGND 0.04199f 
C63103 _0795_/a_81_21# VGND 0.32142f 
C63104 B[11] VGND 0.60737f
C63105 input19/a_75_212# VGND 0.33005f 
C63106 clkbuf_1_1__f__0459_/a_110_47# VGND 2.34765f 
C63107 _0950_/a_75_212# VGND 0.32264f 
C63108 net116 VGND 0.30712f
C63109 _0206_ VGND 0.33721f
C63110 comp0.B\[8\] VGND 0.95878f
C63111 _0547_/a_150_297# VGND 0 
C63112 _0547_/a_68_297# VGND 0.26864f 
C63113 _0240_ VGND 0.85565f
C63114 _0247_ VGND 0.61825f
C63115 _0616_/a_215_47# VGND 0.28928f 
C63116 _0616_/a_78_199# VGND 0.21039f 
C63117 _0145_ VGND 0.24675f
C63118 _1047_/a_1017_47# VGND 0.00447f 
C63119 _1047_/a_592_47# VGND 0.00662f 
C63120 _1047_/a_381_47# VGND 0.06058f 
C63121 _1047_/a_891_413# VGND 0.28426f 
C63122 _1047_/a_1059_315# VGND 0.3947f 
C63123 _1047_/a_466_413# VGND 0.21148f 
C63124 _1047_/a_634_159# VGND 0.2513f 
C63125 _1047_/a_193_47# VGND 0.34453f 
C63126 _1047_/a_27_47# VGND 0.55386f 
C63127 _0215_ VGND 0.42002f
C63128 _0175_ VGND 2.58668f
C63129 _0564_/a_150_297# VGND 0 
C63130 _0564_/a_68_297# VGND 0.26774f 
C63131 _0495_/a_150_297# VGND 0 
C63132 _0495_/a_68_297# VGND 0.26543f 
C63133 _0265_ VGND 0.31928f
C63134 net47 VGND 2.15306f
C63135 _0633_/a_109_297# VGND 0 
C63136 _0334_ VGND 0.61275f
C63137 _0702_/a_113_47# VGND 0.0017f 
C63138 hold7/a_391_47# VGND 0.24431f 
C63139 hold7/a_285_47# VGND 0.41065f 
C63140 hold7/a_49_47# VGND 0.44381f 
C63141 _0097_ VGND 0.3502f
C63142 _0396_ VGND 0.23971f
C63143 _0779_/a_510_47# VGND 0.00857f 
C63144 _0779_/a_215_47# VGND 0.23357f 
C63145 _0779_/a_297_297# VGND 0 
C63146 _0779_/a_79_21# VGND 0.34591f 
C63147 _0451_ VGND 0.59015f
C63148 _0450_ VGND 0.43021f
C63149 _0446_ VGND 0.8886f
C63150 _0848_/a_27_47# VGND 0.1714f 
C63151 _1064_/a_1017_47# VGND 0.00467f 
C63152 _1064_/a_592_47# VGND 0.00777f 
C63153 _1064_/a_975_413# VGND 0 
C63154 _1064_/a_561_413# VGND 0 
C63155 _1064_/a_381_47# VGND 0.07116f 
C63156 _1064_/a_891_413# VGND 0.29902f 
C63157 _1064_/a_1059_315# VGND 0.42011f 
C63158 _1064_/a_466_413# VGND 0.24343f 
C63159 _1064_/a_634_159# VGND 0.28517f 
C63160 _1064_/a_193_47# VGND 0.51196f 
C63161 _1064_/a_27_47# VGND 0.66677f 
C63162 acc0.A\[10\] VGND 2.13721f
C63163 _0650_/a_150_297# VGND 0 
C63164 _0650_/a_68_297# VGND 0.27285f 
C63165 _0116_ VGND 0.29174f
C63166 net206 VGND 1.24165f
C63167 net219 VGND 0.47945f
C63168 _0581_/a_373_47# VGND 0.00216f 
C63169 _0581_/a_109_47# VGND 0.00628f 
C63170 _0581_/a_109_297# VGND 0.00366f 
C63171 _0581_/a_27_297# VGND 0.42589f 
C63172 _0094_ VGND 0.34707f
C63173 _0410_ VGND 0.56048f
C63174 net238 VGND 0.24162f
C63175 _0796_/a_510_47# VGND 0.00782f 
C63176 _0796_/a_215_47# VGND 0.2273f 
C63177 _0796_/a_297_297# VGND 0 
C63178 _0796_/a_79_21# VGND 0.35899f 
C63179 net29 VGND 0.32681f
C63180 B[6] VGND 0.70187f
C63181 input29/a_75_212# VGND 0.35506f 
C63182 B[10] VGND 0.72025f
C63183 input18/a_75_212# VGND 0.36913f 
C63184 comp0.B\[0\] VGND 1.96446f
C63185 _0951_/a_368_53# VGND 0.00258f 
C63186 _0951_/a_296_53# VGND 0 
C63187 _0951_/a_209_311# VGND 0.27444f 
C63188 _0951_/a_109_93# VGND 0.22446f 
C63189 _0617_/a_150_297# VGND 0 
C63190 _0617_/a_68_297# VGND 0.27666f 
C63191 _0138_ VGND 0.39867f
C63192 net173 VGND 0.54686f
C63193 _0548_/a_240_47# VGND 0.16199f 
C63194 _0548_/a_149_47# VGND 0.12675f 
C63195 _0548_/a_245_297# VGND 0 
C63196 _0548_/a_51_297# VGND 0.2918f 
C63197 clkbuf_1_1__f_clk/a_110_47# VGND 2.22889f 
C63198 net134 VGND 0.85051f
C63199 _1048_/a_1017_47# VGND 0.00489f 
C63200 _1048_/a_592_47# VGND 0.00813f 
C63201 _1048_/a_975_413# VGND 0 
C63202 _1048_/a_561_413# VGND 0 
C63203 _1048_/a_381_47# VGND 0.07063f 
C63204 _1048_/a_891_413# VGND 0.29851f 
C63205 _1048_/a_1059_315# VGND 0.41296f 
C63206 _1048_/a_466_413# VGND 0.22503f 
C63207 _1048_/a_634_159# VGND 0.27194f 
C63208 _1048_/a_193_47# VGND 0.39357f 
C63209 _1048_/a_27_47# VGND 0.6346f 
C63210 _0634_/a_113_47# VGND 0.00168f 
C63211 net201 VGND 0.89756f
C63212 _0565_/a_240_47# VGND 0.17795f 
C63213 _0565_/a_149_47# VGND 0.1316f 
C63214 _0565_/a_512_297# VGND 0.00106f 
C63215 _0565_/a_245_297# VGND 0.0012f 
C63216 _0565_/a_51_297# VGND 0.31663f 
C63217 _0176_ VGND 6.05461f
C63218 _0496_/a_27_47# VGND 0.42031f 
C63219 _0703_/a_109_297# VGND 0 
C63220 hold6/a_391_47# VGND 0.26048f 
C63221 hold6/a_285_47# VGND 0.42135f 
C63222 hold6/a_49_47# VGND 0.45414f 
C63223 _0082_ VGND 0.55298f
C63224 net222 VGND 0.21175f
C63225 _0849_/a_510_47# VGND 0.00782f 
C63226 _0849_/a_215_47# VGND 0.23165f 
C63227 _0849_/a_297_297# VGND 0 
C63228 _0849_/a_79_21# VGND 0.3597f 
C63229 control0.reset VGND 1.22221f
C63230 _1065_/a_1017_47# VGND 0.00414f 
C63231 _1065_/a_592_47# VGND 0.00684f 
C63232 _1065_/a_975_413# VGND 0 
C63233 _1065_/a_561_413# VGND 0 
C63234 _1065_/a_381_47# VGND 0.06193f 
C63235 _1065_/a_891_413# VGND 0.27689f 
C63236 _1065_/a_1059_315# VGND 0.38856f 
C63237 _1065_/a_466_413# VGND 0.21395f 
C63238 _1065_/a_634_159# VGND 0.25351f 
C63239 _1065_/a_193_47# VGND 0.34816f 
C63240 _1065_/a_27_47# VGND 0.59322f 
C63241 net83 VGND 0.64853f
C63242 _0115_ VGND 1.00122f
C63243 net221 VGND 0.29836f
C63244 _0582_/a_373_47# VGND 0.00344f 
C63245 _0582_/a_109_47# VGND 0.0076f 
C63246 _0582_/a_109_297# VGND 0.00468f 
C63247 _0582_/a_27_297# VGND 0.45958f 
C63248 _0282_ VGND 0.34973f
C63249 _0651_/a_113_47# VGND 0.00164f 
C63250 net239 VGND 0.55827f
C63251 _0720_/a_150_297# VGND 0 
C63252 _0720_/a_68_297# VGND 0.28601f 
C63253 _0797_/a_297_47# VGND 0.00517f 
C63254 _0797_/a_207_413# VGND 0.25803f 
C63255 _0797_/a_27_413# VGND 0.29145f 
C63256 _0465_ VGND 2.33599f
C63257 _0935_/a_27_47# VGND 0.3102f 
C63258 clknet_0__0460_ VGND 3.3065f
C63259 clkbuf_1_0__f__0460_/a_110_47# VGND 2.27242f 
C63260 net28 VGND 0.28213f
C63261 B[5] VGND 0.57787f
C63262 input28/a_75_212# VGND 0.36298f 
C63263 net17 VGND 3.92106f
C63264 B[0] VGND 0.76187f
C63265 input17/a_75_212# VGND 0.36723f 
C63266 net102 VGND 0.29545f
C63267 _0471_ VGND 0.47902f
C63268 _0207_ VGND 0.35056f
C63269 net171 VGND 0.90108f
C63270 _0549_/a_150_297# VGND 0 
C63271 _0549_/a_68_297# VGND 0.26135f 
C63272 _0250_ VGND 1.20079f
C63273 _0249_ VGND 0.47035f
C63274 _0618_/a_510_47# VGND 0.00607f 
C63275 _0618_/a_215_47# VGND 0.21784f 
C63276 _0618_/a_297_297# VGND 0 
C63277 _0618_/a_79_21# VGND 0.33492f 
C63278 acc0.A\[3\] VGND 0.87279f
C63279 _0147_ VGND 0.69157f
C63280 net135 VGND 0.44123f
C63281 _1049_/a_1017_47# VGND 0.00461f 
C63282 _1049_/a_592_47# VGND 0.00785f 
C63283 _1049_/a_975_413# VGND 0 
C63284 _1049_/a_561_413# VGND 0 
C63285 _1049_/a_381_47# VGND 0.06082f 
C63286 _1049_/a_891_413# VGND 0.28608f 
C63287 _1049_/a_1059_315# VGND 0.39723f 
C63288 _1049_/a_466_413# VGND 0.22098f 
C63289 _1049_/a_634_159# VGND 0.26311f 
C63290 _1049_/a_193_47# VGND 0.3529f 
C63291 _1049_/a_27_47# VGND 0.59324f 
C63292 _0177_ VGND 0.31933f
C63293 _0497_/a_150_297# VGND 0 
C63294 _0497_/a_68_297# VGND 0.25974f 
C63295 acc0.A\[30\] VGND 1.17969f
C63296 _0704_/a_150_297# VGND 0.00127f 
C63297 _0704_/a_68_297# VGND 0.2941f 
C63298 _0267_ VGND 1.1419f
C63299 _0635_/a_27_47# VGND 0.17593f 
C63300 _0635_/a_109_297# VGND 0 
C63301 _0566_/a_27_47# VGND 0.69422f 
C63302 hold5/a_391_47# VGND 0.25833f 
C63303 hold5/a_285_47# VGND 0.41656f 
C63304 hold5/a_49_47# VGND 0.46166f 
C63305 control0.sh VGND 2.77958f
C63306 clknet_1_1__leaf_clk VGND 2.48371f
C63307 _1066_/a_1017_47# VGND 0.00404f 
C63308 _1066_/a_592_47# VGND 0.00662f 
C63309 _1066_/a_381_47# VGND 0.06058f 
C63310 _1066_/a_891_413# VGND 0.29466f 
C63311 _1066_/a_1059_315# VGND 0.42073f 
C63312 _1066_/a_466_413# VGND 0.21622f 
C63313 _1066_/a_634_159# VGND 0.25325f 
C63314 _1066_/a_193_47# VGND 0.36303f 
C63315 _1066_/a_27_47# VGND 0.57532f 
C63316 _0114_ VGND 0.20841f
C63317 net165 VGND 0.54506f
C63318 _0583_/a_373_47# VGND 0.00288f 
C63319 _0583_/a_109_47# VGND 0.0076f 
C63320 _0583_/a_109_297# VGND 0.00279f 
C63321 _0583_/a_27_297# VGND 0.43925f 
C63322 _0721_/a_27_47# VGND 0.69704f 
C63323 _0798_/a_199_47# VGND 0.00406f 
C63324 _0798_/a_113_297# VGND 0.04057f 
C63325 clknet_0__0461_ VGND 2.76465f
C63326 clkbuf_1_0__f__0461_/a_110_47# VGND 2.19452f 
C63327 net27 VGND 0.40933f
C63328 B[4] VGND 0.77292f
C63329 input27/a_75_212# VGND 0.31265f 
C63330 A[9] VGND 0.65135f
C63331 input16/a_75_212# VGND 0.33594f 
C63332 comp0.B\[10\] VGND 0.77676f
C63333 _0953_/a_304_297# VGND 0.00172f 
C63334 _0953_/a_220_297# VGND 0.00236f 
C63335 _0953_/a_114_297# VGND 0.00538f 
C63336 _0953_/a_32_297# VGND 0.78418f 
C63337 _0162_ VGND 0.82216f
C63338 _0487_ VGND 2.46634f
C63339 _0485_ VGND 0.66138f
C63340 _0484_ VGND 1.13847f
C63341 _0970_/a_285_47# VGND 0.00375f 
C63342 _0970_/a_114_47# VGND 0.01078f 
C63343 _0970_/a_27_297# VGND 0.06485f 
C63344 _0619_/a_150_297# VGND 0 
C63345 _0619_/a_68_297# VGND 0.27316f 
C63346 net143 VGND 0.40951f
C63347 _0567_/a_373_47# VGND 0.00339f 
C63348 _0567_/a_109_47# VGND 0.00698f 
C63349 _0567_/a_109_297# VGND 0.01623f 
C63350 _0567_/a_27_297# VGND 0.45533f 
C63351 _0159_ VGND 0.60928f
C63352 net7 VGND 0.33528f
C63353 net247 VGND 0.38228f
C63354 _0498_/a_240_47# VGND 0.17221f 
C63355 _0498_/a_149_47# VGND 0.13206f 
C63356 _0498_/a_512_297# VGND 0 
C63357 _0498_/a_245_297# VGND 0 
C63358 _0498_/a_51_297# VGND 0.28548f 
C63359 _0336_ VGND 0.85582f
C63360 _0220_ VGND 1.91038f
C63361 _0705_/a_145_75# VGND 0.00491f 
C63362 _0705_/a_59_75# VGND 0.2873f 
C63363 _0636_/a_145_75# VGND 0.00528f 
C63364 _0636_/a_59_75# VGND 0.32737f 
C63365 hold4/a_391_47# VGND 0.27999f 
C63366 hold4/a_285_47# VGND 0.43211f 
C63367 hold4/a_49_47# VGND 0.44326f 
C63368 control0.add VGND 1.28068f
C63369 _1067_/a_1017_47# VGND 0.00404f 
C63370 _1067_/a_592_47# VGND 0.00662f 
C63371 _1067_/a_381_47# VGND 0.06058f 
C63372 _1067_/a_891_413# VGND 0.27785f 
C63373 _1067_/a_1059_315# VGND 0.3948f 
C63374 _1067_/a_466_413# VGND 0.21294f 
C63375 _1067_/a_634_159# VGND 0.25176f 
C63376 _1067_/a_193_47# VGND 0.34279f 
C63377 _1067_/a_27_47# VGND 0.58378f 
C63378 net157 VGND 1.87159f
C63379 _0584_/a_373_47# VGND 0.00302f 
C63380 _0584_/a_109_47# VGND 0.00767f 
C63381 _0584_/a_109_297# VGND 0.00371f 
C63382 _0584_/a_27_297# VGND 0.43939f 
C63383 _0110_ VGND 0.54374f
C63384 _0351_ VGND 0.36295f
C63385 _0722_/a_510_47# VGND 0.0078f 
C63386 _0722_/a_215_47# VGND 0.23702f 
C63387 _0722_/a_297_297# VGND 0 
C63388 _0722_/a_79_21# VGND 0.3684f 
C63389 acc0.A\[11\] VGND 2.32132f
C63390 net38 VGND 1.85176f
C63391 _0653_/a_113_47# VGND 0.002f 
C63392 _0411_ VGND 0.37406f
C63393 _0799_/a_303_47# VGND 0.00692f 
C63394 _0799_/a_209_47# VGND 0.01091f 
C63395 _0799_/a_209_297# VGND 0.01608f 
C63396 _0799_/a_80_21# VGND 0.43801f 
C63397 _0302_ VGND 0.49689f
C63398 _0670_/a_510_47# VGND 0.00785f 
C63399 _0670_/a_215_47# VGND 0.23174f 
C63400 _0670_/a_297_297# VGND 0 
C63401 _0670_/a_79_21# VGND 0.38513f 
C63402 clknet_0__0462_ VGND 2.32372f
C63403 clkbuf_1_0__f__0462_/a_110_47# VGND 2.26058f 
C63404 net26 VGND 1.01428f
C63405 B[3] VGND 0.7204f
C63406 input26/a_75_212# VGND 0.38037f 
C63407 A[8] VGND 0.63589f
C63408 input15/a_75_212# VGND 0.30916f 
C63409 comp0.B\[12\] VGND 1.20908f
C63410 comp0.B\[11\] VGND 1.6952f
C63411 _0954_/a_304_297# VGND 0 
C63412 _0954_/a_114_297# VGND 0.00172f 
C63413 _0954_/a_32_297# VGND 0.75758f 
C63414 _0163_ VGND 0.40716f
C63415 _0181_ VGND 6.82649f
C63416 _0971_/a_384_47# VGND 0.00334f 
C63417 _0971_/a_299_297# VGND 0.03862f 
C63418 _0971_/a_81_21# VGND 0.31199f 
C63419 _0178_ VGND 1.186f
C63420 _0499_/a_145_75# VGND 0.00468f 
C63421 _0499_/a_59_75# VGND 0.29039f 
C63422 _0128_ VGND 0.41645f
C63423 net208 VGND 0.27491f
C63424 _0568_/a_373_47# VGND 0.00329f 
C63425 _0568_/a_109_47# VGND 0.00737f 
C63426 _0568_/a_109_297# VGND 0.00396f 
C63427 _0568_/a_27_297# VGND 0.45498f 
C63428 _0269_ VGND 0.84308f
C63429 _0268_ VGND 1.44716f
C63430 _0637_/a_139_47# VGND 0.00381f 
C63431 _0637_/a_311_297# VGND 0 
C63432 _0637_/a_56_297# VGND 0.03665f 
C63433 hold3/a_391_47# VGND 0.23934f 
C63434 hold3/a_285_47# VGND 0.40275f 
C63435 hold3/a_49_47# VGND 0.4598f 
C63436 _0166_ VGND 0.26695f
C63437 _1068_/a_1017_47# VGND 0.00418f 
C63438 _1068_/a_592_47# VGND 0.00728f 
C63439 _1068_/a_975_413# VGND 0 
C63440 _1068_/a_561_413# VGND 0 
C63441 _1068_/a_381_47# VGND 0.06343f 
C63442 _1068_/a_891_413# VGND 0.28013f 
C63443 _1068_/a_1059_315# VGND 0.40871f 
C63444 _1068_/a_466_413# VGND 0.21637f 
C63445 _1068_/a_634_159# VGND 0.2586f 
C63446 _1068_/a_193_47# VGND 0.35461f 
C63447 _1068_/a_27_47# VGND 0.5672f 
C63448 _0112_ VGND 0.47795f
C63449 net149 VGND 2.32726f
C63450 _0585_/a_373_47# VGND 0.00344f 
C63451 _0585_/a_109_47# VGND 0.00753f 
C63452 _0585_/a_109_297# VGND 0.00309f 
C63453 _0585_/a_27_297# VGND 0.43819f 
C63454 _0654_/a_297_47# VGND 0.00504f 
C63455 _0654_/a_207_413# VGND 0.24989f 
C63456 _0654_/a_27_413# VGND 0.28469f 
C63457 _0723_/a_297_47# VGND 0.00516f 
C63458 _0723_/a_207_413# VGND 0.25062f 
C63459 _0723_/a_27_413# VGND 0.28606f 
C63460 clknet_1_0__leaf__0460_ VGND 5.17634f
C63461 _0459_ VGND 2.5979f
C63462 _0869_/a_27_47# VGND 0.31749f 
C63463 _0303_ VGND 0.32902f
C63464 _0671_/a_199_47# VGND 0.00395f 
C63465 _0671_/a_113_297# VGND 0.03968f 
C63466 clkbuf_1_0__f__0463_/a_110_47# VGND 2.25134f 
C63467 net25 VGND 0.30662f
C63468 B[2] VGND 0.55323f
C63469 input25/a_75_212# VGND 0.33063f 
C63470 A[7] VGND 0.52737f
C63471 input14/a_75_212# VGND 0.34512f 
C63472 _0324_ VGND 0.92486f
C63473 _0359_ VGND 1.06311f
C63474 _0740_/a_113_47# VGND 0.00207f 
C63475 _0474_ VGND 0.76287f
C63476 comp0.B\[6\] VGND 1.27968f
C63477 comp0.B\[5\] VGND 0.68752f
C63478 comp0.B\[3\] VGND 0.54535f
C63479 _0955_/a_304_297# VGND 0 
C63480 _0955_/a_220_297# VGND 0 
C63481 _0955_/a_114_297# VGND 0 
C63482 _0955_/a_32_297# VGND 0.77185f 
C63483 _0164_ VGND 0.23852f
C63484 net231 VGND 0.43507f
C63485 _0972_/a_584_47# VGND 0.00536f 
C63486 _0972_/a_346_47# VGND 0.0034f 
C63487 _0972_/a_256_47# VGND 0.00243f 
C63488 _0972_/a_250_297# VGND 0.03198f 
C63489 _0972_/a_93_21# VGND 0.38307f 
C63490 net62 VGND 3.07912f
C63491 _0638_/a_109_297# VGND 0 
C63492 _0127_ VGND 0.44351f
C63493 acc0.A\[29\] VGND 2.46452f
C63494 _0569_/a_373_47# VGND 0.00344f 
C63495 _0569_/a_109_47# VGND 0.00797f 
C63496 _0569_/a_109_297# VGND 0.00401f 
C63497 _0569_/a_27_297# VGND 0.44589f 
C63498 _0339_ VGND 1.29148f
C63499 _0338_ VGND 0.8388f
C63500 _0335_ VGND 0.98812f
C63501 _0707_/a_315_47# VGND 0.00119f 
C63502 _0707_/a_208_47# VGND 0.00287f 
C63503 _0707_/a_544_297# VGND 0 
C63504 _0707_/a_201_297# VGND 0.00506f 
C63505 _0707_/a_75_199# VGND 0.54908f 
C63506 hold2/a_391_47# VGND 0.26787f 
C63507 hold2/a_285_47# VGND 0.46255f 
C63508 hold2/a_49_47# VGND 0.47602f 
C63509 control0.count\[0\] VGND 0.95977f
C63510 _0167_ VGND 0.34744f
C63511 clknet_1_0__leaf_clk VGND 4.58201f
C63512 _1069_/a_1017_47# VGND 0.00447f 
C63513 _1069_/a_592_47# VGND 0.00748f 
C63514 _1069_/a_381_47# VGND 0.06759f 
C63515 _1069_/a_891_413# VGND 0.28365f 
C63516 _1069_/a_1059_315# VGND 0.39312f 
C63517 _1069_/a_466_413# VGND 0.22445f 
C63518 _1069_/a_634_159# VGND 0.26887f 
C63519 _1069_/a_193_47# VGND 0.45636f 
C63520 _1069_/a_27_47# VGND 0.61528f 
C63521 _0724_/a_199_47# VGND 0.00397f 
C63522 _0724_/a_113_297# VGND 0.03849f 
C63523 _0218_ VGND 9.75844f
C63524 _0586_/a_27_47# VGND 0.40444f 
C63525 _0286_ VGND 1.05361f
C63526 _0283_ VGND 0.97971f
C63527 _0655_/a_369_297# VGND 0 
C63528 _0655_/a_109_93# VGND 0.24874f 
C63529 _0655_/a_215_53# VGND 0.36898f 
C63530 _0296_ VGND 0.63402f
C63531 _0672_/a_510_47# VGND 0.00892f 
C63532 _0672_/a_215_47# VGND 0.23792f 
C63533 _0672_/a_297_297# VGND 0 
C63534 _0672_/a_79_21# VGND 0.38639f 
C63535 _0367_ VGND 0.27291f
C63536 _0315_ VGND 1.64946f
C63537 _0366_ VGND 1.13427f
C63538 _0741_/a_109_297# VGND 0 
C63539 clkbuf_1_0__f__0464_/a_110_47# VGND 2.22128f 
C63540 net24 VGND 0.29373f
C63541 B[1] VGND 0.90129f
C63542 input24/a_75_212# VGND 0.31695f 
C63543 A[6] VGND 0.72386f
C63544 input13/a_75_212# VGND 0.35f 
C63545 _0421_ VGND 0.30167f
C63546 _0810_/a_113_47# VGND 0.00187f 
C63547 comp0.B\[15\] VGND 1.06799f
C63548 _0956_/a_304_297# VGND 0 
C63549 _0956_/a_220_297# VGND 0 
C63550 _0956_/a_114_297# VGND 0 
C63551 _0956_/a_32_297# VGND 0.80286f 
C63552 _0165_ VGND 0.34746f
C63553 net240 VGND 0.24205f
C63554 _0973_/a_373_47# VGND 0.00288f 
C63555 _0973_/a_109_47# VGND 0.00795f 
C63556 _0973_/a_109_297# VGND 0.00274f 
C63557 _0973_/a_27_297# VGND 0.4554f 
C63558 net118 VGND 0.42862f
C63559 _0088_ VGND 0.49693f
C63560 _0990_/a_1017_47# VGND 0.00404f 
C63561 _0990_/a_592_47# VGND 0.00748f 
C63562 _0990_/a_381_47# VGND 0.06538f 
C63563 _0990_/a_891_413# VGND 0.27546f 
C63564 _0990_/a_1059_315# VGND 0.38594f 
C63565 _0990_/a_466_413# VGND 0.21702f 
C63566 _0990_/a_634_159# VGND 0.25246f 
C63567 _0990_/a_193_47# VGND 0.36721f 
C63568 _0990_/a_27_47# VGND 0.59468f 
C63569 _0271_ VGND 1.03267f
C63570 _0256_ VGND 0.74903f
C63571 _0270_ VGND 0.59571f
C63572 _0639_/a_109_297# VGND 0 
C63573 net60 VGND 0.98547f
C63574 _0708_/a_150_297# VGND 0 
C63575 _0708_/a_68_297# VGND 0.28051f 
C63576 hold1/a_391_47# VGND 0.25927f 
C63577 hold1/a_285_47# VGND 0.41776f 
C63578 hold1/a_49_47# VGND 0.46256f 
C63579 _0187_ VGND 1.20017f
C63580 net4 VGND 0.4303f
C63581 _0510_/a_373_47# VGND 0.00234f 
C63582 _0510_/a_109_47# VGND 0.00638f 
C63583 _0510_/a_109_297# VGND 0.0051f 
C63584 _0510_/a_27_297# VGND 0.43454f 
C63585 _0587_/a_27_47# VGND 0.68116f 
C63586 _0288_ VGND 0.73415f
C63587 acc0.A\[9\] VGND 1.60083f
C63588 _0656_/a_145_75# VGND 0.00544f 
C63589 _0656_/a_59_75# VGND 0.32412f 
C63590 _0353_ VGND 0.83667f
C63591 _0725_/a_303_47# VGND 0.00665f 
C63592 _0725_/a_209_47# VGND 0.00729f 
C63593 _0725_/a_209_297# VGND 0.00923f 
C63594 _0725_/a_80_21# VGND 0.4368f 
C63595 net96 VGND 0.6013f
C63596 _1010_/a_1017_47# VGND 0.00404f 
C63597 _1010_/a_592_47# VGND 0.00748f 
C63598 _1010_/a_381_47# VGND 0.06508f 
C63599 _1010_/a_891_413# VGND 0.27442f 
C63600 _1010_/a_1059_315# VGND 0.38311f 
C63601 _1010_/a_466_413# VGND 0.21842f 
C63602 _1010_/a_634_159# VGND 0.25661f 
C63603 _1010_/a_193_47# VGND 0.3474f 
C63604 _1010_/a_27_47# VGND 0.59926f 
C63605 _0811_/a_384_47# VGND 0.00338f 
C63606 _0811_/a_299_297# VGND 0.03819f 
C63607 _0811_/a_81_21# VGND 0.30046f 
C63608 _0368_ VGND 0.64063f
C63609 _0742_/a_384_47# VGND 0.00373f 
C63610 _0742_/a_299_297# VGND 0.03987f 
C63611 _0742_/a_81_21# VGND 0.31983f 
C63612 clkbuf_1_0__f__0465_/a_110_47# VGND 2.29506f 
C63613 net23 VGND 4.43404f
C63614 B[15] VGND 0.93101f
C63615 input23/a_75_212# VGND 0.35175f 
C63616 rst VGND 0.71082f
C63617 input34/a_27_47# VGND 0.38435f 
C63618 A[5] VGND 0.60915f
C63619 input12/a_75_212# VGND 0.31292f 
C63620 _0304_ VGND 0.67208f
C63621 _0295_ VGND 0.64695f
C63622 _0673_/a_253_47# VGND 0.21301f 
C63623 _0673_/a_337_297# VGND 0 
C63624 _0673_/a_253_297# VGND 0 
C63625 _0673_/a_103_199# VGND 0.41107f 
C63626 _0475_ VGND 0.51799f
C63627 _0472_ VGND 0.70175f
C63628 _0473_ VGND 1.20362f
C63629 _0957_/a_304_297# VGND 0.00149f 
C63630 _0957_/a_220_297# VGND 0.00238f 
C63631 _0957_/a_114_297# VGND 0.003f 
C63632 _0957_/a_32_297# VGND 0.74267f 
C63633 _0690_/a_150_297# VGND 0 
C63634 _0690_/a_68_297# VGND 0.26076f 
C63635 net159 VGND 0.56238f
C63636 _0974_/a_448_47# VGND 0.20236f 
C63637 _0974_/a_544_297# VGND 0 
C63638 _0974_/a_222_93# VGND 0.22795f 
C63639 _0974_/a_79_199# VGND 0.22706f 
C63640 A[2] VGND 0.92823f
C63641 input9/a_27_47# VGND 0.38061f 
C63642 net67 VGND 2.21599f
C63643 _0089_ VGND 0.52812f
C63644 net77 VGND 0.64672f
C63645 _0991_/a_1017_47# VGND 0.00447f 
C63646 _0991_/a_592_47# VGND 0.00769f 
C63647 _0991_/a_975_413# VGND 0 
C63648 _0991_/a_561_413# VGND 0 
C63649 _0991_/a_381_47# VGND 0.06911f 
C63650 _0991_/a_891_413# VGND 0.31333f 
C63651 _0991_/a_1059_315# VGND 0.45181f 
C63652 _0991_/a_466_413# VGND 0.22346f 
C63653 _0991_/a_634_159# VGND 0.27665f 
C63654 _0991_/a_193_47# VGND 0.43949f 
C63655 _0991_/a_27_47# VGND 0.6201f 
C63656 _0709_/a_113_47# VGND 0.0017f 
C63657 net80 VGND 0.57884f
C63658 _0156_ VGND 0.49338f
C63659 net192 VGND 0.56792f
C63660 _0511_/a_384_47# VGND 0.00332f 
C63661 _0511_/a_299_297# VGND 0.06989f 
C63662 _0511_/a_81_21# VGND 0.34056f 
C63663 _0657_/a_109_297# VGND 0 
C63664 _0588_/a_113_47# VGND 0.00211f 
C63665 _0109_ VGND 0.90808f
C63666 net227 VGND 0.54466f
C63667 _0355_ VGND 0.41772f
C63668 _0354_ VGND 0.52997f
C63669 _0726_/a_240_47# VGND 0.18113f 
C63670 _0726_/a_149_47# VGND 0.14675f 
C63671 _0726_/a_512_297# VGND 0 
C63672 _0726_/a_245_297# VGND 0.00401f 
C63673 _0726_/a_51_297# VGND 0.38754f 
C63674 net57 VGND 1.33481f
C63675 net97 VGND 0.58594f
C63676 _1011_/a_1017_47# VGND 0.00496f 
C63677 _1011_/a_592_47# VGND 0.01067f 
C63678 _1011_/a_975_413# VGND 0 
C63679 _1011_/a_561_413# VGND 0.00179f 
C63680 _1011_/a_381_47# VGND 0.06634f 
C63681 _1011_/a_891_413# VGND 0.29818f 
C63682 _1011_/a_1059_315# VGND 0.41292f 
C63683 _1011_/a_466_413# VGND 0.24685f 
C63684 _1011_/a_634_159# VGND 0.28518f 
C63685 _1011_/a_193_47# VGND 0.38976f 
C63686 _1011_/a_27_47# VGND 0.60498f 
C63687 net99 VGND 0.39284f
C63688 clknet_0_clk VGND 2.93635f
C63689 clkbuf_1_0__f_clk/a_110_47# VGND 2.22027f 
C63690 net43 VGND 3.66702f
C63691 _0674_/a_113_47# VGND 0.00208f 
C63692 _0090_ VGND 0.55747f
C63693 _0422_ VGND 0.22123f
C63694 net217 VGND 0.56992f
C63695 _0812_/a_510_47# VGND 0.00928f 
C63696 _0812_/a_215_47# VGND 0.23443f 
C63697 _0812_/a_297_297# VGND 0 
C63698 _0812_/a_79_21# VGND 0.39408f 
C63699 net33 VGND 2.09498f
C63700 init VGND 0.5892f
C63701 input33/a_75_212# VGND 0.36707f 
C63702 net22 VGND 0.46645f
C63703 B[14] VGND 0.52346f
C63704 input22/a_75_212# VGND 0.373f 
C63705 A[4] VGND 0.55324f
C63706 input11/a_75_212# VGND 0.31112f 
C63707 net237 VGND 0.22969f
C63708 _0743_/a_240_47# VGND 0.16227f 
C63709 _0743_/a_149_47# VGND 0.1273f 
C63710 _0743_/a_245_297# VGND 0 
C63711 _0743_/a_51_297# VGND 0.28239f 
C63712 _0477_ VGND 0.68199f
C63713 _0958_/a_303_47# VGND 0.00352f 
C63714 _0958_/a_197_47# VGND 0.00361f 
C63715 _0958_/a_109_47# VGND 0.0017f 
C63716 _0958_/a_27_47# VGND 0.29617f 
C63717 _0691_/a_150_297# VGND 0 
C63718 _0691_/a_68_297# VGND 0.28276f 
C63719 _0382_ VGND 0.30668f
C63720 _0237_ VGND 1.54671f
C63721 _0381_ VGND 0.47026f
C63722 _0760_/a_285_47# VGND 0.21374f 
C63723 _0760_/a_129_47# VGND 0.00589f 
C63724 _0760_/a_377_297# VGND 0 
C63725 _0760_/a_47_47# VGND 0.32573f 
C63726 _0486_ VGND 0.63679f
C63727 control0.state\[2\] VGND 1.37225f
C63728 _0975_/a_145_75# VGND 0.00405f 
C63729 _0975_/a_59_75# VGND 0.31049f 
C63730 A[1] VGND 0.54412f
C63731 input8/a_75_212# VGND 0.37099f 
C63732 clkbuf_0__0460_/a_110_47# VGND 2.22613f 
C63733 _0992_/a_1017_47# VGND 0.00447f 
C63734 _0992_/a_592_47# VGND 0.0076f 
C63735 _0992_/a_561_413# VGND 0 
C63736 _0992_/a_381_47# VGND 0.06837f 
C63737 _0992_/a_891_413# VGND 0.29239f 
C63738 _0992_/a_1059_315# VGND 0.40499f 
C63739 _0992_/a_466_413# VGND 0.23994f 
C63740 _0992_/a_634_159# VGND 0.28307f 
C63741 _0992_/a_193_47# VGND 0.45166f 
C63742 _0992_/a_27_47# VGND 0.59267f 
C63743 net3 VGND 1.0183f
C63744 _0512_/a_373_47# VGND 0.00362f 
C63745 _0512_/a_109_47# VGND 0.00639f 
C63746 _0512_/a_109_297# VGND 0.00274f 
C63747 _0512_/a_27_297# VGND 0.43627f 
C63748 _0221_ VGND 1.49253f
C63749 _0589_/a_113_47# VGND 0.0019f 
C63750 _0658_/a_113_47# VGND 0.00171f 
C63751 _0356_ VGND 0.38836f
C63752 _0727_/a_277_47# VGND 0.00289f 
C63753 _0727_/a_193_47# VGND 0.0017f 
C63754 _0727_/a_109_47# VGND 0.00279f 
C63755 _1012_/a_1017_47# VGND 0.00447f 
C63756 _1012_/a_592_47# VGND 0.00748f 
C63757 _1012_/a_975_413# VGND 0 
C63758 _1012_/a_381_47# VGND 0.06714f 
C63759 _1012_/a_891_413# VGND 0.31504f 
C63760 _1012_/a_1059_315# VGND 0.44003f 
C63761 _1012_/a_466_413# VGND 0.22886f 
C63762 _1012_/a_634_159# VGND 0.28173f 
C63763 _1012_/a_193_47# VGND 0.49567f 
C63764 _1012_/a_27_47# VGND 0.65275f 
C63765 _0675_/a_150_297# VGND 0 
C63766 _0675_/a_68_297# VGND 0.2599f 
C63767 _0744_/a_27_47# VGND 0.81045f 
C63768 _0813_/a_109_297# VGND 0 
C63769 B[9] VGND 0.56438f
C63770 input32/a_75_212# VGND 0.35404f 
C63771 B[13] VGND 0.9596f
C63772 input21/a_75_212# VGND 0.36701f 
C63773 A[3] VGND 0.63297f
C63774 input10/a_75_212# VGND 0.37323f 
C63775 net95 VGND 0.40277f
C63776 _0470_ VGND 0.28323f
C63777 _0959_/a_300_47# VGND 0.0045f 
C63778 _0959_/a_472_297# VGND 0.00205f 
C63779 _0959_/a_217_297# VGND 0.00768f 
C63780 _0959_/a_80_21# VGND 0.55314f 
C63781 _0692_/a_113_47# VGND 0.00198f 
C63782 _0761_/a_113_47# VGND 0.002f 
C63783 _0087_ VGND 0.43464f
C63784 _0437_ VGND 0.97403f
C63785 net212 VGND 0.23762f
C63786 _0830_/a_510_47# VGND 0.00884f 
C63787 _0830_/a_215_47# VGND 0.22725f 
C63788 _0830_/a_297_297# VGND 0.00246f 
C63789 _0830_/a_79_21# VGND 0.35394f 
C63790 _0466_ VGND 3.12994f
C63791 _0488_ VGND 1.99945f
C63792 _0976_/a_439_47# VGND 0.00339f 
C63793 _0976_/a_218_47# VGND 0.00361f 
C63794 _0976_/a_535_374# VGND 0.00152f 
C63795 _0976_/a_218_374# VGND 0 
C63796 _0976_/a_505_21# VGND 0.38709f 
C63797 _0976_/a_76_199# VGND 0.2944f 
C63798 A[15] VGND 0.59553f
C63799 input7/a_75_212# VGND 0.36138f 
C63800 clkbuf_0__0461_/a_110_47# VGND 2.3496f 
C63801 _0993_/a_1017_47# VGND 0.00681f 
C63802 _0993_/a_592_47# VGND 0.00794f 
C63803 _0993_/a_975_413# VGND 0.00299f 
C63804 _0993_/a_561_413# VGND 0 
C63805 _0993_/a_381_47# VGND 0.06978f 
C63806 _0993_/a_891_413# VGND 0.35333f 
C63807 _0993_/a_1059_315# VGND 0.45083f 
C63808 _0993_/a_466_413# VGND 0.24555f 
C63809 _0993_/a_634_159# VGND 0.29f 
C63810 _0993_/a_193_47# VGND 0.52932f 
C63811 _0993_/a_27_47# VGND 0.66112f 
C63812 _0155_ VGND 0.20207f
C63813 _0188_ VGND 0.31741f
C63814 _0513_/a_384_47# VGND 0.00362f 
C63815 _0513_/a_299_297# VGND 0.05564f 
C63816 _0513_/a_81_21# VGND 0.31482f 
C63817 _0291_ VGND 1.20876f
C63818 acc0.A\[8\] VGND 2.39512f
C63819 net66 VGND 1.71835f
C63820 _0659_/a_150_297# VGND 0 
C63821 _0659_/a_68_297# VGND 0.26894f 
C63822 _0728_/a_145_75# VGND 0.00468f 
C63823 _0728_/a_59_75# VGND 0.2812f 
C63824 _1013_/a_1017_47# VGND 0.0049f 
C63825 _1013_/a_592_47# VGND 0.0082f 
C63826 _1013_/a_975_413# VGND 0 
C63827 _1013_/a_561_413# VGND 0 
C63828 _1013_/a_381_47# VGND 0.08425f 
C63829 _1013_/a_891_413# VGND 0.31874f 
C63830 _1013_/a_1059_315# VGND 0.43061f 
C63831 _1013_/a_466_413# VGND 0.23726f 
C63832 _1013_/a_634_159# VGND 0.27555f 
C63833 _1013_/a_193_47# VGND 0.44433f 
C63834 _1013_/a_27_47# VGND 0.67523f 
C63835 _0197_ VGND 0.27351f
C63836 _0530_/a_384_47# VGND 0.00332f 
C63837 _0530_/a_299_297# VGND 0.04007f 
C63838 _0530_/a_81_21# VGND 0.31758f 
C63839 _0307_ VGND 1.3395f
C63840 _0676_/a_113_47# VGND 0.00212f 
C63841 _0370_ VGND 0.47717f
C63842 _0745_/a_193_47# VGND 0.00118f 
C63843 _0745_/a_109_47# VGND 0 
C63844 _0814_/a_181_47# VGND 0.00276f 
C63845 _0814_/a_109_47# VGND 0.00215f 
C63846 _0814_/a_27_47# VGND 0.33641f 
C63847 net31 VGND 1.20673f
C63848 B[8] VGND 0.60926f
C63849 input31/a_75_212# VGND 0.358f 
C63850 B[12] VGND 0.52455f
C63851 input20/a_75_212# VGND 0.32734f 
C63852 _1030_/a_1017_47# VGND 0.00474f 
C63853 _1030_/a_592_47# VGND 0.00684f 
C63854 _1030_/a_975_413# VGND 0 
C63855 _1030_/a_561_413# VGND 0 
C63856 _1030_/a_381_47# VGND 0.08207f 
C63857 _1030_/a_891_413# VGND 0.28131f 
C63858 _1030_/a_1059_315# VGND 0.39576f 
C63859 _1030_/a_466_413# VGND 0.22428f 
C63860 _1030_/a_634_159# VGND 0.25447f 
C63861 _1030_/a_193_47# VGND 0.36929f 
C63862 _1030_/a_27_47# VGND 0.62217f 
C63863 _0693_/a_150_297# VGND 0 
C63864 _0693_/a_68_297# VGND 0.26794f 
C63865 _0383_ VGND 0.55681f
C63866 _0369_ VGND 10.68824f
C63867 _0762_/a_510_47# VGND 0.00993f 
C63868 _0762_/a_215_47# VGND 0.2446f 
C63869 _0762_/a_297_297# VGND 0.0033f 
C63870 _0762_/a_79_21# VGND 0.37018f 
C63871 _0253_ VGND 0.89715f
C63872 _0831_/a_285_47# VGND 0.0043f 
C63873 _0831_/a_285_297# VGND 0.00581f 
C63874 _0831_/a_117_297# VGND 0.00145f 
C63875 _0831_/a_35_297# VGND 0.41383f 
C63876 _0489_ VGND 0.29333f
C63877 _0977_/a_75_212# VGND 0.3309f 
C63878 A[14] VGND 0.72111f
C63879 input6/a_75_212# VGND 0.36415f 
C63880 _0462_ VGND 2.2254f
C63881 clkbuf_0__0462_/a_110_47# VGND 2.25327f 
C63882 _0994_/a_1017_47# VGND 0.00429f 
C63883 _0994_/a_592_47# VGND 0.00706f 
C63884 _0994_/a_975_413# VGND 0 
C63885 _0994_/a_561_413# VGND 0 
C63886 _0994_/a_381_47# VGND 0.06576f 
C63887 _0994_/a_891_413# VGND 0.29769f 
C63888 _0994_/a_1059_315# VGND 0.40354f 
C63889 _0994_/a_466_413# VGND 0.23443f 
C63890 _0994_/a_634_159# VGND 0.27168f 
C63891 _0994_/a_193_47# VGND 0.37722f 
C63892 _0994_/a_27_47# VGND 0.65838f 
C63893 net122 VGND 0.71283f
C63894 clknet_1_1__leaf__0463_ VGND 4.19661f
C63895 _0189_ VGND 0.46949f
C63896 net2 VGND 0.43236f
C63897 _0514_/a_373_47# VGND 0.00333f 
C63898 _0514_/a_109_47# VGND 0.00853f 
C63899 _0514_/a_109_297# VGND 0.01389f 
C63900 _0514_/a_27_297# VGND 0.47838f 
C63901 net71 VGND 0.79349f
C63902 clkbuf_1_1__f__0460_/a_110_47# VGND 2.22167f 
C63903 net242 VGND 0.30165f
C63904 _0729_/a_150_297# VGND 0 
C63905 _0729_/a_68_297# VGND 0.26173f 
C63906 acc0.A\[0\] VGND 0.38176f
C63907 net100 VGND 0.31302f
C63908 _1014_/a_1017_47# VGND 0.00429f 
C63909 _1014_/a_592_47# VGND 0.00858f 
C63910 _1014_/a_975_413# VGND 0 
C63911 _1014_/a_561_413# VGND 0 
C63912 _1014_/a_381_47# VGND 0.06121f 
C63913 _1014_/a_891_413# VGND 0.28305f 
C63914 _1014_/a_1059_315# VGND 0.38954f 
C63915 _1014_/a_466_413# VGND 0.23047f 
C63916 _1014_/a_634_159# VGND 0.28925f 
C63917 _1014_/a_193_47# VGND 0.37003f 
C63918 _1014_/a_27_47# VGND 0.61599f 
C63919 net9 VGND 5.21919f
C63920 net175 VGND 1.1309f
C63921 _0531_/a_373_47# VGND 0.00344f 
C63922 _0531_/a_109_47# VGND 0.00792f 
C63923 _0531_/a_109_297# VGND 0.00425f 
C63924 _0531_/a_27_297# VGND 0.44568f 
C63925 _0232_ VGND 0.48923f
C63926 _0223_ VGND 0.47267f
C63927 _0600_/a_253_47# VGND 0.21042f 
C63928 _0600_/a_337_297# VGND 0 
C63929 _0600_/a_253_297# VGND 0 
C63930 _0600_/a_103_199# VGND 0.29763f 
C63931 acc0.A\[17\] VGND 1.1082f
C63932 _0677_/a_285_47# VGND 0.22854f 
C63933 _0677_/a_129_47# VGND 0.0061f 
C63934 _0677_/a_377_297# VGND 0 
C63935 _0677_/a_47_47# VGND 0.35428f 
C63936 _0425_ VGND 0.17148f
C63937 _0401_ VGND 2.44242f
C63938 _0290_ VGND 1.77385f
C63939 _0423_ VGND 0.70412f
C63940 _0815_/a_199_47# VGND 0.00374f 
C63941 _0815_/a_113_297# VGND 0.04136f 
C63942 _0346_ VGND 9.61039f
C63943 _0746_/a_384_47# VGND 0.00355f 
C63944 _0746_/a_299_297# VGND 0.044f 
C63945 _0746_/a_81_21# VGND 0.30159f 
C63946 B[7] VGND 0.55007f
C63947 input30/a_75_212# VGND 0.37312f 
C63948 _1031_/a_1017_47# VGND 0.00415f 
C63949 _1031_/a_592_47# VGND 0.00734f 
C63950 _1031_/a_975_413# VGND 0 
C63951 _1031_/a_561_413# VGND 0 
C63952 _1031_/a_381_47# VGND 0.06938f 
C63953 _1031_/a_891_413# VGND 0.2896f 
C63954 _1031_/a_1059_315# VGND 0.4208f 
C63955 _1031_/a_466_413# VGND 0.21691f 
C63956 _1031_/a_634_159# VGND 0.25903f 
C63957 _1031_/a_193_47# VGND 0.38108f 
C63958 _1031_/a_27_47# VGND 0.63204f 
C63959 _0326_ VGND 0.77167f
C63960 _0325_ VGND 0.36139f
C63961 _0694_/a_113_47# VGND 0.00172f 
C63962 _0439_ VGND 0.31452f
C63963 _0438_ VGND 0.77699f
C63964 _0832_/a_113_47# VGND 0.00196f 
C63965 _0384_ VGND 0.40724f
C63966 _0763_/a_193_47# VGND 0.00139f 
C63967 _0763_/a_109_47# VGND 0 
C63968 _0978_/a_373_47# VGND 0.00231f 
C63969 _0978_/a_109_47# VGND 0.01133f 
C63970 _0978_/a_109_297# VGND 0.00998f 
C63971 _0978_/a_27_297# VGND 0.45497f 
C63972 A[13] VGND 0.6515f
C63973 input5/a_75_212# VGND 0.37617f 
C63974 _0397_ VGND 1.08682f
C63975 _0780_/a_285_47# VGND 0.00684f 
C63976 _0780_/a_285_297# VGND 0.00562f 
C63977 _0780_/a_117_297# VGND 0.00141f 
C63978 _0780_/a_35_297# VGND 0.4604f 
C63979 _0463_ VGND 0.82437f
C63980 clkbuf_0__0463_/a_110_47# VGND 2.2263f 
C63981 _0995_/a_1017_47# VGND 0.00456f 
C63982 _0995_/a_592_47# VGND 0.00782f 
C63983 _0995_/a_975_413# VGND 0 
C63984 _0995_/a_561_413# VGND 0 
C63985 _0995_/a_381_47# VGND 0.06253f 
C63986 _0995_/a_891_413# VGND 0.29352f 
C63987 _0995_/a_1059_315# VGND 0.41217f 
C63988 _0995_/a_466_413# VGND 0.22177f 
C63989 _0995_/a_634_159# VGND 0.27008f 
C63990 _0995_/a_193_47# VGND 0.44494f 
C63991 _0995_/a_27_47# VGND 0.56988f 
C63992 net181 VGND 0.58829f
C63993 _0515_/a_384_47# VGND 0.00346f 
C63994 _0515_/a_299_297# VGND 0.04058f 
C63995 _0515_/a_81_21# VGND 0.30488f 
C63996 clkbuf_1_1__f__0461_/a_110_47# VGND 2.1993f 
C63997 _0113_ VGND 0.62415f
C63998 _1015_/a_1017_47# VGND 0.00457f 
C63999 _1015_/a_592_47# VGND 0.00774f 
C64000 _1015_/a_975_413# VGND 0 
C64001 _1015_/a_561_413# VGND 0 
C64002 _1015_/a_381_47# VGND 0.06665f 
C64003 _1015_/a_891_413# VGND 0.28864f 
C64004 _1015_/a_1059_315# VGND 0.40121f 
C64005 _1015_/a_466_413# VGND 0.22056f 
C64006 _1015_/a_634_159# VGND 0.26079f 
C64007 _1015_/a_193_47# VGND 0.35656f 
C64008 _1015_/a_27_47# VGND 0.60414f 
C64009 _0146_ VGND 0.52547f
C64010 _0198_ VGND 0.27778f
C64011 _0532_/a_384_47# VGND 0.00322f 
C64012 _0532_/a_299_297# VGND 0.03897f 
C64013 _0532_/a_81_21# VGND 0.31294f 
C64014 _0601_/a_150_297# VGND 0 
C64015 _0601_/a_68_297# VGND 0.29465f 
C64016 _0309_ VGND 0.72881f
C64017 _0678_/a_150_297# VGND 0 
C64018 _0678_/a_68_297# VGND 0.27014f 
C64019 _0104_ VGND 0.40492f
C64020 _0371_ VGND 0.17873f
C64021 net216 VGND 0.2071f
C64022 _0747_/a_510_47# VGND 0.00777f 
C64023 _0747_/a_215_47# VGND 0.23162f 
C64024 _0747_/a_79_21# VGND 0.34218f 
C64025 _0426_ VGND 0.28601f
C64026 _0816_/a_150_297# VGND 0 
C64027 _0816_/a_68_297# VGND 0.28709f 
C64028 net202 VGND 0.5579f
C64029 _1032_/a_1017_47# VGND 0.00475f 
C64030 _1032_/a_592_47# VGND 0.00822f 
C64031 _1032_/a_975_413# VGND 0 
C64032 _1032_/a_561_413# VGND 0 
C64033 _1032_/a_381_47# VGND 0.07121f 
C64034 _1032_/a_891_413# VGND 0.3032f 
C64035 _1032_/a_1059_315# VGND 0.42805f 
C64036 _1032_/a_466_413# VGND 0.24381f 
C64037 _1032_/a_634_159# VGND 0.2767f 
C64038 _1032_/a_193_47# VGND 0.49416f 
C64039 _1032_/a_27_47# VGND 0.61192f 
C64040 _0327_ VGND 0.5261f
C64041 _0323_ VGND 0.28963f
C64042 _0312_ VGND 1.48639f
C64043 _0695_/a_300_47# VGND 0.00413f 
C64044 _0695_/a_217_297# VGND 0.00163f 
C64045 _0695_/a_80_21# VGND 0.50928f 
C64046 _0764_/a_384_47# VGND 0.00349f 
C64047 _0764_/a_299_297# VGND 0.04595f 
C64048 _0764_/a_81_21# VGND 0.34427f 
C64049 _0086_ VGND 0.40771f
C64050 net235 VGND 0.42469f
C64051 _0833_/a_510_47# VGND 0.00842f 
C64052 _0833_/a_215_47# VGND 0.23755f 
C64053 _0833_/a_297_297# VGND 0 
C64054 _0833_/a_79_21# VGND 0.35369f 
C64055 _0902_/a_27_47# VGND 0.38601f 
C64056 _0169_ VGND 0.47402f
C64057 net164 VGND 0.2156f
C64058 _0480_ VGND 0.71838f
C64059 _0979_/a_373_47# VGND 0.00227f 
C64060 _0979_/a_109_47# VGND 0.00712f 
C64061 _0979_/a_109_297# VGND 0.00773f 
C64062 _0979_/a_27_297# VGND 0.45722f 
C64063 A[12] VGND 0.23364f
C64064 input4/a_75_212# VGND 0.34588f 
C64065 _0781_/a_150_297# VGND 0 
C64066 _0781_/a_68_297# VGND 0.27826f 
C64067 _0850_/a_150_297# VGND 0 
C64068 _0850_/a_68_297# VGND 0.26497f 
C64069 clknet_0__0464_ VGND 3.38749f
C64070 clkbuf_0__0464_/a_110_47# VGND 2.26156f 
C64071 _0996_/a_1017_47# VGND 0.00404f 
C64072 _0996_/a_592_47# VGND 0.0074f 
C64073 _0996_/a_381_47# VGND 0.06538f 
C64074 _0996_/a_891_413# VGND 0.29152f 
C64075 _0996_/a_1059_315# VGND 0.40031f 
C64076 _0996_/a_466_413# VGND 0.21922f 
C64077 _0996_/a_634_159# VGND 0.25465f 
C64078 _0996_/a_193_47# VGND 0.34928f 
C64079 _0996_/a_27_47# VGND 0.59414f 
C64080 _0190_ VGND 0.38111f
C64081 net16 VGND 0.58926f
C64082 _0516_/a_373_47# VGND 0.00288f 
C64083 _0516_/a_109_47# VGND 0.00863f 
C64084 _0516_/a_109_297# VGND 0.00604f 
C64085 _0516_/a_27_297# VGND 0.45062f 
C64086 clkbuf_1_1__f__0462_/a_110_47# VGND 2.2613f 
C64087 net166 VGND 0.30499f
C64088 _1016_/a_1017_47# VGND 0.00447f 
C64089 _1016_/a_592_47# VGND 0.01067f 
C64090 _1016_/a_975_413# VGND 0 
C64091 _1016_/a_561_413# VGND 0.00179f 
C64092 _1016_/a_381_47# VGND 0.06182f 
C64093 _1016_/a_891_413# VGND 0.28472f 
C64094 _1016_/a_1059_315# VGND 0.3951f 
C64095 _1016_/a_466_413# VGND 0.24966f 
C64096 _1016_/a_634_159# VGND 0.2853f 
C64097 _1016_/a_193_47# VGND 0.36988f 
C64098 _1016_/a_27_47# VGND 0.61745f 
C64099 _0199_ VGND 0.80853f
C64100 net8 VGND 1.36639f
C64101 _0180_ VGND 4.07923f
C64102 _0182_ VGND 1.53365f
C64103 acc0.A\[1\] VGND 1.98373f
C64104 _0533_/a_373_47# VGND 0.00212f 
C64105 _0533_/a_109_47# VGND 0.00618f 
C64106 _0533_/a_109_297# VGND 0.00274f 
C64107 _0533_/a_27_297# VGND 0.4245f 
C64108 _0602_/a_113_47# VGND 0.00195f 
C64109 _0310_ VGND 0.58489f
C64110 _0679_/a_150_297# VGND 0 
C64111 _0679_/a_68_297# VGND 0.28066f 
C64112 _0294_ VGND 2.08514f
C64113 _0748_/a_384_47# VGND 0.00325f 
C64114 _0748_/a_299_297# VGND 0.05528f 
C64115 _0748_/a_81_21# VGND 0.30898f 
C64116 _0424_ VGND 0.37956f
C64117 _0817_/a_585_47# VGND 0 
C64118 _0817_/a_266_47# VGND 0.20397f 
C64119 _0817_/a_368_297# VGND 0 
C64120 _0817_/a_266_297# VGND 0 
C64121 _0817_/a_81_21# VGND 0.35942f 
C64122 comp0.B\[1\] VGND 0.63772f
C64123 _0131_ VGND 0.86733f
C64124 net119 VGND 0.43955f
C64125 _1033_/a_1017_47# VGND 0.00486f 
C64126 _1033_/a_592_47# VGND 0.00816f 
C64127 _1033_/a_975_413# VGND 0 
C64128 _1033_/a_561_413# VGND 0 
C64129 _1033_/a_381_47# VGND 0.07048f 
C64130 _1033_/a_891_413# VGND 0.29774f 
C64131 _1033_/a_1059_315# VGND 0.41178f 
C64132 _1033_/a_466_413# VGND 0.22741f 
C64133 _1033_/a_634_159# VGND 0.27232f 
C64134 _1033_/a_193_47# VGND 0.47621f 
C64135 _1033_/a_27_47# VGND 0.588f 
C64136 _0137_ VGND 0.40869f
C64137 _0172_ VGND 5.47054f
C64138 net30 VGND 0.29811f
C64139 net180 VGND 0.35187f
C64140 _0550_/a_240_47# VGND 0.16106f 
C64141 _0550_/a_149_47# VGND 0.12503f 
C64142 _0550_/a_51_297# VGND 0.28961f 
C64143 net106 VGND 0.87016f
C64144 _0385_ VGND 0.60255f
C64145 net220 VGND 0.43998f
C64146 _0765_/a_510_47# VGND 0.00636f 
C64147 _0765_/a_215_47# VGND 0.22534f 
C64148 _0765_/a_297_297# VGND 0 
C64149 _0765_/a_79_21# VGND 0.36326f 
C64150 _0328_ VGND 2.74593f
C64151 _0696_/a_109_297# VGND 0 
C64152 _0433_ VGND 0.78765f
C64153 _0834_/a_109_297# VGND 0 
C64154 acc0.A\[4\] VGND 2.57858f
C64155 net136 VGND 0.30832f
C64156 _1050_/a_1017_47# VGND 0.00404f 
C64157 _1050_/a_592_47# VGND 0.00662f 
C64158 _1050_/a_381_47# VGND 0.06058f 
C64159 _1050_/a_891_413# VGND 0.27478f 
C64160 _1050_/a_1059_315# VGND 0.38365f 
C64161 _1050_/a_466_413# VGND 0.21262f 
C64162 _1050_/a_634_159# VGND 0.25177f 
C64163 _1050_/a_193_47# VGND 0.34318f 
C64164 _1050_/a_27_47# VGND 0.58466f 
C64165 A[11] VGND 0.42991f
C64166 input3/a_75_212# VGND 0.35867f 
C64167 net111 VGND 0.78902f
C64168 _0782_/a_27_47# VGND 0.67831f 
C64169 _0453_ VGND 0.49928f
C64170 _0266_ VGND 0.48385f
C64171 _0452_ VGND 0.48601f
C64172 _0851_/a_113_47# VGND 0.00198f 
C64173 clknet_0__0465_ VGND 3.00041f
C64174 clkbuf_0__0465_/a_110_47# VGND 2.25243f 
C64175 _0997_/a_1017_47# VGND 0.00681f 
C64176 _0997_/a_592_47# VGND 0.00789f 
C64177 _0997_/a_975_413# VGND 0.00238f 
C64178 _0997_/a_561_413# VGND 0 
C64179 _0997_/a_381_47# VGND 0.06346f 
C64180 _0997_/a_891_413# VGND 0.31555f 
C64181 _0997_/a_1059_315# VGND 0.43043f 
C64182 _0997_/a_466_413# VGND 0.22499f 
C64183 _0997_/a_634_159# VGND 0.27536f 
C64184 _0997_/a_193_47# VGND 0.4023f 
C64185 _0997_/a_27_47# VGND 0.62367f 
C64186 _0153_ VGND 0.36106f
C64187 _0517_/a_384_47# VGND 0.00372f 
C64188 _0517_/a_299_297# VGND 0.04064f 
C64189 _0517_/a_81_21# VGND 0.31467f 
C64190 clknet_0__0463_ VGND 3.3157f
C64191 clkbuf_1_1__f__0463_/a_110_47# VGND 2.24289f 
C64192 net103 VGND 0.74285f
C64193 _1017_/a_1017_47# VGND 0.00447f 
C64194 _1017_/a_592_47# VGND 0.00824f 
C64195 _1017_/a_561_413# VGND 0.00129f 
C64196 _1017_/a_381_47# VGND 0.08287f 
C64197 _1017_/a_891_413# VGND 0.28597f 
C64198 _1017_/a_1059_315# VGND 0.40099f 
C64199 _1017_/a_466_413# VGND 0.23642f 
C64200 _1017_/a_634_159# VGND 0.26442f 
C64201 _1017_/a_193_47# VGND 0.39658f 
C64202 _1017_/a_27_47# VGND 0.60924f 
C64203 _0603_/a_150_297# VGND 0 
C64204 _0603_/a_68_297# VGND 0.29647f 
C64205 _0534_/a_384_47# VGND 0.00328f 
C64206 _0534_/a_299_297# VGND 0.03802f 
C64207 _0534_/a_81_21# VGND 0.2982f 
C64208 _0372_ VGND 1.04148f
C64209 _0248_ VGND 1.21429f
C64210 _0749_/a_384_47# VGND 0.00343f 
C64211 _0749_/a_299_297# VGND 0.04522f 
C64212 _0749_/a_81_21# VGND 0.31932f 
C64213 _0818_/a_193_47# VGND 0 
C64214 _0818_/a_109_47# VGND 0 
C64215 comp0.B\[2\] VGND 0.94557f
C64216 _1034_/a_1017_47# VGND 0.00662f 
C64217 _1034_/a_592_47# VGND 0.00832f 
C64218 _1034_/a_975_413# VGND 0.00167f 
C64219 _1034_/a_561_413# VGND 0 
C64220 _1034_/a_381_47# VGND 0.06993f 
C64221 _1034_/a_891_413# VGND 0.32021f 
C64222 _1034_/a_1059_315# VGND 0.42265f 
C64223 _1034_/a_466_413# VGND 0.22558f 
C64224 _1034_/a_634_159# VGND 0.27435f 
C64225 _1034_/a_193_47# VGND 0.50185f 
C64226 _1034_/a_27_47# VGND 0.60958f 
C64227 _0551_/a_27_47# VGND 0.40162f 
C64228 _0252_ VGND 0.92227f
C64229 acc0.A\[7\] VGND 0.82411f
C64230 net65 VGND 2.32682f
C64231 _0620_/a_113_47# VGND 0.00173f 
C64232 _0329_ VGND 0.42485f
C64233 _0322_ VGND 0.77152f
C64234 _0697_/a_300_47# VGND 0.0057f 
C64235 _0697_/a_472_297# VGND 0 
C64236 _0697_/a_217_297# VGND 0.00197f 
C64237 _0697_/a_80_21# VGND 0.54489f 
C64238 _0766_/a_109_297# VGND 0 
C64239 _0255_ VGND 1.03463f
C64240 _0835_/a_215_47# VGND 0.3027f 
C64241 _0835_/a_493_297# VGND 0 
C64242 _0835_/a_292_297# VGND 0.00162f 
C64243 _0835_/a_78_199# VGND 0.26286f 
C64244 acc0.A\[5\] VGND 1.7864f
C64245 _0149_ VGND 0.39208f
C64246 net137 VGND 0.47064f
C64247 _1051_/a_1017_47# VGND 0.00447f 
C64248 _1051_/a_592_47# VGND 0.00748f 
C64249 _1051_/a_381_47# VGND 0.06139f 
C64250 _1051_/a_891_413# VGND 0.28312f 
C64251 _1051_/a_1059_315# VGND 0.40616f 
C64252 _1051_/a_466_413# VGND 0.21771f 
C64253 _1051_/a_634_159# VGND 0.25863f 
C64254 _1051_/a_193_47# VGND 0.34676f 
C64255 _1051_/a_27_47# VGND 0.59067f 
C64256 A[10] VGND 0.91296f
C64257 input2/a_75_212# VGND 0.33019f 
C64258 _0096_ VGND 0.59978f
C64259 _0399_ VGND 7.75486f
C64260 _0398_ VGND 0.48397f
C64261 _0783_/a_510_47# VGND 0.00622f 
C64262 _0783_/a_215_47# VGND 0.22879f 
C64263 _0783_/a_297_297# VGND 0 
C64264 _0783_/a_79_21# VGND 0.40769f 
C64265 _0852_/a_285_47# VGND 0.00527f 
C64266 _0852_/a_285_297# VGND 0.00137f 
C64267 _0852_/a_117_297# VGND 0 
C64268 _0852_/a_35_297# VGND 0.42171f 
C64269 net84 VGND 0.66308f
C64270 _0998_/a_1017_47# VGND 0.00447f 
C64271 _0998_/a_592_47# VGND 0.00748f 
C64272 _0998_/a_975_413# VGND 0 
C64273 _0998_/a_381_47# VGND 0.06542f 
C64274 _0998_/a_891_413# VGND 0.29071f 
C64275 _0998_/a_1059_315# VGND 0.41229f 
C64276 _0998_/a_466_413# VGND 0.22037f 
C64277 _0998_/a_634_159# VGND 0.26943f 
C64278 _0998_/a_193_47# VGND 0.4032f 
C64279 _0998_/a_27_47# VGND 0.59856f 
C64280 _0191_ VGND 0.40856f
C64281 net15 VGND 0.39002f
C64282 _0518_/a_373_47# VGND 0.00257f 
C64283 _0518_/a_109_47# VGND 0.00812f 
C64284 _0518_/a_109_297# VGND 0.01035f 
C64285 _0518_/a_27_297# VGND 0.45329f 
C64286 clkbuf_1_1__f__0464_/a_110_47# VGND 2.46855f 
C64287 net104 VGND 0.78899f
C64288 _1018_/a_1017_47# VGND 0.00404f 
C64289 _1018_/a_592_47# VGND 0.00662f 
C64290 _1018_/a_381_47# VGND 0.06079f 
C64291 _1018_/a_891_413# VGND 0.27607f 
C64292 _1018_/a_1059_315# VGND 0.40156f 
C64293 _1018_/a_466_413# VGND 0.21592f 
C64294 _1018_/a_634_159# VGND 0.2536f 
C64295 _1018_/a_193_47# VGND 0.36279f 
C64296 _1018_/a_27_47# VGND 0.59374f 
C64297 comp0.B\[14\] VGND 0.90608f
C64298 _0535_/a_150_297# VGND 0 
C64299 _0535_/a_68_297# VGND 0.26834f 
C64300 _0235_ VGND 0.38562f
C64301 _0604_/a_113_47# VGND 0.00178f 
C64302 _0428_ VGND 0.30121f
C64303 _0427_ VGND 0.43549f
C64304 _0819_/a_384_47# VGND 0.00366f 
C64305 _0819_/a_299_297# VGND 0.03805f 
C64306 _0819_/a_81_21# VGND 0.31875f 
C64307 _0133_ VGND 1.01935f
C64308 net121 VGND 0.53746f
C64309 _1035_/a_1017_47# VGND 0.00475f 
C64310 _1035_/a_592_47# VGND 0.00822f 
C64311 _1035_/a_975_413# VGND 0 
C64312 _1035_/a_561_413# VGND 0 
C64313 _1035_/a_381_47# VGND 0.07235f 
C64314 _1035_/a_891_413# VGND 0.30037f 
C64315 _1035_/a_1059_315# VGND 0.41311f 
C64316 _1035_/a_466_413# VGND 0.22692f 
C64317 _1035_/a_634_159# VGND 0.2757f 
C64318 _1035_/a_193_47# VGND 0.39373f 
C64319 _1035_/a_27_47# VGND 0.6241f 
C64320 _0209_ VGND 0.28274f
C64321 _0552_/a_150_297# VGND 0 
C64322 _0552_/a_68_297# VGND 0.26988f 
C64323 _0621_/a_285_47# VGND 0.0055f 
C64324 _0621_/a_285_297# VGND 0.00238f 
C64325 _0621_/a_117_297# VGND 0 
C64326 _0621_/a_35_297# VGND 0.44723f 
C64327 _0330_ VGND 0.42645f
C64328 _0317_ VGND 1.26103f
C64329 _0698_/a_199_47# VGND 0.00394f 
C64330 _0698_/a_113_297# VGND 0.03986f 
C64331 _0387_ VGND 1.34549f
C64332 _0767_/a_145_75# VGND 0.00504f 
C64333 _0767_/a_59_75# VGND 0.33933f 
C64334 _0836_/a_150_297# VGND 0 
C64335 _0836_/a_68_297# VGND 0.2654f 
C64336 _1052_/a_1017_47# VGND 0.00423f 
C64337 _1052_/a_592_47# VGND 0.00685f 
C64338 _1052_/a_975_413# VGND 0 
C64339 _1052_/a_561_413# VGND 0 
C64340 _1052_/a_381_47# VGND 0.06285f 
C64341 _1052_/a_891_413# VGND 0.2832f 
C64342 _1052_/a_1059_315# VGND 0.39533f 
C64343 _1052_/a_466_413# VGND 0.21526f 
C64344 _1052_/a_634_159# VGND 0.25636f 
C64345 _1052_/a_193_47# VGND 0.36111f 
C64346 _1052_/a_27_47# VGND 0.60872f 
C64347 net1 VGND 4.2664f
C64348 A[0] VGND 0.69385f
C64349 input1/a_27_47# VGND 0.37778f 
C64350 _0784_/a_113_47# VGND 0.00194f 
C64351 _0853_/a_150_297# VGND 0 
C64352 _0853_/a_68_297# VGND 0.28056f 
C64353 net85 VGND 0.62029f
C64354 _0999_/a_1017_47# VGND 0.00465f 
C64355 _0999_/a_592_47# VGND 0.00774f 
C64356 _0999_/a_975_413# VGND 0 
C64357 _0999_/a_561_413# VGND 0 
C64358 _0999_/a_381_47# VGND 0.06648f 
C64359 _0999_/a_891_413# VGND 0.30444f 
C64360 _0999_/a_1059_315# VGND 0.40374f 
C64361 _0999_/a_466_413# VGND 0.22046f 
C64362 _0999_/a_634_159# VGND 0.26094f 
C64363 _0999_/a_193_47# VGND 0.35456f 
C64364 _0999_/a_27_47# VGND 0.6017f 
C64365 _0152_ VGND 0.19684f
C64366 _0519_/a_384_47# VGND 0.00326f 
C64367 _0519_/a_299_297# VGND 0.03826f 
C64368 _0519_/a_81_21# VGND 0.30012f 
C64369 clkbuf_1_1__f__0465_/a_110_47# VGND 2.38613f 
C64370 net207 VGND 0.42165f
C64371 net105 VGND 0.70406f
C64372 _1019_/a_1017_47# VGND 0.00468f 
C64373 _1019_/a_592_47# VGND 0.00808f 
C64374 _1019_/a_975_413# VGND 0 
C64375 _1019_/a_561_413# VGND 0 
C64376 _1019_/a_381_47# VGND 0.06819f 
C64377 _1019_/a_891_413# VGND 0.29765f 
C64378 _1019_/a_1059_315# VGND 0.4093f 
C64379 _1019_/a_466_413# VGND 0.22483f 
C64380 _1019_/a_634_159# VGND 0.27192f 
C64381 _1019_/a_193_47# VGND 0.4492f 
C64382 _1019_/a_27_47# VGND 0.60665f 
C64383 _0228_ VGND 0.6602f
C64384 _0605_/a_109_297# VGND 0 
C64385 _0144_ VGND 0.45525f
C64386 _0200_ VGND 0.34635f
C64387 _0536_/a_240_47# VGND 0.18211f 
C64388 _0536_/a_149_47# VGND 0.13453f 
C64389 _0536_/a_512_297# VGND 0 
C64390 _0536_/a_245_297# VGND 0.00123f 
C64391 _0536_/a_51_297# VGND 0.29962f 
C64392 comp0.B\[4\] VGND 1.38442f
C64393 net161 VGND 0.39974f
C64394 _1036_/a_1017_47# VGND 0.00486f 
C64395 _1036_/a_592_47# VGND 0.00791f 
C64396 _1036_/a_975_413# VGND 0 
C64397 _1036_/a_561_413# VGND 0 
C64398 _1036_/a_381_47# VGND 0.06665f 
C64399 _1036_/a_891_413# VGND 0.29891f 
C64400 _1036_/a_1059_315# VGND 0.40929f 
C64401 _1036_/a_466_413# VGND 0.22558f 
C64402 _1036_/a_634_159# VGND 0.2713f 
C64403 _1036_/a_193_47# VGND 0.46747f 
C64404 _1036_/a_27_47# VGND 0.6122f 
C64405 _0136_ VGND 1.1608f
C64406 _0174_ VGND 2.52485f
C64407 _0553_/a_240_47# VGND 0.16104f 
C64408 _0553_/a_149_47# VGND 0.125f 
C64409 _0553_/a_51_297# VGND 0.28349f 
C64410 _0622_/a_193_47# VGND 0.00171f 
C64411 _0622_/a_109_47# VGND 0.00108f 
C64412 _0331_ VGND 0.6693f
C64413 net56 VGND 1.00535f
C64414 _0699_/a_150_297# VGND 0 
C64415 _0699_/a_68_297# VGND 0.28232f 
C64416 _0768_/a_27_47# VGND 0.22545f 
C64417 _0768_/a_109_297# VGND 0 
C64418 _0442_ VGND 0.53822f
C64419 _0441_ VGND 0.21998f
C64420 _0440_ VGND 0.5235f
C64421 _0837_/a_585_47# VGND 0.00111f 
C64422 _0837_/a_266_47# VGND 0.20836f 
C64423 _0837_/a_266_297# VGND 0 
C64424 _0837_/a_81_21# VGND 0.34878f 
C64425 net139 VGND 0.56645f
C64426 _1053_/a_1017_47# VGND 0.00462f 
C64427 _1053_/a_592_47# VGND 0.0077f 
C64428 _1053_/a_975_413# VGND 0 
C64429 _1053_/a_561_413# VGND 0 
C64430 _1053_/a_381_47# VGND 0.0685f 
C64431 _1053_/a_891_413# VGND 0.29203f 
C64432 _1053_/a_1059_315# VGND 0.38982f 
C64433 _1053_/a_466_413# VGND 0.2256f 
C64434 _1053_/a_634_159# VGND 0.2693f 
C64435 _1053_/a_193_47# VGND 0.46832f 
C64436 _1053_/a_27_47# VGND 0.61057f 
C64437 _0126_ VGND 0.22729f
C64438 net190 VGND 1.27814f
C64439 net197 VGND 0.43004f
C64440 _0570_/a_373_47# VGND 0.00288f 
C64441 _0570_/a_109_47# VGND 0.00764f 
C64442 _0570_/a_109_297# VGND 0.00274f 
C64443 _0570_/a_27_297# VGND 0.43687f 
C64444 hold19/a_391_47# VGND 0.2666f 
C64445 hold19/a_285_47# VGND 0.4548f 
C64446 hold19/a_49_47# VGND 0.47666f 
C64447 _0785_/a_384_47# VGND 0.00324f 
C64448 _0785_/a_299_297# VGND 0.03806f 
C64449 _0785_/a_81_21# VGND 0.29836f 
C64450 _0081_ VGND 0.52878f
C64451 _0455_ VGND 0.39509f
C64452 _0454_ VGND 0.38737f
C64453 _0854_/a_510_47# VGND 0.00781f 
C64454 _0854_/a_215_47# VGND 0.23164f 
C64455 _0854_/a_79_21# VGND 0.35052f 
C64456 net133 VGND 0.77101f
C64457 clknet_1_0__leaf__0464_ VGND 3.80095f
C64458 control0.count\[1\] VGND 1.83271f
C64459 _0168_ VGND 0.73707f
C64460 VPWR VGND 1.40324p
C64461 _1070_/a_1017_47# VGND 0.00447f 
C64462 _1070_/a_592_47# VGND 0.00748f 
C64463 _1070_/a_975_413# VGND 0 
C64464 _1070_/a_381_47# VGND 0.07232f 
C64465 _1070_/a_891_413# VGND 0.30918f 
C64466 _1070_/a_1059_315# VGND 0.42448f 
C64467 _1070_/a_466_413# VGND 0.22374f 
C64468 _1070_/a_634_159# VGND 0.26919f 
C64469 _1070_/a_193_47# VGND 0.50781f 
C64470 _1070_/a_27_47# VGND 0.65183f 
C64471 net138 VGND 0.40277f
C64472 net76 VGND 0.6065f
C64473 _0537_/a_150_297# VGND 0 
C64474 _0537_/a_68_297# VGND 0.27283f 
C64475 _0238_ VGND 2.04588f
C64476 _0236_ VGND 0.73332f
C64477 _0606_/a_465_297# VGND 0 
C64478 _0606_/a_392_297# VGND 0 
C64479 _0606_/a_297_297# VGND 0 
C64480 _0606_/a_109_53# VGND 0.27354f 
C64481 _0606_/a_215_297# VGND 0.39719f 
C64482 net87 VGND 0.37982f
C64483 clknet_1_0__leaf__0459_ VGND 4.31124f
C64484 _0135_ VGND 0.62713f
C64485 _1037_/a_1017_47# VGND 0.00447f 
C64486 _1037_/a_592_47# VGND 0.00748f 
C64487 _1037_/a_975_413# VGND 0 
C64488 _1037_/a_381_47# VGND 0.06718f 
C64489 _1037_/a_891_413# VGND 0.2872f 
C64490 _1037_/a_1059_315# VGND 0.39719f 
C64491 _1037_/a_466_413# VGND 0.21939f 
C64492 _1037_/a_634_159# VGND 0.26786f 
C64493 _1037_/a_193_47# VGND 0.3723f 
C64494 _1037_/a_27_47# VGND 0.6177f 
C64495 _0210_ VGND 0.36893f
C64496 net160 VGND 0.6635f
C64497 _0554_/a_150_297# VGND 0 
C64498 _0554_/a_68_297# VGND 0.27388f 
C64499 net63 VGND 1.3306f
C64500 _0623_/a_109_297# VGND 0 
C64501 _0838_/a_109_297# VGND 0 
C64502 _0388_ VGND 0.47237f
C64503 _0386_ VGND 0.56959f
C64504 _0244_ VGND 2.24061f
C64505 _0769_/a_384_47# VGND 0.00362f 
C64506 _0769_/a_299_297# VGND 0.03991f 
C64507 _0769_/a_81_21# VGND 0.30746f 
C64508 net169 VGND 0.27738f
C64509 net140 VGND 0.45608f
C64510 _1054_/a_1017_47# VGND 0.004f 
C64511 _1054_/a_592_47# VGND 0.00688f 
C64512 _1054_/a_975_413# VGND 0 
C64513 _1054_/a_561_413# VGND 0 
C64514 _1054_/a_381_47# VGND 0.06157f 
C64515 _1054_/a_891_413# VGND 0.27999f 
C64516 _1054_/a_1059_315# VGND 0.39859f 
C64517 _1054_/a_466_413# VGND 0.21501f 
C64518 _1054_/a_634_159# VGND 0.25413f 
C64519 _1054_/a_193_47# VGND 0.34957f 
C64520 _1054_/a_27_47# VGND 0.56017f 
C64521 _0125_ VGND 0.48932f
C64522 acc0.A\[27\] VGND 2.84831f
C64523 _0571_/a_373_47# VGND 0.00288f 
C64524 _0571_/a_109_47# VGND 0.00795f 
C64525 _0571_/a_109_297# VGND 0.00274f 
C64526 _0571_/a_27_297# VGND 0.43808f 
C64527 _0254_ VGND 0.80745f
C64528 _0640_/a_465_297# VGND 0 
C64529 _0640_/a_392_297# VGND 0 
C64530 _0640_/a_297_297# VGND 0 
C64531 _0640_/a_109_53# VGND 0.26762f 
C64532 _0640_/a_215_297# VGND 0.3569f 
C64533 net176 VGND 0.29688f
C64534 hold29/a_391_47# VGND 0.24706f 
C64535 hold29/a_285_47# VGND 0.40884f 
C64536 hold29/a_49_47# VGND 0.47988f 
C64537 hold18/a_391_47# VGND 0.25403f 
C64538 hold18/a_285_47# VGND 0.42276f 
C64539 hold18/a_49_47# VGND 0.47023f 
C64540 _0402_ VGND 1.47601f
C64541 _0786_/a_300_47# VGND 0.00431f 
C64542 _0786_/a_472_297# VGND 0 
C64543 _0786_/a_217_297# VGND 0.00194f 
C64544 _0786_/a_80_21# VGND 0.49142f 
C64545 _0456_ VGND 0.23635f
C64546 net234 VGND 0.27181f
C64547 _0855_/a_384_47# VGND 0.00329f 
C64548 _0855_/a_299_297# VGND 0.03893f 
C64549 _0855_/a_81_21# VGND 0.30156f 
C64550 _0464_ VGND 1.05948f
C64551 _0924_/a_27_47# VGND 0.30579f 
C64552 _1071_/a_1017_47# VGND 0.00404f 
C64553 _1071_/a_592_47# VGND 0.00677f 
C64554 _1071_/a_975_413# VGND 0 
C64555 _1071_/a_561_413# VGND 0 
C64556 _1071_/a_381_47# VGND 0.06186f 
C64557 _1071_/a_891_413# VGND 0.27622f 
C64558 _1071_/a_1059_315# VGND 0.39552f 
C64559 _1071_/a_466_413# VGND 0.21841f 
C64560 _1071_/a_634_159# VGND 0.25457f 
C64561 _1071_/a_193_47# VGND 0.35097f 
C64562 _1071_/a_27_47# VGND 0.5607f 
C64563 net81 VGND 0.53734f
C64564 acc0.A\[16\] VGND 1.54615f
C64565 _0607_/a_373_47# VGND 0.00399f 
C64566 _0607_/a_109_47# VGND 0.00827f 
C64567 _0607_/a_109_297# VGND 0.00551f 
C64568 _0607_/a_27_297# VGND 0.4506f 
C64569 _0143_ VGND 1.10298f
C64570 net21 VGND 0.58611f
C64571 net183 VGND 0.34507f
C64572 _0201_ VGND 0.54729f
C64573 _0538_/a_240_47# VGND 0.17453f 
C64574 _0538_/a_149_47# VGND 0.13313f 
C64575 _0538_/a_512_297# VGND 0 
C64576 _0538_/a_245_297# VGND 0 
C64577 _0538_/a_51_297# VGND 0.31925f 
C64578 net172 VGND 0.43937f
C64579 net124 VGND 0.63832f
C64580 _1038_/a_1017_47# VGND 0.00397f 
C64581 _1038_/a_592_47# VGND 0.00662f 
C64582 _1038_/a_975_413# VGND 0 
C64583 _1038_/a_381_47# VGND 0.06264f 
C64584 _1038_/a_891_413# VGND 0.27481f 
C64585 _1038_/a_1059_315# VGND 0.38391f 
C64586 _1038_/a_466_413# VGND 0.21185f 
C64587 _1038_/a_634_159# VGND 0.25198f 
C64588 _1038_/a_193_47# VGND 0.35971f 
C64589 _1038_/a_27_47# VGND 0.5669f 
C64590 net204 VGND 0.42005f
C64591 _0555_/a_240_47# VGND 0.16126f 
C64592 _0555_/a_149_47# VGND 0.125f 
C64593 _0555_/a_51_297# VGND 0.29165f 
C64594 _0624_/a_145_75# VGND 0.00763f 
C64595 _0624_/a_59_75# VGND 0.34464f 
C64596 _0432_ VGND 2.2712f
C64597 _0443_ VGND 0.40335f
C64598 net179 VGND 0.62547f
C64599 net141 VGND 0.59407f
C64600 _1055_/a_1017_47# VGND 0.00475f 
C64601 _1055_/a_592_47# VGND 0.0077f 
C64602 _1055_/a_975_413# VGND 0 
C64603 _1055_/a_561_413# VGND 0 
C64604 _1055_/a_381_47# VGND 0.06657f 
C64605 _1055_/a_891_413# VGND 0.29676f 
C64606 _1055_/a_1059_315# VGND 0.41413f 
C64607 _1055_/a_466_413# VGND 0.22195f 
C64608 _1055_/a_634_159# VGND 0.26391f 
C64609 _1055_/a_193_47# VGND 0.421f 
C64610 _1055_/a_27_47# VGND 0.62987f 
C64611 _0124_ VGND 0.43577f
C64612 _0216_ VGND 7.27173f
C64613 net155 VGND 1.19163f
C64614 _0195_ VGND 3.97286f
C64615 net210 VGND 0.3598f
C64616 _0572_/a_373_47# VGND 0.00313f 
C64617 _0572_/a_109_47# VGND 0.00862f 
C64618 _0572_/a_109_297# VGND 0.00788f 
C64619 _0572_/a_27_297# VGND 0.46107f 
C64620 _0641_/a_113_47# VGND 0.00199f 
C64621 _0342_ VGND 0.4425f
C64622 _0340_ VGND 0.75353f
C64623 _0341_ VGND 0.68099f
C64624 _0710_/a_381_47# VGND 0 
C64625 _0710_/a_109_47# VGND 0.00519f 
C64626 _0710_/a_109_297# VGND 0.00408f 
C64627 net186 VGND 0.45162f
C64628 hold39/a_391_47# VGND 0.26023f 
C64629 hold39/a_285_47# VGND 0.40763f 
C64630 hold39/a_49_47# VGND 0.45266f 
C64631 hold28/a_391_47# VGND 0.23969f 
C64632 hold28/a_285_47# VGND 0.39863f 
C64633 hold28/a_49_47# VGND 0.4697f 
C64634 control0.count\[2\] VGND 1.75255f
C64635 hold17/a_391_47# VGND 0.26764f 
C64636 hold17/a_285_47# VGND 0.45879f 
C64637 hold17/a_49_47# VGND 0.53069f 
C64638 _0856_/a_510_47# VGND 0.00832f 
C64639 _0856_/a_215_47# VGND 0.23328f 
C64640 _0856_/a_297_297# VGND 0 
C64641 _0856_/a_79_21# VGND 0.36471f 
C64642 _0787_/a_303_47# VGND 0.0063f 
C64643 _0787_/a_209_47# VGND 0.00666f 
C64644 _0787_/a_209_297# VGND 0.01024f 
C64645 _0787_/a_80_21# VGND 0.42091f 
C64646 _1072_/a_1017_47# VGND 0.00447f 
C64647 _1072_/a_592_47# VGND 0.00748f 
C64648 _1072_/a_975_413# VGND 0 
C64649 _1072_/a_381_47# VGND 0.06831f 
C64650 _1072_/a_891_413# VGND 0.2951f 
C64651 _1072_/a_1059_315# VGND 0.41687f 
C64652 _1072_/a_466_413# VGND 0.22266f 
C64653 _1072_/a_634_159# VGND 0.26919f 
C64654 _1072_/a_193_47# VGND 0.46656f 
C64655 _1072_/a_27_47# VGND 0.5759f 
C64656 clknet_1_0__leaf__0465_ VGND 5.83354f
C64657 _0539_/a_150_297# VGND 0 
C64658 _0539_/a_68_297# VGND 0.28134f 
C64659 _0239_ VGND 0.19797f
C64660 _0608_/a_27_47# VGND 0.175f 
C64661 _0608_/a_109_297# VGND 0 
C64662 net125 VGND 0.43989f
C64663 _1039_/a_1017_47# VGND 0.00429f 
C64664 _1039_/a_592_47# VGND 0.00691f 
C64665 _1039_/a_975_413# VGND 0 
C64666 _1039_/a_561_413# VGND 0 
C64667 _1039_/a_381_47# VGND 0.06191f 
C64668 _1039_/a_891_413# VGND 0.28651f 
C64669 _1039_/a_1059_315# VGND 0.39561f 
C64670 _1039_/a_466_413# VGND 0.22393f 
C64671 _1039_/a_634_159# VGND 0.27384f 
C64672 _1039_/a_193_47# VGND 0.37569f 
C64673 _1039_/a_27_47# VGND 0.58787f 
C64674 _0211_ VGND 0.66875f
C64675 _0556_/a_150_297# VGND 0 
C64676 _0556_/a_68_297# VGND 0.26547f 
C64677 _0625_/a_145_75# VGND 0.00731f 
C64678 _0625_/a_59_75# VGND 0.3092f 
C64679 pp[12] VGND 0.75564f
C64680 output39/a_27_47# VGND 0.44167f 
C64681 net182 VGND 0.38684f
C64682 _1056_/a_1017_47# VGND 0.00425f 
C64683 _1056_/a_592_47# VGND 0.00832f 
C64684 _1056_/a_975_413# VGND 0 
C64685 _1056_/a_561_413# VGND 0 
C64686 _1056_/a_381_47# VGND 0.08598f 
C64687 _1056_/a_891_413# VGND 0.2818f 
C64688 _1056_/a_1059_315# VGND 0.39201f 
C64689 _1056_/a_466_413# VGND 0.23345f 
C64690 _1056_/a_634_159# VGND 0.26582f 
C64691 _1056_/a_193_47# VGND 0.39053f 
C64692 _1056_/a_27_47# VGND 0.62991f 
C64693 net108 VGND 0.31855f
C64694 clknet_1_0__leaf__0462_ VGND 5.07795f
C64695 _0573_/a_27_47# VGND 0.70368f 
C64696 _0273_ VGND 0.44636f
C64697 _0642_/a_382_47# VGND 0.00386f 
C64698 _0642_/a_298_297# VGND 0.00684f 
C64699 _0642_/a_215_297# VGND 0.41064f 
C64700 _0642_/a_27_413# VGND 0.26869f 
C64701 hold49/a_391_47# VGND 0.23647f 
C64702 hold49/a_285_47# VGND 0.3943f 
C64703 hold49/a_49_47# VGND 0.43434f 
C64704 hold38/a_391_47# VGND 0.26043f 
C64705 hold38/a_285_47# VGND 0.41214f 
C64706 hold38/a_49_47# VGND 0.46072f 
C64707 hold27/a_391_47# VGND 0.25713f 
C64708 hold27/a_285_47# VGND 0.42026f 
C64709 hold27/a_49_47# VGND 0.4869f 
C64710 net163 VGND 0.34029f
C64711 _0129_ VGND 0.29929f
C64712 hold16/a_391_47# VGND 0.2422f 
C64713 hold16/a_285_47# VGND 0.39879f 
C64714 hold16/a_49_47# VGND 0.44076f 
C64715 _0403_ VGND 0.61927f
C64716 _0788_/a_150_297# VGND 0 
C64717 _0788_/a_68_297# VGND 0.28251f 
C64718 _0457_ VGND 1.67165f
C64719 _0857_/a_27_47# VGND 0.36593f 
C64720 _0222_ VGND 1.91479f
C64721 _0590_/a_113_47# VGND 0.00202f 
C64722 clkload4/Y VGND 0.20088f
C64723 clkload4/a_268_47# VGND 0.008f 
C64724 clkload4/a_110_47# VGND 0.00176f 
C64725 _0461_ VGND 1.47382f
C64726 _0891_/a_27_47# VGND 0.30796f 
C64727 _0478_ VGND 0.609f
C64728 _0960_/a_181_47# VGND 0.00227f 
C64729 _0960_/a_109_47# VGND 0 
C64730 _0960_/a_27_47# VGND 0.2977f 
C64731 _0241_ VGND 0.71266f
C64732 net248 VGND 0.61823f
C64733 hold101/a_391_47# VGND 0.28979f 
C64734 hold101/a_285_47# VGND 0.44236f 
C64735 hold101/a_49_47# VGND 0.45419f 
C64736 _0258_ VGND 0.704f
C64737 _0257_ VGND 0.84676f
C64738 _0626_/a_150_297# VGND 0 
C64739 _0626_/a_68_297# VGND 0.27006f 
C64740 _0134_ VGND 0.30887f
C64741 _0557_/a_240_47# VGND 0.16146f 
C64742 _0557_/a_149_47# VGND 0.12557f 
C64743 _0557_/a_512_297# VGND 0 
C64744 _0557_/a_245_297# VGND 0 
C64745 _0557_/a_51_297# VGND 0.27646f 
C64746 clk VGND 3.26277f
C64747 clkbuf_0_clk/a_110_47# VGND 2.28072f 
C64748 pp[11] VGND 0.97513f
C64749 output38/a_27_47# VGND 0.42145f 
C64750 pp[21] VGND 1.07843f
C64751 net49 VGND 1.35221f
C64752 output49/a_27_47# VGND 0.45649f 
C64753 net189 VGND 0.35659f
C64754 _1057_/a_1017_47# VGND 0.00414f 
C64755 _1057_/a_592_47# VGND 0.00689f 
C64756 _1057_/a_975_413# VGND 0 
C64757 _1057_/a_561_413# VGND 0 
C64758 _1057_/a_381_47# VGND 0.06388f 
C64759 _1057_/a_891_413# VGND 0.30291f 
C64760 _1057_/a_1059_315# VGND 0.42895f 
C64761 _1057_/a_466_413# VGND 0.23635f 
C64762 _1057_/a_634_159# VGND 0.27199f 
C64763 _1057_/a_193_47# VGND 0.38791f 
C64764 _1057_/a_27_47# VGND 0.6241f 
C64765 _0574_/a_373_47# VGND 0.00344f 
C64766 _0574_/a_109_47# VGND 0.00792f 
C64767 _0574_/a_109_297# VGND 0.00274f 
C64768 _0574_/a_27_297# VGND 0.45278f 
C64769 _0344_ VGND 0.26001f
C64770 _0712_/a_561_47# VGND 0.00684f 
C64771 _0712_/a_465_47# VGND 0.00452f 
C64772 _0712_/a_381_47# VGND 0.00243f 
C64773 _0712_/a_297_297# VGND 0.04669f 
C64774 _0712_/a_79_21# VGND 0.28506f 
C64775 _0275_ VGND 0.68241f
C64776 _0274_ VGND 0.64645f
C64777 _0272_ VGND 0.1744f
C64778 _0643_/a_253_47# VGND 0.20955f 
C64779 _0643_/a_337_297# VGND 0 
C64780 _0643_/a_253_297# VGND 0 
C64781 _0643_/a_103_199# VGND 0.31224f 
C64782 hold59/a_391_47# VGND 0.24008f 
C64783 hold59/a_285_47# VGND 0.39644f 
C64784 hold59/a_49_47# VGND 0.46434f 
C64785 hold48/a_391_47# VGND 0.26886f 
C64786 hold48/a_285_47# VGND 0.44804f 
C64787 hold48/a_49_47# VGND 0.51027f 
C64788 hold37/a_391_47# VGND 0.25911f 
C64789 hold37/a_285_47# VGND 0.42633f 
C64790 hold37/a_49_47# VGND 0.4625f 
C64791 hold26/a_391_47# VGND 0.25969f 
C64792 hold26/a_285_47# VGND 0.42662f 
C64793 hold26/a_49_47# VGND 0.49418f 
C64794 net162 VGND 0.47033f
C64795 acc0.A\[31\] VGND 1.37294f
C64796 hold15/a_391_47# VGND 0.26253f 
C64797 hold15/a_285_47# VGND 0.42408f 
C64798 hold15/a_49_47# VGND 0.47482f 
C64799 _0458_ VGND 1.4954f
C64800 _0858_/a_27_47# VGND 0.36449f 
C64801 _0299_ VGND 0.73341f
C64802 _0298_ VGND 1.09531f
C64803 _0404_ VGND 1.50589f
C64804 _0789_/a_315_47# VGND 0 
C64805 _0789_/a_208_47# VGND 0.00254f 
C64806 _0789_/a_544_297# VGND 0.00152f 
C64807 _0789_/a_201_297# VGND 0.00894f 
C64808 _0789_/a_75_199# VGND 0.56116f 
C64809 _0591_/a_109_297# VGND 0 
C64810 _0660_/a_113_47# VGND 0.00271f 
C64811 clkload3/Y VGND 0.20457f
C64812 clkload3/a_268_47# VGND 0.00802f 
C64813 clkload3/a_110_47# VGND 0.00176f 
C64814 net123 VGND 0.69521f
C64815 clknet_1_0__leaf__0463_ VGND 5.31876f
C64816 _0479_ VGND 0.27744f
C64817 _0961_/a_199_47# VGND 0.00396f 
C64818 _0961_/a_113_297# VGND 0.04031f 
C64819 acc0.A\[14\] VGND 4.26862f
C64820 hold100/a_391_47# VGND 0.24805f 
C64821 hold100/a_285_47# VGND 0.4077f 
C64822 hold100/a_49_47# VGND 0.44049f 
C64823 _0212_ VGND 0.46387f
C64824 net185 VGND 1.0641f
C64825 _0558_/a_150_297# VGND 0 
C64826 _0558_/a_68_297# VGND 0.28598f 
C64827 _0627_/a_109_93# VGND 0.23879f 
C64828 _0627_/a_215_53# VGND 0.39213f 
C64829 pp[10] VGND 0.78082f
C64830 output37/a_27_47# VGND 0.69272f 
C64831 pp[20] VGND 0.95933f
C64832 net48 VGND 2.02472f
C64833 output48/a_27_47# VGND 0.48176f 
C64834 pp[30] VGND 0.78583f
C64835 net59 VGND 1.06036f
C64836 output59/a_27_47# VGND 0.42713f 
C64837 net144 VGND 0.59679f
C64838 _1058_/a_1017_47# VGND 0.00422f 
C64839 _1058_/a_592_47# VGND 0.00684f 
C64840 _1058_/a_975_413# VGND 0 
C64841 _1058_/a_561_413# VGND 0 
C64842 _1058_/a_381_47# VGND 0.0621f 
C64843 _1058_/a_891_413# VGND 0.27825f 
C64844 _1058_/a_1059_315# VGND 0.38799f 
C64845 _1058_/a_466_413# VGND 0.21311f 
C64846 _1058_/a_634_159# VGND 0.2552f 
C64847 _1058_/a_193_47# VGND 0.35198f 
C64848 _1058_/a_27_47# VGND 0.56754f 
C64849 net199 VGND 0.60788f
C64850 _0575_/a_373_47# VGND 0.00236f 
C64851 _0575_/a_109_47# VGND 0.00756f 
C64852 _0575_/a_109_297# VGND 0.00277f 
C64853 _0575_/a_27_297# VGND 0.43018f 
C64854 _0276_ VGND 0.64554f
C64855 _0644_/a_285_47# VGND 0.22969f 
C64856 _0644_/a_129_47# VGND 0.00587f 
C64857 _0644_/a_377_297# VGND 0 
C64858 _0644_/a_47_47# VGND 0.31551f 
C64859 _0713_/a_27_47# VGND 0.7553f 
C64860 net117 VGND 0.31742f
C64861 hold69/a_391_47# VGND 0.2362f 
C64862 hold69/a_285_47# VGND 0.3927f 
C64863 hold69/a_49_47# VGND 0.43299f 
C64864 net205 VGND 0.27462f
C64865 hold58/a_391_47# VGND 0.25758f 
C64866 hold58/a_285_47# VGND 0.41608f 
C64867 hold58/a_49_47# VGND 0.44442f 
C64868 net194 VGND 0.47199f
C64869 hold47/a_391_47# VGND 0.25504f 
C64870 hold47/a_285_47# VGND 0.41565f 
C64871 hold47/a_49_47# VGND 0.47868f 
C64872 hold36/a_391_47# VGND 0.24054f 
C64873 hold36/a_285_47# VGND 0.39652f 
C64874 hold36/a_49_47# VGND 0.46528f 
C64875 hold25/a_391_47# VGND 0.24507f 
C64876 hold25/a_285_47# VGND 0.40383f 
C64877 hold25/a_49_47# VGND 0.43876f 
C64878 hold14/a_391_47# VGND 0.25843f 
C64879 hold14/a_285_47# VGND 0.41424f 
C64880 hold14/a_49_47# VGND 0.44494f 
C64881 _0592_/a_150_297# VGND 0 
C64882 _0592_/a_68_297# VGND 0.28374f 
C64883 _0108_ VGND 0.36544f
C64884 _0358_ VGND 0.22484f
C64885 _0357_ VGND 0.93891f
C64886 _0730_/a_510_47# VGND 0.0058f 
C64887 _0730_/a_215_47# VGND 0.21837f 
C64888 _0730_/a_79_21# VGND 0.32721f 
C64889 _0293_ VGND 0.44807f
C64890 _0287_ VGND 0.56432f
C64891 _0289_ VGND 1.15814f
C64892 _0292_ VGND 1.36993f
C64893 _0661_/a_277_297# VGND 0 
C64894 _0661_/a_205_297# VGND 0 
C64895 _0661_/a_109_297# VGND 0 
C64896 _0661_/a_27_297# VGND 0.40159f 
C64897 clkload2/Y VGND 0.20674f
C64898 clkload2/a_268_47# VGND 0.00821f 
C64899 clkload2/a_110_47# VGND 0.00196f 
C64900 _0962_/a_109_297# VGND 0.00109f 
C64901 clknet_1_1__leaf__0459_ VGND 5.88592f
C64902 _0559_/a_240_47# VGND 0.17319f 
C64903 _0559_/a_149_47# VGND 0.12982f 
C64904 _0559_/a_512_297# VGND 0 
C64905 _0559_/a_245_297# VGND 0 
C64906 _0559_/a_51_297# VGND 0.2761f 
C64907 _0260_ VGND 1.01195f
C64908 _0628_/a_109_297# VGND 0.0051f 
C64909 pp[1] VGND 0.63149f
C64910 output47/a_27_47# VGND 0.72077f 
C64911 pp[2] VGND 0.64598f
C64912 output58/a_27_47# VGND 0.74047f 
C64913 pp[0] VGND 0.4746f
C64914 net36 VGND 3.62455f
C64915 output36/a_27_47# VGND 0.41674f 
C64916 _0157_ VGND 0.44392f
C64917 net145 VGND 0.76088f
C64918 _1059_/a_1017_47# VGND 0.00506f 
C64919 _1059_/a_592_47# VGND 0.00785f 
C64920 _1059_/a_975_413# VGND 0 
C64921 _1059_/a_561_413# VGND 0 
C64922 _1059_/a_381_47# VGND 0.06637f 
C64923 _1059_/a_891_413# VGND 0.29801f 
C64924 _1059_/a_1059_315# VGND 0.41012f 
C64925 _1059_/a_466_413# VGND 0.21761f 
C64926 _1059_/a_634_159# VGND 0.27536f 
C64927 _1059_/a_193_47# VGND 0.37935f 
C64928 _1059_/a_27_47# VGND 0.61769f 
C64929 _0576_/a_373_47# VGND 0.00344f 
C64930 _0576_/a_109_47# VGND 0.00806f 
C64931 _0576_/a_109_297# VGND 0.00298f 
C64932 _0576_/a_27_297# VGND 0.44222f 
C64933 _0645_/a_285_47# VGND 0.22763f 
C64934 _0645_/a_129_47# VGND 0.00554f 
C64935 _0645_/a_377_297# VGND 0 
C64936 _0645_/a_47_47# VGND 0.32635f 
C64937 _0111_ VGND 0.71867f
C64938 net225 VGND 0.26707f
C64939 _0714_/a_240_47# VGND 0.18015f 
C64940 _0714_/a_149_47# VGND 0.1454f 
C64941 _0714_/a_512_297# VGND 0 
C64942 _0714_/a_245_297# VGND 0.00232f 
C64943 _0714_/a_51_297# VGND 0.30976f 
C64944 net226 VGND 0.4392f
C64945 hold79/a_391_47# VGND 0.25911f 
C64946 hold79/a_285_47# VGND 0.42331f 
C64947 hold79/a_49_47# VGND 0.48764f 
C64948 net215 VGND 0.24528f
C64949 hold68/a_391_47# VGND 0.2456f 
C64950 hold68/a_285_47# VGND 0.40486f 
C64951 hold68/a_49_47# VGND 0.43857f 
C64952 hold57/a_391_47# VGND 0.24912f 
C64953 hold57/a_285_47# VGND 0.40963f 
C64954 hold57/a_49_47# VGND 0.53479f 
C64955 net193 VGND 0.5104f
C64956 comp0.B\[13\] VGND 1.19251f
C64957 hold46/a_391_47# VGND 0.23868f 
C64958 hold46/a_285_47# VGND 0.40425f 
C64959 hold46/a_49_47# VGND 0.46284f 
C64960 _0154_ VGND 0.20545f
C64961 hold35/a_391_47# VGND 0.30523f 
C64962 hold35/a_285_47# VGND 0.447f 
C64963 hold35/a_49_47# VGND 0.45656f 
C64964 comp0.B\[7\] VGND 0.70619f
C64965 hold24/a_391_47# VGND 0.23505f 
C64966 hold24/a_285_47# VGND 0.39339f 
C64967 hold24/a_49_47# VGND 0.4617f 
C64968 hold13/a_391_47# VGND 0.28288f 
C64969 hold13/a_285_47# VGND 0.49179f 
C64970 hold13/a_49_47# VGND 0.47196f 
C64971 _0259_ VGND 1.31421f
C64972 _0662_/a_384_47# VGND 0.00328f 
C64973 _0662_/a_299_297# VGND 0.03806f 
C64974 _0662_/a_81_21# VGND 0.30014f 
C64975 _0225_ VGND 1.29712f
C64976 _0224_ VGND 0.31786f
C64977 _0593_/a_113_47# VGND 0.00192f 
C64978 _0731_/a_384_47# VGND 0.00357f 
C64979 _0731_/a_299_297# VGND 0.0382f 
C64980 _0731_/a_81_21# VGND 0.33466f 
C64981 _0093_ VGND 0.35407f
C64982 _0413_ VGND 0.28155f
C64983 _0412_ VGND 0.18647f
C64984 _0800_/a_240_47# VGND 0.18047f 
C64985 _0800_/a_149_47# VGND 0.13269f 
C64986 _0800_/a_512_297# VGND 0.00235f 
C64987 _0800_/a_245_297# VGND 0 
C64988 _0800_/a_51_297# VGND 0.33296f 
C64989 clkload1/Y VGND 0.21918f
C64990 clkload1/a_268_47# VGND 0.00846f 
C64991 clkload1/a_110_47# VGND 0.00187f 
C64992 _0946_/a_184_297# VGND 0 
C64993 _0946_/a_112_297# VGND 0 
C64994 _0946_/a_30_53# VGND 0.49711f 
C64995 _0481_ VGND 1.10112f
C64996 _0963_/a_285_47# VGND 0.00552f 
C64997 _0963_/a_285_297# VGND 0.00138f 
C64998 _0963_/a_117_297# VGND 0 
C64999 _0963_/a_35_297# VGND 0.42738f 
C65000 net58 VGND 2.20971f
C65001 acc0.A\[2\] VGND 0.87555f
C65002 _0629_/a_145_75# VGND 0.00359f 
C65003 _0629_/a_59_75# VGND 0.30473f 
C65004 _0179_ VGND 7.87854f
C65005 _0500_/a_27_47# VGND 0.66714f 
C65006 done VGND 1.28379f
C65007 net35 VGND 1.5436f
C65008 output35/a_27_47# VGND 0.48119f 
C65009 pp[19] VGND 0.87087f
C65010 net46 VGND 2.08886f
C65011 output46/a_27_47# VGND 0.44846f 
C65012 pp[29] VGND 0.82574f
C65013 output57/a_27_47# VGND 0.48285f 
C65014 _0646_/a_285_47# VGND 0.23002f 
C65015 _0646_/a_129_47# VGND 0.00608f 
C65016 _0646_/a_377_297# VGND 0 
C65017 _0646_/a_47_47# VGND 0.31851f 
C65018 _0120_ VGND 0.21954f
C65019 _0183_ VGND 4.07066f
C65020 acc0.A\[22\] VGND 0.76476f
C65021 _0217_ VGND 4.77978f
C65022 net150 VGND 1.07627f
C65023 _0577_/a_373_47# VGND 0.00328f 
C65024 _0577_/a_109_47# VGND 0.00768f 
C65025 _0577_/a_109_297# VGND 0.00376f 
C65026 _0577_/a_27_297# VGND 0.44259f 
C65027 _0715_/a_27_47# VGND 0.68771f 
C65028 net45 VGND 2.22653f
C65029 _0098_ VGND 0.34652f
C65030 net86 VGND 0.6128f
C65031 _1000_/a_1017_47# VGND 0.00407f 
C65032 _1000_/a_592_47# VGND 0.00703f 
C65033 _1000_/a_975_413# VGND 0 
C65034 _1000_/a_561_413# VGND 0 
C65035 _1000_/a_381_47# VGND 0.06191f 
C65036 _1000_/a_891_413# VGND 0.28073f 
C65037 _1000_/a_1059_315# VGND 0.4014f 
C65038 _1000_/a_466_413# VGND 0.21433f 
C65039 _1000_/a_634_159# VGND 0.256f 
C65040 _1000_/a_193_47# VGND 0.35148f 
C65041 _1000_/a_27_47# VGND 0.59444f 
C65042 hold89/a_391_47# VGND 0.24479f 
C65043 hold89/a_285_47# VGND 0.40323f 
C65044 hold89/a_49_47# VGND 0.44685f 
C65045 hold78/a_391_47# VGND 0.26859f 
C65046 hold78/a_285_47# VGND 0.42868f 
C65047 hold78/a_49_47# VGND 0.4682f 
C65048 hold67/a_391_47# VGND 0.29208f 
C65049 hold67/a_285_47# VGND 0.46085f 
C65050 hold67/a_49_47# VGND 0.52664f 
C65051 net203 VGND 0.46596f
C65052 hold56/a_391_47# VGND 0.26269f 
C65053 hold56/a_285_47# VGND 0.4377f 
C65054 hold56/a_49_47# VGND 0.49582f 
C65055 hold45/a_391_47# VGND 0.24804f 
C65056 hold45/a_285_47# VGND 0.41692f 
C65057 hold45/a_49_47# VGND 0.49621f 
C65058 hold34/a_391_47# VGND 0.26188f 
C65059 hold34/a_285_47# VGND 0.42747f 
C65060 hold34/a_49_47# VGND 0.45779f 
C65061 hold23/a_391_47# VGND 0.24714f 
C65062 hold23/a_285_47# VGND 0.40927f 
C65063 hold23/a_49_47# VGND 0.44094f 
C65064 hold12/a_391_47# VGND 0.28113f 
C65065 hold12/a_285_47# VGND 0.46039f 
C65066 hold12/a_49_47# VGND 0.50646f 
C65067 net126 VGND 0.35673f
C65068 acc0.A\[20\] VGND 1.40631f
C65069 _0594_/a_113_47# VGND 0.00194f 
C65070 _0732_/a_303_47# VGND 0.00651f 
C65071 _0732_/a_209_47# VGND 0.00701f 
C65072 _0732_/a_209_297# VGND 0.00804f 
C65073 _0732_/a_80_21# VGND 0.43077f 
C65074 _0663_/a_297_47# VGND 0.00423f 
C65075 _0663_/a_207_413# VGND 0.26529f 
C65076 _0663_/a_27_413# VGND 0.28749f 
C65077 _0414_ VGND 0.28592f
C65078 _0801_/a_113_47# VGND 0.00226f 
C65079 clkload0/X VGND 0.31257f
C65080 clkload0/a_27_47# VGND 0.76255f 
C65081 _0467_ VGND 1.17179f
C65082 _0947_/a_109_297# VGND 0 
C65083 net78 VGND 0.58596f
C65084 _0311_ VGND 0.56951f
C65085 _0305_ VGND 2.3739f
C65086 _0680_/a_300_47# VGND 0.00418f 
C65087 _0680_/a_217_297# VGND 0.00355f 
C65088 _0680_/a_80_21# VGND 0.5379f 
C65089 _0482_ VGND 0.30394f
C65090 _0964_/a_109_297# VGND 0.00118f 
C65091 _0170_ VGND 0.35199f
C65092 net167 VGND 0.96109f
C65093 _0490_ VGND 0.30743f
C65094 _0981_/a_373_47# VGND 0.00245f 
C65095 _0981_/a_109_47# VGND 0.00748f 
C65096 _0981_/a_109_297# VGND 0.006f 
C65097 _0981_/a_27_297# VGND 0.43467f 
C65098 _0501_/a_27_47# VGND 0.40272f 
C65099 pp[9] VGND 0.43888f
C65100 output67/a_27_47# VGND 0.66769f 
C65101 pp[18] VGND 0.66663f
C65102 output45/a_27_47# VGND 0.45433f 
C65103 pp[28] VGND 0.53195f
C65104 output56/a_27_47# VGND 0.42838f 
C65105 _0647_/a_285_47# VGND 0.22263f 
C65106 _0647_/a_129_47# VGND 0.00518f 
C65107 _0647_/a_377_297# VGND 0 
C65108 _0647_/a_47_47# VGND 0.32228f 
C65109 net187 VGND 0.9393f
C65110 _0578_/a_373_47# VGND 0.00344f 
C65111 _0578_/a_109_47# VGND 0.00806f 
C65112 _0578_/a_109_297# VGND 0.00275f 
C65113 _0578_/a_27_297# VGND 0.44311f 
C65114 _0716_/a_27_47# VGND 0.72254f 
C65115 _1001_/a_1017_47# VGND 0.00417f 
C65116 _1001_/a_592_47# VGND 0.00816f 
C65117 _1001_/a_975_413# VGND 0 
C65118 _1001_/a_561_413# VGND 0 
C65119 _1001_/a_381_47# VGND 0.06808f 
C65120 _1001_/a_891_413# VGND 0.28444f 
C65121 _1001_/a_1059_315# VGND 0.38996f 
C65122 _1001_/a_466_413# VGND 0.22555f 
C65123 _1001_/a_634_159# VGND 0.27325f 
C65124 _1001_/a_193_47# VGND 0.4043f 
C65125 _1001_/a_27_47# VGND 0.58484f 
C65126 hold99/a_391_47# VGND 0.27654f 
C65127 hold99/a_285_47# VGND 0.46575f 
C65128 hold99/a_49_47# VGND 0.48922f 
C65129 hold88/a_391_47# VGND 0.26432f 
C65130 hold88/a_285_47# VGND 0.42509f 
C65131 hold88/a_49_47# VGND 0.50336f 
C65132 hold77/a_391_47# VGND 0.27232f 
C65133 hold77/a_285_47# VGND 0.46173f 
C65134 hold77/a_49_47# VGND 0.52959f 
C65135 net213 VGND 0.26899f
C65136 hold66/a_391_47# VGND 0.24137f 
C65137 hold66/a_285_47# VGND 0.39339f 
C65138 hold66/a_49_47# VGND 0.43602f 
C65139 _0130_ VGND 0.33359f
C65140 hold55/a_391_47# VGND 0.24199f 
C65141 hold55/a_285_47# VGND 0.39915f 
C65142 hold55/a_49_47# VGND 0.46934f 
C65143 hold44/a_391_47# VGND 0.27853f 
C65144 hold44/a_285_47# VGND 0.46598f 
C65145 hold44/a_49_47# VGND 0.52243f 
C65146 hold33/a_391_47# VGND 0.25775f 
C65147 hold33/a_285_47# VGND 0.43839f 
C65148 hold33/a_49_47# VGND 0.45345f 
C65149 hold22/a_391_47# VGND 0.23877f 
C65150 hold22/a_285_47# VGND 0.39596f 
C65151 hold22/a_49_47# VGND 0.43146f 
C65152 net158 VGND 0.29779f
C65153 hold11/a_391_47# VGND 0.26137f 
C65154 hold11/a_285_47# VGND 0.4263f 
C65155 hold11/a_49_47# VGND 0.50905f 
C65156 _0227_ VGND 1.83481f
C65157 acc0.A\[21\] VGND 1.18188f
C65158 _0595_/a_109_297# VGND 0 
C65159 _0361_ VGND 0.63378f
C65160 _0733_/a_448_47# VGND 0.23174f 
C65161 _0733_/a_544_297# VGND 0.0014f 
C65162 _0733_/a_222_93# VGND 0.22735f 
C65163 _0733_/a_79_199# VGND 0.2272f 
C65164 _0284_ VGND 0.90451f
C65165 _0285_ VGND 0.61004f
C65166 _0664_/a_297_47# VGND 0.15308f 
C65167 _0664_/a_79_21# VGND 0.2685f 
C65168 _0802_/a_145_75# VGND 0.00361f 
C65169 _0802_/a_59_75# VGND 0.3061f 
C65170 _0948_/a_109_297# VGND 0.0022f 
C65171 _0750_/a_181_47# VGND 0.00243f 
C65172 _0750_/a_109_47# VGND 0.00158f 
C65173 _0750_/a_27_47# VGND 0.33039f 
C65174 _0681_/a_113_47# VGND 0.00207f 
C65175 _0483_ VGND 0.45049f
C65176 control0.count\[3\] VGND 0.70142f
C65177 _0965_/a_285_47# VGND 0.21554f 
C65178 _0965_/a_129_47# VGND 0.00382f 
C65179 _0965_/a_377_297# VGND 0 
C65180 _0965_/a_47_47# VGND 0.29774f 
C65181 _0080_ VGND 0.3906f
C65182 net68 VGND 0.56921f
C65183 _0982_/a_1017_47# VGND 0.0042f 
C65184 _0982_/a_592_47# VGND 0.00689f 
C65185 _0982_/a_975_413# VGND 0 
C65186 _0982_/a_561_413# VGND 0 
C65187 _0982_/a_381_47# VGND 0.06243f 
C65188 _0982_/a_891_413# VGND 0.27882f 
C65189 _0982_/a_1059_315# VGND 0.38735f 
C65190 _0982_/a_466_413# VGND 0.21528f 
C65191 _0982_/a_634_159# VGND 0.25556f 
C65192 _0982_/a_193_47# VGND 0.36807f 
C65193 _0982_/a_27_47# VGND 0.61389f 
C65194 clknet_1_1__leaf__0460_ VGND 4.91902f
C65195 _0502_/a_27_47# VGND 0.67073f 
C65196 clknet_1_0__leaf__0458_ VGND 3.77418f
C65197 pp[8] VGND 0.43331f
C65198 output66/a_27_47# VGND 0.69582f 
C65199 pp[17] VGND 0.97972f
C65200 net44 VGND 2.08295f
C65201 output44/a_27_47# VGND 0.41823f 
C65202 pp[27] VGND 0.54895f
C65203 output55/a_27_47# VGND 0.3945f 
C65204 net211 VGND 0.49948f
C65205 _0579_/a_373_47# VGND 0.0029f 
C65206 _0579_/a_109_47# VGND 0.00869f 
C65207 _0579_/a_109_297# VGND 0.01611f 
C65208 _0579_/a_27_297# VGND 0.4547f 
C65209 _0348_ VGND 0.30057f
C65210 _0717_/a_303_47# VGND 0.00609f 
C65211 _0717_/a_209_47# VGND 0.00568f 
C65212 _0717_/a_209_297# VGND 0.00737f 
C65213 _0717_/a_80_21# VGND 0.42241f 
C65214 _0280_ VGND 0.65297f
C65215 _0278_ VGND 0.65802f
C65216 _0279_ VGND 0.97297f
C65217 _0648_/a_277_297# VGND 0 
C65218 _0648_/a_205_297# VGND 0 
C65219 _0648_/a_109_297# VGND 0 
C65220 _0648_/a_27_297# VGND 0.39659f 
C65221 _0100_ VGND 0.46488f
C65222 net88 VGND 0.50663f
C65223 _1002_/a_1017_47# VGND 0.00447f 
C65224 _1002_/a_592_47# VGND 0.00748f 
C65225 _1002_/a_381_47# VGND 0.06744f 
C65226 _1002_/a_891_413# VGND 0.29021f 
C65227 _1002_/a_1059_315# VGND 0.40825f 
C65228 _1002_/a_466_413# VGND 0.23811f 
C65229 _1002_/a_634_159# VGND 0.28161f 
C65230 _1002_/a_193_47# VGND 0.38245f 
C65231 _1002_/a_27_47# VGND 0.5947f 
C65232 net245 VGND 0.99985f
C65233 net40 VGND 2.32604f
C65234 hold98/a_391_47# VGND 0.26072f 
C65235 hold98/a_285_47# VGND 0.42731f 
C65236 hold98/a_49_47# VGND 0.48792f 
C65237 hold87/a_391_47# VGND 0.24475f 
C65238 hold87/a_285_47# VGND 0.40431f 
C65239 hold87/a_49_47# VGND 0.44166f 
C65240 hold76/a_391_47# VGND 0.25793f 
C65241 hold76/a_285_47# VGND 0.41473f 
C65242 hold76/a_49_47# VGND 0.45263f 
C65243 hold65/a_391_47# VGND 0.25879f 
C65244 hold65/a_285_47# VGND 0.42684f 
C65245 hold65/a_49_47# VGND 0.45045f 
C65246 hold54/a_391_47# VGND 0.25367f 
C65247 hold54/a_285_47# VGND 0.4567f 
C65248 hold54/a_49_47# VGND 0.48752f 
C65249 hold43/a_391_47# VGND 0.27651f 
C65250 hold43/a_285_47# VGND 0.4719f 
C65251 hold43/a_49_47# VGND 0.56416f 
C65252 hold32/a_391_47# VGND 0.25564f 
C65253 hold32/a_285_47# VGND 0.41763f 
C65254 hold32/a_49_47# VGND 0.43666f 
C65255 hold21/a_391_47# VGND 0.25252f 
C65256 hold21/a_285_47# VGND 0.40976f 
C65257 hold21/a_49_47# VGND 0.46464f 
C65258 hold10/a_391_47# VGND 0.23796f 
C65259 hold10/a_285_47# VGND 0.39287f 
C65260 hold10/a_49_47# VGND 0.43075f 
C65261 _0596_/a_145_75# VGND 0.00376f 
C65262 _0596_/a_59_75# VGND 0.30508f 
C65263 _0362_ VGND 0.33684f
C65264 _0734_/a_285_47# VGND 0.23057f 
C65265 _0734_/a_129_47# VGND 0.00583f 
C65266 _0734_/a_377_297# VGND 0 
C65267 _0734_/a_47_47# VGND 0.36613f 
C65268 _0665_/a_109_297# VGND 0 
C65269 clknet_0__0457_ VGND 3.76362f
C65270 clkbuf_1_0__f__0457_/a_110_47# VGND 2.31019f 
C65271 _0803_/a_150_297# VGND 0 
C65272 _0803_/a_68_297# VGND 0.2676f 
C65273 _0469_ VGND 0.24553f
C65274 _0949_/a_145_75# VGND 0.00355f 
C65275 _0949_/a_59_75# VGND 0.27539f 
C65276 _0682_/a_150_297# VGND 0 
C65277 _0682_/a_68_297# VGND 0.28458f 
C65278 net214 VGND 0.43036f
C65279 _0820_/a_510_47# VGND 0.01135f 
C65280 _0820_/a_215_47# VGND 0.2302f 
C65281 _0820_/a_297_297# VGND 0.00648f 
C65282 _0820_/a_79_21# VGND 0.40376f 
C65283 _0751_/a_183_297# VGND 0 
C65284 _0751_/a_111_297# VGND 0 
C65285 _0751_/a_29_53# VGND 0.40176f 
C65286 net236 VGND 0.34798f
C65287 _0966_/a_27_47# VGND 0.18214f 
C65288 _0966_/a_109_297# VGND 0 
C65289 net69 VGND 0.3204f
C65290 _0983_/a_1017_47# VGND 0.00404f 
C65291 _0983_/a_592_47# VGND 0.00662f 
C65292 _0983_/a_381_47# VGND 0.06058f 
C65293 _0983_/a_891_413# VGND 0.29564f 
C65294 _0983_/a_1059_315# VGND 0.42461f 
C65295 _0983_/a_466_413# VGND 0.2296f 
C65296 _0983_/a_634_159# VGND 0.26703f 
C65297 _0983_/a_193_47# VGND 0.3727f 
C65298 _0983_/a_27_47# VGND 0.58643f 
C65299 pp[7] VGND 0.70653f
C65300 output65/a_27_47# VGND 0.7166f 
C65301 pp[16] VGND 0.74957f
C65302 output43/a_27_47# VGND 0.45302f 
C65303 pp[26] VGND 1.10533f
C65304 net54 VGND 1.3571f
C65305 output54/a_27_47# VGND 0.44458f 
C65306 _0649_/a_113_47# VGND 0.002f 
C65307 _0349_ VGND 1.56811f
C65308 _0337_ VGND 1.29909f
C65309 _0718_/a_285_47# VGND 0.23274f 
C65310 _0718_/a_129_47# VGND 0.0056f 
C65311 _0718_/a_377_297# VGND 0 
C65312 _0718_/a_47_47# VGND 0.304f 
C65313 _0101_ VGND 0.58632f
C65314 net89 VGND 0.69869f
C65315 _1003_/a_1017_47# VGND 0.00467f 
C65316 _1003_/a_592_47# VGND 0.00777f 
C65317 _1003_/a_975_413# VGND 0 
C65318 _1003_/a_561_413# VGND 0 
C65319 _1003_/a_381_47# VGND 0.07048f 
C65320 _1003_/a_891_413# VGND 0.29171f 
C65321 _1003_/a_1059_315# VGND 0.40075f 
C65322 _1003_/a_466_413# VGND 0.22819f 
C65323 _1003_/a_634_159# VGND 0.28198f 
C65324 _1003_/a_193_47# VGND 0.40137f 
C65325 _1003_/a_27_47# VGND 0.65168f 
C65326 net14 VGND 0.38823f
C65327 net168 VGND 1.51992f
C65328 _0520_/a_373_47# VGND 0.00395f 
C65329 _0520_/a_109_47# VGND 0.00627f 
C65330 _0520_/a_109_297# VGND 0.00735f 
C65331 _0520_/a_27_297# VGND 0.44421f 
C65332 hold97/a_391_47# VGND 0.25232f 
C65333 hold97/a_285_47# VGND 0.40287f 
C65334 hold97/a_49_47# VGND 0.47545f 
C65335 net233 VGND 0.44964f
C65336 net61 VGND 1.8036f
C65337 hold86/a_391_47# VGND 0.24074f 
C65338 hold86/a_285_47# VGND 0.40371f 
C65339 hold86/a_49_47# VGND 0.43812f 
C65340 hold75/a_391_47# VGND 0.25423f 
C65341 hold75/a_285_47# VGND 0.42033f 
C65342 hold75/a_49_47# VGND 0.46641f 
C65343 hold64/a_391_47# VGND 0.26257f 
C65344 hold64/a_285_47# VGND 0.41775f 
C65345 hold64/a_49_47# VGND 0.44922f 
C65346 net200 VGND 0.61454f
C65347 _0123_ VGND 0.55633f
C65348 hold53/a_391_47# VGND 0.2724f 
C65349 hold53/a_285_47# VGND 0.42949f 
C65350 hold53/a_49_47# VGND 0.47103f 
C65351 hold42/a_391_47# VGND 0.23877f 
C65352 hold42/a_285_47# VGND 0.39798f 
C65353 hold42/a_49_47# VGND 0.43626f 
C65354 net178 VGND 0.70397f
C65355 hold31/a_391_47# VGND 0.24042f 
C65356 hold31/a_285_47# VGND 0.39899f 
C65357 hold31/a_49_47# VGND 0.44143f 
C65358 hold20/a_391_47# VGND 0.26716f 
C65359 hold20/a_285_47# VGND 0.42944f 
C65360 hold20/a_49_47# VGND 0.49642f 
C65361 acc0.A\[12\] VGND 2.01292f
C65362 net39 VGND 2.62651f
C65363 _0666_/a_113_47# VGND 0.00206f 
C65364 _0092_ VGND 0.34166f
C65365 _0416_ VGND 0.30641f
C65366 _0415_ VGND 0.25266f
C65367 _0804_/a_510_47# VGND 0.00581f 
C65368 _0804_/a_215_47# VGND 0.21884f 
C65369 _0804_/a_79_21# VGND 0.34387f 
C65370 net224 VGND 0.5329f
C65371 _0735_/a_109_297# VGND 0 
C65372 clknet_0__0458_ VGND 2.93881f
C65373 clkbuf_1_0__f__0458_/a_110_47# VGND 2.28137f 
C65374 _0118_ VGND 0.62935f
C65375 _1020_/a_1017_47# VGND 0.00422f 
C65376 _1020_/a_592_47# VGND 0.00793f 
C65377 _1020_/a_975_413# VGND 0 
C65378 _1020_/a_561_413# VGND 0 
C65379 _1020_/a_381_47# VGND 0.07081f 
C65380 _1020_/a_891_413# VGND 0.27915f 
C65381 _1020_/a_1059_315# VGND 0.38622f 
C65382 _1020_/a_466_413# VGND 0.22848f 
C65383 _1020_/a_634_159# VGND 0.27723f 
C65384 _1020_/a_193_47# VGND 0.39561f 
C65385 _1020_/a_27_47# VGND 0.60952f 
C65386 net120 VGND 0.51483f
C65387 _0313_ VGND 0.88522f
C65388 _0314_ VGND 0.7827f
C65389 _0683_/a_113_47# VGND 0.00177f 
C65390 _0429_ VGND 0.48576f
C65391 _0251_ VGND 1.44693f
C65392 _0821_/a_113_47# VGND 0.00214f 
C65393 _0376_ VGND 0.25248f
C65394 _0375_ VGND 0.79819f
C65395 _0234_ VGND 0.80652f
C65396 _0752_/a_384_47# VGND 0.00456f 
C65397 _0752_/a_300_297# VGND 0.04228f 
C65398 _0752_/a_27_413# VGND 0.35675f 
C65399 _0476_ VGND 1.41277f
C65400 _0967_/a_487_297# VGND 0 
C65401 _0967_/a_403_297# VGND 0 
C65402 _0967_/a_297_297# VGND 0 
C65403 _0967_/a_215_297# VGND 0.70745f 
C65404 _0967_/a_109_93# VGND 0.25385f 
C65405 net70 VGND 0.94546f
C65406 _0984_/a_1017_47# VGND 0.0047f 
C65407 _0984_/a_592_47# VGND 0.00813f 
C65408 _0984_/a_975_413# VGND 0 
C65409 _0984_/a_561_413# VGND 0 
C65410 _0984_/a_381_47# VGND 0.07172f 
C65411 _0984_/a_891_413# VGND 0.30009f 
C65412 _0984_/a_1059_315# VGND 0.41393f 
C65413 _0984_/a_466_413# VGND 0.24689f 
C65414 _0984_/a_634_159# VGND 0.29028f 
C65415 _0984_/a_193_47# VGND 0.426f 
C65416 _0984_/a_27_47# VGND 0.6694f 
C65417 _0504_/a_27_47# VGND 0.72055f 
C65418 pp[6] VGND 0.63597f
C65419 output64/a_27_47# VGND 0.68744f 
C65420 pp[15] VGND 0.65295f
C65421 output42/a_27_47# VGND 0.47085f 
C65422 pp[25] VGND 1.16018f
C65423 net53 VGND 1.71913f
C65424 output53/a_27_47# VGND 0.45352f 
C65425 _0719_/a_27_47# VGND 0.46145f 
C65426 _1004_/a_1017_47# VGND 0.00397f 
C65427 _1004_/a_592_47# VGND 0.00748f 
C65428 _1004_/a_381_47# VGND 0.0689f 
C65429 _1004_/a_891_413# VGND 0.27807f 
C65430 _1004_/a_1059_315# VGND 0.3836f 
C65431 _1004_/a_466_413# VGND 0.21991f 
C65432 _1004_/a_634_159# VGND 0.26333f 
C65433 _1004_/a_193_47# VGND 0.37942f 
C65434 _1004_/a_27_47# VGND 0.63536f 
C65435 _0151_ VGND 0.4111f
C65436 net230 VGND 0.34255f
C65437 _0192_ VGND 0.49655f
C65438 _0521_/a_384_47# VGND 0.0036f 
C65439 _0521_/a_299_297# VGND 0.04636f 
C65440 _0521_/a_81_21# VGND 0.34022f 
C65441 net243 VGND 0.54038f
C65442 hold96/a_391_47# VGND 0.25177f 
C65443 hold96/a_285_47# VGND 0.41064f 
C65444 hold96/a_49_47# VGND 0.45678f 
C65445 net232 VGND 0.33145f
C65446 hold85/a_391_47# VGND 0.24554f 
C65447 hold85/a_285_47# VGND 0.43338f 
C65448 hold85/a_49_47# VGND 0.48735f 
C65449 hold74/a_391_47# VGND 0.25162f 
C65450 hold74/a_285_47# VGND 0.41498f 
C65451 hold74/a_49_47# VGND 0.50385f 
C65452 hold63/a_391_47# VGND 0.25722f 
C65453 hold63/a_285_47# VGND 0.42832f 
C65454 hold63/a_49_47# VGND 0.50553f 
C65455 hold52/a_391_47# VGND 0.25863f 
C65456 hold52/a_285_47# VGND 0.40503f 
C65457 hold52/a_49_47# VGND 0.46236f 
C65458 net188 VGND 0.43673f
C65459 hold41/a_391_47# VGND 0.23944f 
C65460 hold41/a_285_47# VGND 0.39641f 
C65461 hold41/a_49_47# VGND 0.44195f 
C65462 _0121_ VGND 0.26675f
C65463 hold30/a_391_47# VGND 0.2563f 
C65464 hold30/a_285_47# VGND 0.41347f 
C65465 hold30/a_49_47# VGND 0.45939f 
C65466 clknet_0__0459_ VGND 2.58104f
C65467 clkbuf_1_0__f__0459_/a_110_47# VGND 2.22211f 
C65468 _0667_/a_113_47# VGND 0.00179f 
C65469 _0230_ VGND 0.71015f
C65470 _0226_ VGND 2.36076f
C65471 _0229_ VGND 0.39412f
C65472 _0598_/a_297_47# VGND 0.17721f 
C65473 _0598_/a_382_297# VGND 0.00208f 
C65474 _0598_/a_79_21# VGND 0.28908f 
C65475 _0107_ VGND 0.55091f
C65476 _0363_ VGND 0.26863f
C65477 _0736_/a_139_47# VGND 0.00309f 
C65478 _0736_/a_311_297# VGND 0 
C65479 _0736_/a_56_297# VGND 0.03725f 
C65480 _0805_/a_181_47# VGND 0.00208f 
C65481 _0805_/a_109_47# VGND 0 
C65482 _0805_/a_27_47# VGND 0.30077f 
C65483 _0119_ VGND 0.38394f
C65484 _1021_/a_1017_47# VGND 0.00447f 
C65485 _1021_/a_592_47# VGND 0.00748f 
C65486 _1021_/a_975_413# VGND 0 
C65487 _1021_/a_381_47# VGND 0.06684f 
C65488 _1021_/a_891_413# VGND 0.29303f 
C65489 _1021_/a_1059_315# VGND 0.40649f 
C65490 _1021_/a_466_413# VGND 0.22181f 
C65491 _1021_/a_634_159# VGND 0.26701f 
C65492 _1021_/a_193_47# VGND 0.4152f 
C65493 _1021_/a_27_47# VGND 0.61626f 
C65494 _0316_ VGND 0.681f
C65495 net55 VGND 2.59879f
C65496 _0684_/a_145_75# VGND 0.00488f 
C65497 _0684_/a_59_75# VGND 0.31307f 
C65498 _0231_ VGND 1.44108f
C65499 _0233_ VGND 0.51006f
C65500 _0343_ VGND 5.07927f
C65501 _0753_/a_561_47# VGND 0.00694f 
C65502 _0753_/a_465_47# VGND 0.00338f 
C65503 _0753_/a_381_47# VGND 0.00382f 
C65504 _0753_/a_297_297# VGND 0.04362f 
C65505 _0753_/a_79_21# VGND 0.28141f 
C65506 _0430_ VGND 0.59296f
C65507 net64 VGND 2.93003f
C65508 net34 VGND 1.14325f
C65509 control0.state\[1\] VGND 1.27804f
C65510 control0.state\[0\] VGND 2.46948f
C65511 _0968_/a_193_297# VGND 0 
C65512 _0968_/a_109_297# VGND 0 
C65513 net82 VGND 0.31547f
C65514 _0390_ VGND 0.44111f
C65515 _0243_ VGND 0.70025f
C65516 _0389_ VGND 0.32744f
C65517 _0770_/a_297_47# VGND 0.21079f 
C65518 _0770_/a_382_297# VGND 0 
C65519 _0770_/a_79_21# VGND 0.29056f 
C65520 _0083_ VGND 0.36761f
C65521 _0985_/a_1017_47# VGND 0.00448f 
C65522 _0985_/a_592_47# VGND 0.00835f 
C65523 _0985_/a_975_413# VGND 0 
C65524 _0985_/a_561_413# VGND 0 
C65525 _0985_/a_381_47# VGND 0.0632f 
C65526 _0985_/a_891_413# VGND 0.2848f 
C65527 _0985_/a_1059_315# VGND 0.39164f 
C65528 _0985_/a_466_413# VGND 0.22926f 
C65529 _0985_/a_634_159# VGND 0.27464f 
C65530 _0985_/a_193_47# VGND 0.36715f 
C65531 _0985_/a_27_47# VGND 0.60831f 
C65532 net101 VGND 0.82375f
